module fake_jpeg_7864_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_41),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_1),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_51),
.B1(n_20),
.B2(n_17),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_36),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_34),
.B(n_42),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_55),
.B(n_19),
.C(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_54),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_37),
.B1(n_34),
.B2(n_28),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_57),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_69),
.B(n_64),
.C(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_70),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_89),
.B(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_86),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_21),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_72),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_1),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_101),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_46),
.C(n_42),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_107),
.C(n_104),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_113),
.B(n_120),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_82),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_111),
.B(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_123),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_119),
.C(n_83),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_90),
.C(n_79),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_93),
.B(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_125),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_81),
.CI(n_29),
.CON(n_123),
.SN(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_75),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

OAI322xp33_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_99),
.A3(n_96),
.B1(n_106),
.B2(n_109),
.C1(n_110),
.C2(n_29),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_129),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_96),
.B(n_95),
.C(n_18),
.D(n_31),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_95),
.B1(n_97),
.B2(n_75),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_134),
.B1(n_94),
.B2(n_18),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_23),
.C(n_3),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_83),
.B1(n_94),
.B2(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_117),
.C(n_119),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_142),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_116),
.C(n_113),
.Y(n_142)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_123),
.B(n_116),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_123),
.C(n_121),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_56),
.C(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_143),
.B1(n_136),
.B2(n_147),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_23),
.C(n_14),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_149),
.B(n_14),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_128),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_13),
.C(n_12),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_130),
.B1(n_137),
.B2(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_132),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_11),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_11),
.C(n_3),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_5),
.C(n_6),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_154),
.B1(n_153),
.B2(n_151),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_158),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_2),
.C(n_5),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_161),
.B(n_159),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_163),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.C(n_169),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_172),
.C(n_167),
.Y(n_177)
);


endmodule