module fake_aes_2381_n_44 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_44);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx6_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
OA21x2_ASAP7_75t_L g13 ( .A1(n_1), .A2(n_4), .B(n_2), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_7), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_4), .B(n_5), .Y(n_18) );
OR2x6_ASAP7_75t_L g19 ( .A(n_18), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_15), .B(n_6), .Y(n_21) );
NOR2xp33_ASAP7_75t_R g22 ( .A(n_12), .B(n_0), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_11), .Y(n_24) );
INVx4_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
AOI22xp33_ASAP7_75t_SL g26 ( .A1(n_19), .A2(n_14), .B1(n_16), .B2(n_13), .Y(n_26) );
CKINVDCx11_ASAP7_75t_R g27 ( .A(n_19), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_20), .A2(n_17), .B1(n_13), .B2(n_5), .C(n_6), .Y(n_28) );
AO21x2_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_21), .B(n_22), .Y(n_29) );
OAI22xp5_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_24), .B1(n_13), .B2(n_17), .Y(n_30) );
INVx1_ASAP7_75t_SL g31 ( .A(n_27), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_25), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B(n_25), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI211xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_31), .B(n_17), .C(n_23), .Y(n_37) );
O2A1O1Ixp33_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_11), .B(n_3), .C(n_2), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_36), .Y(n_39) );
HB1xp67_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
NOR2x1_ASAP7_75t_L g41 ( .A(n_38), .B(n_23), .Y(n_41) );
OR2x2_ASAP7_75t_L g42 ( .A(n_40), .B(n_23), .Y(n_42) );
BUFx2_ASAP7_75t_L g43 ( .A(n_41), .Y(n_43) );
AOI22xp5_ASAP7_75t_L g44 ( .A1(n_43), .A2(n_11), .B1(n_37), .B2(n_42), .Y(n_44) );
endmodule