module fake_jpeg_2297_n_76 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_76);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_22;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_5),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_32),
.B1(n_19),
.B2(n_20),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_42),
.C(n_35),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_11),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_44),
.B1(n_46),
.B2(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_57),
.B1(n_32),
.B2(n_31),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_22),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_34),
.B(n_35),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_56),
.B(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_64),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_63),
.B(n_26),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp67_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_62),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_72),
.B(n_22),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_65),
.A3(n_67),
.B1(n_20),
.B2(n_21),
.C1(n_16),
.C2(n_22),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.B1(n_22),
.B2(n_70),
.C(n_12),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_12),
.Y(n_76)
);


endmodule