module real_aes_8586_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g185 ( .A1(n_0), .A2(n_186), .B(n_187), .C(n_191), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_1), .B(n_181), .Y(n_192) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_3), .B(n_146), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_4), .A2(n_127), .B(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_5), .A2(n_132), .B(n_137), .C(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_6), .A2(n_127), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_7), .B(n_181), .Y(n_477) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_8), .A2(n_160), .B(n_210), .Y(n_209) );
AND2x6_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_10), .A2(n_132), .B(n_137), .C(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g532 ( .A(n_11), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_12), .B(n_40), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_13), .B(n_190), .Y(n_509) );
INVx1_ASAP7_75t_L g156 ( .A(n_14), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_15), .B(n_146), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_16), .A2(n_147), .B(n_517), .C(n_519), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_17), .B(n_181), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_18), .B(n_174), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_19), .A2(n_137), .B(n_168), .C(n_173), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_20), .A2(n_189), .B(n_204), .C(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_21), .B(n_190), .Y(n_462) );
OAI222xp33_ASAP7_75t_L g442 ( .A1(n_22), .A2(n_443), .B1(n_725), .B2(n_726), .C1(n_732), .C2(n_736), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_22), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_23), .B(n_190), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_24), .Y(n_458) );
INVx1_ASAP7_75t_L g483 ( .A(n_25), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_26), .A2(n_137), .B(n_173), .C(n_213), .Y(n_212) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_27), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_28), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_29), .Y(n_736) );
INVx1_ASAP7_75t_L g559 ( .A(n_30), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_31), .A2(n_127), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g130 ( .A(n_32), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_33), .A2(n_135), .B(n_140), .C(n_150), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_34), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_35), .A2(n_189), .B(n_474), .C(n_476), .Y(n_473) );
INVxp67_ASAP7_75t_L g560 ( .A(n_36), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_37), .B(n_215), .Y(n_214) );
CKINVDCx14_ASAP7_75t_R g472 ( .A(n_38), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_39), .A2(n_137), .B(n_173), .C(n_482), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_41), .A2(n_191), .B(n_530), .C(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_42), .B(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_43), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_44), .B(n_146), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_45), .B(n_127), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_46), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_47), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_48), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_49), .A2(n_135), .B(n_150), .C(n_224), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_50), .A2(n_118), .B1(n_119), .B2(n_437), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g188 ( .A(n_51), .Y(n_188) );
INVx1_ASAP7_75t_L g225 ( .A(n_52), .Y(n_225) );
INVx1_ASAP7_75t_L g495 ( .A(n_53), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_54), .B(n_127), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_55), .Y(n_177) );
CKINVDCx14_ASAP7_75t_R g528 ( .A(n_56), .Y(n_528) );
INVx1_ASAP7_75t_L g133 ( .A(n_57), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_58), .B(n_127), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_59), .B(n_181), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_60), .A2(n_172), .B(n_235), .C(n_237), .Y(n_234) );
INVx1_ASAP7_75t_L g155 ( .A(n_61), .Y(n_155) );
INVx1_ASAP7_75t_SL g475 ( .A(n_62), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_64), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_65), .B(n_181), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_66), .B(n_147), .Y(n_201) );
INVx1_ASAP7_75t_L g461 ( .A(n_67), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_68), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_69), .B(n_143), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_70), .A2(n_137), .B(n_150), .C(n_261), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_71), .Y(n_233) );
INVx1_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_73), .A2(n_127), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_74), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_75), .A2(n_127), .B(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_76), .A2(n_166), .B(n_555), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_77), .Y(n_480) );
INVx1_ASAP7_75t_L g515 ( .A(n_78), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_79), .B(n_142), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_80), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_81), .A2(n_127), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g518 ( .A(n_82), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_83), .A2(n_100), .B1(n_111), .B2(n_739), .Y(n_99) );
INVx2_ASAP7_75t_L g153 ( .A(n_84), .Y(n_153) );
INVx1_ASAP7_75t_L g508 ( .A(n_85), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_86), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_87), .B(n_190), .Y(n_202) );
OR2x2_ASAP7_75t_L g106 ( .A(n_88), .B(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g445 ( .A(n_88), .B(n_108), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_88), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_89), .A2(n_137), .B(n_150), .C(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_90), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
INVxp67_ASAP7_75t_L g238 ( .A(n_92), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_93), .B(n_160), .Y(n_533) );
INVx2_ASAP7_75t_L g498 ( .A(n_94), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_95), .B(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g197 ( .A(n_96), .Y(n_197) );
INVx1_ASAP7_75t_L g262 ( .A(n_97), .Y(n_262) );
AND2x2_ASAP7_75t_L g227 ( .A(n_98), .B(n_152), .Y(n_227) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g740 ( .A(n_101), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_105), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_106), .Y(n_438) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_107), .B(n_448), .Y(n_735) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g447 ( .A(n_108), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OAI21x1_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_116), .B(n_441), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g738 ( .A(n_114), .Y(n_738) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_438), .B(n_439), .Y(n_116) );
INVx2_ASAP7_75t_L g437 ( .A(n_119), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_119), .A2(n_727), .B1(n_730), .B2(n_731), .Y(n_726) );
OR3x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_351), .C(n_394), .Y(n_119) );
NAND5xp2_ASAP7_75t_L g120 ( .A(n_121), .B(n_278), .C(n_308), .D(n_325), .E(n_340), .Y(n_120) );
AOI221xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_193), .B1(n_240), .B2(n_246), .C(n_250), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_162), .Y(n_122) );
OR2x2_ASAP7_75t_L g255 ( .A(n_123), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g295 ( .A(n_123), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_123), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_123), .B(n_248), .Y(n_330) );
OR2x2_ASAP7_75t_L g342 ( .A(n_123), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_123), .B(n_301), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_123), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_123), .B(n_279), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_123), .B(n_287), .Y(n_393) );
AND2x2_ASAP7_75t_L g425 ( .A(n_123), .B(n_179), .Y(n_425) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_123), .Y(n_433) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_124), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g252 ( .A(n_124), .B(n_228), .Y(n_252) );
BUFx2_ASAP7_75t_L g275 ( .A(n_124), .Y(n_275) );
AND2x2_ASAP7_75t_L g304 ( .A(n_124), .B(n_163), .Y(n_304) );
AND2x2_ASAP7_75t_L g359 ( .A(n_124), .B(n_256), .Y(n_359) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_157), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_134), .B(n_152), .Y(n_125) );
BUFx2_ASAP7_75t_L g166 ( .A(n_127), .Y(n_166) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_128), .B(n_132), .Y(n_198) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
INVx1_ASAP7_75t_L g205 ( .A(n_130), .Y(n_205) );
INVx1_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
INVx3_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
INVx1_ASAP7_75t_L g215 ( .A(n_131), .Y(n_215) );
INVx4_ASAP7_75t_SL g151 ( .A(n_132), .Y(n_151) );
BUFx3_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_SL g183 ( .A1(n_136), .A2(n_151), .B(n_184), .C(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_136), .A2(n_151), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_136), .A2(n_151), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_136), .A2(n_151), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_136), .A2(n_151), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_136), .A2(n_151), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_136), .A2(n_151), .B(n_556), .C(n_557), .Y(n_555) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx3_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_138), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_145), .C(n_148), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_142), .A2(n_148), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_142), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
O2A1O1Ixp5_ASAP7_75t_L g507 ( .A1(n_142), .A2(n_463), .B(n_508), .C(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g236 ( .A(n_144), .Y(n_236) );
INVx2_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_146), .B(n_238), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_146), .A2(n_171), .B(n_483), .C(n_484), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_146), .A2(n_236), .B1(n_559), .B2(n_560), .Y(n_558) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_147), .B(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx1_ASAP7_75t_L g519 ( .A(n_149), .Y(n_519) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
INVx1_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_152), .A2(n_222), .B(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_152), .A2(n_198), .B(n_480), .C(n_481), .Y(n_479) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_152), .A2(n_526), .B(n_533), .Y(n_525) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_153), .B(n_154), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx3_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_159), .A2(n_196), .B(n_206), .Y(n_195) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_159), .A2(n_259), .B(n_267), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_159), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_159), .A2(n_457), .B(n_464), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_159), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_159), .B(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_211), .B(n_212), .Y(n_210) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_162), .B(n_313), .Y(n_322) );
OAI32xp33_ASAP7_75t_L g336 ( .A1(n_162), .A2(n_272), .A3(n_337), .B1(n_338), .B2(n_339), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_162), .B(n_338), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_162), .B(n_255), .Y(n_379) );
INVx1_ASAP7_75t_SL g408 ( .A(n_162), .Y(n_408) );
NAND4xp25_ASAP7_75t_L g417 ( .A(n_162), .B(n_195), .C(n_359), .D(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_179), .Y(n_162) );
INVx5_ASAP7_75t_L g249 ( .A(n_163), .Y(n_249) );
AND2x2_ASAP7_75t_L g279 ( .A(n_163), .B(n_180), .Y(n_279) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_163), .Y(n_358) );
AND2x2_ASAP7_75t_L g428 ( .A(n_163), .B(n_375), .Y(n_428) );
OR2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_176), .Y(n_163) );
AOI21xp5_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_167), .B(n_174), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .Y(n_168) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_172), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_175), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_178), .A2(n_504), .B(n_510), .Y(n_503) );
AND2x4_ASAP7_75t_L g301 ( .A(n_179), .B(n_249), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_179), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g335 ( .A(n_179), .B(n_256), .Y(n_335) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g248 ( .A(n_180), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g287 ( .A(n_180), .B(n_258), .Y(n_287) );
AND2x2_ASAP7_75t_L g296 ( .A(n_180), .B(n_257), .Y(n_296) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_192), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_189), .B(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g530 ( .A(n_190), .Y(n_530) );
INVx2_ASAP7_75t_L g463 ( .A(n_191), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_193), .A2(n_365), .B1(n_367), .B2(n_369), .C1(n_372), .C2(n_373), .Y(n_364) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_217), .Y(n_193) );
AND2x2_ASAP7_75t_L g297 ( .A(n_194), .B(n_298), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_194), .B(n_275), .C(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_209), .Y(n_194) );
INVx5_ASAP7_75t_SL g245 ( .A(n_195), .Y(n_245) );
OAI322xp33_ASAP7_75t_L g250 ( .A1(n_195), .A2(n_251), .A3(n_253), .B1(n_254), .B2(n_269), .C1(n_272), .C2(n_274), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_195), .B(n_243), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_195), .B(n_229), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_198), .A2(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_198), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_203), .A2(n_214), .B(n_216), .Y(n_213) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g553 ( .A(n_208), .Y(n_553) );
INVx2_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_209), .B(n_219), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_217), .B(n_282), .Y(n_337) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g316 ( .A(n_218), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
OR2x2_ASAP7_75t_L g244 ( .A(n_219), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_219), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g284 ( .A(n_219), .B(n_229), .Y(n_284) );
AND2x2_ASAP7_75t_L g307 ( .A(n_219), .B(n_243), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_219), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g323 ( .A(n_219), .B(n_282), .Y(n_323) );
AND2x2_ASAP7_75t_L g331 ( .A(n_219), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_219), .B(n_291), .Y(n_381) );
INVx5_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g271 ( .A(n_220), .B(n_245), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_220), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g298 ( .A(n_220), .B(n_229), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_220), .B(n_345), .Y(n_386) );
OR2x2_ASAP7_75t_L g402 ( .A(n_220), .B(n_346), .Y(n_402) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_220), .B(n_363), .Y(n_409) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_220), .Y(n_416) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
AND2x2_ASAP7_75t_L g270 ( .A(n_228), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g320 ( .A(n_228), .B(n_243), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_228), .B(n_245), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_228), .B(n_282), .Y(n_404) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_229), .B(n_245), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_229), .B(n_243), .Y(n_292) );
OR2x2_ASAP7_75t_L g346 ( .A(n_229), .B(n_243), .Y(n_346) );
AND2x2_ASAP7_75t_L g363 ( .A(n_229), .B(n_242), .Y(n_363) );
INVxp67_ASAP7_75t_L g385 ( .A(n_229), .Y(n_385) );
AND2x2_ASAP7_75t_L g412 ( .A(n_229), .B(n_282), .Y(n_412) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_229), .Y(n_419) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_230), .A2(n_470), .B(n_477), .Y(n_469) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_230), .A2(n_493), .B(n_499), .Y(n_492) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_230), .A2(n_513), .B(n_520), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_235), .A2(n_262), .B(n_263), .C(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_236), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_236), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_242), .B(n_293), .Y(n_366) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g282 ( .A(n_243), .B(n_245), .Y(n_282) );
OR2x2_ASAP7_75t_L g349 ( .A(n_243), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g293 ( .A(n_244), .Y(n_293) );
OR2x2_ASAP7_75t_L g354 ( .A(n_244), .B(n_346), .Y(n_354) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g253 ( .A(n_248), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_248), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g254 ( .A(n_249), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_249), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_249), .B(n_256), .Y(n_289) );
INVx2_ASAP7_75t_L g334 ( .A(n_249), .Y(n_334) );
AND2x2_ASAP7_75t_L g347 ( .A(n_249), .B(n_287), .Y(n_347) );
AND2x2_ASAP7_75t_L g372 ( .A(n_249), .B(n_296), .Y(n_372) );
INVx1_ASAP7_75t_L g324 ( .A(n_254), .Y(n_324) );
INVx2_ASAP7_75t_SL g311 ( .A(n_255), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g375 ( .A(n_258), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_266), .Y(n_259) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g476 ( .A(n_265), .Y(n_476) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g344 ( .A(n_271), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g350 ( .A(n_271), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_271), .A2(n_353), .B1(n_355), .B2(n_360), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_271), .B(n_363), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_272), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g306 ( .A(n_273), .Y(n_306) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g288 ( .A(n_275), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_275), .B(n_279), .Y(n_339) );
AND2x2_ASAP7_75t_L g362 ( .A(n_275), .B(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g338 ( .A(n_277), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_285), .C(n_299), .Y(n_278) );
INVx1_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_279), .A2(n_411), .B1(n_413), .B2(n_414), .C(n_417), .Y(n_410) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g429 ( .A(n_282), .Y(n_429) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g378 ( .A(n_284), .B(n_317), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B(n_290), .C(n_294), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI32xp33_ASAP7_75t_L g403 ( .A1(n_292), .A2(n_293), .A3(n_356), .B1(n_393), .B2(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x2_ASAP7_75t_L g435 ( .A(n_295), .B(n_334), .Y(n_435) );
AND2x2_ASAP7_75t_L g382 ( .A(n_296), .B(n_334), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_296), .B(n_304), .Y(n_400) );
AOI31xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .A3(n_303), .B(n_305), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_301), .B(n_313), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_301), .B(n_311), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_301), .A2(n_331), .B1(n_421), .B2(n_424), .C(n_426), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g326 ( .A(n_306), .B(n_327), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_315), .B1(n_318), .B2(n_321), .C1(n_323), .C2(n_324), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g391 ( .A(n_310), .Y(n_391) );
INVx1_ASAP7_75t_L g413 ( .A(n_313), .Y(n_413) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_316), .A2(n_427), .B1(n_429), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g332 ( .A(n_317), .Y(n_332) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_336), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g370 ( .A(n_328), .B(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g422 ( .A(n_328), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g397 ( .A(n_333), .Y(n_397) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g361 ( .A(n_334), .Y(n_361) );
INVx1_ASAP7_75t_L g343 ( .A(n_335), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_338), .B(n_425), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_347), .B2(n_348), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g434 ( .A(n_347), .Y(n_434) );
INVxp33_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_349), .B(n_393), .Y(n_392) );
OAI32xp33_ASAP7_75t_L g383 ( .A1(n_350), .A2(n_384), .A3(n_385), .B1(n_386), .B2(n_387), .Y(n_383) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_364), .C(n_376), .D(n_388), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
NAND2xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_359), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
CKINVDCx16_ASAP7_75t_R g369 ( .A(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_373), .A2(n_389), .B1(n_406), .B2(n_409), .C(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g424 ( .A(n_375), .B(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B1(n_380), .B2(n_382), .C(n_383), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_385), .B(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_405), .C(n_420), .D(n_431), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B(n_401), .C(n_403), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g436 ( .A(n_423), .Y(n_436) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_436), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_437), .A2(n_444), .B1(n_446), .B2(n_449), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g439 ( .A(n_438), .B(n_440), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_439), .A2(n_442), .B(n_737), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g729 ( .A(n_445), .Y(n_729) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx6_ASAP7_75t_L g730 ( .A(n_447), .Y(n_730) );
INVx3_ASAP7_75t_L g731 ( .A(n_449), .Y(n_731) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_450), .B(n_680), .Y(n_449) );
NOR4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_617), .C(n_651), .D(n_667), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_546), .C(n_581), .D(n_597), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_487), .B1(n_521), .B2(n_534), .C1(n_539), .C2(n_545), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI31xp33_ASAP7_75t_L g713 ( .A1(n_454), .A2(n_714), .A3(n_715), .B(n_717), .Y(n_713) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
AND2x2_ASAP7_75t_L g688 ( .A(n_455), .B(n_468), .Y(n_688) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g538 ( .A(n_456), .Y(n_538) );
AND2x2_ASAP7_75t_L g545 ( .A(n_456), .B(n_478), .Y(n_545) );
AND2x2_ASAP7_75t_L g602 ( .A(n_456), .B(n_469), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_466), .B(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_467), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_467), .B(n_549), .Y(n_592) );
AND2x2_ASAP7_75t_L g685 ( .A(n_467), .B(n_625), .Y(n_685) );
OAI321xp33_ASAP7_75t_L g719 ( .A1(n_467), .A2(n_538), .A3(n_692), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g723 ( .A(n_467), .B(n_524), .C(n_632), .D(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g587 ( .A(n_468), .B(n_536), .Y(n_587) );
AND2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_538), .Y(n_606) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g537 ( .A(n_469), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g562 ( .A(n_469), .B(n_478), .Y(n_562) );
AND2x2_ASAP7_75t_L g648 ( .A(n_469), .B(n_536), .Y(n_648) );
INVx3_ASAP7_75t_SL g536 ( .A(n_478), .Y(n_536) );
AND2x2_ASAP7_75t_L g580 ( .A(n_478), .B(n_567), .Y(n_580) );
OR2x2_ASAP7_75t_L g613 ( .A(n_478), .B(n_538), .Y(n_613) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_478), .Y(n_620) );
AND2x2_ASAP7_75t_L g649 ( .A(n_478), .B(n_537), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_478), .B(n_622), .Y(n_664) );
AND2x2_ASAP7_75t_L g696 ( .A(n_478), .B(n_688), .Y(n_696) );
AND2x2_ASAP7_75t_L g705 ( .A(n_478), .B(n_550), .Y(n_705) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_485), .Y(n_478) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
INVx1_ASAP7_75t_SL g673 ( .A(n_489), .Y(n_673) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g541 ( .A(n_490), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g523 ( .A(n_491), .B(n_502), .Y(n_523) );
AND2x2_ASAP7_75t_L g609 ( .A(n_491), .B(n_525), .Y(n_609) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_512), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_492), .B(n_525), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_492), .B(n_525), .Y(n_616) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_492), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_500), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_500), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g589 ( .A(n_501), .B(n_590), .Y(n_589) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_501), .A2(n_579), .A3(n_585), .B1(n_616), .B2(n_666), .C1(n_676), .C2(n_678), .Y(n_675) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_502), .B(n_524), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_502), .B(n_525), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_502), .B(n_542), .Y(n_596) );
AND2x2_ASAP7_75t_L g650 ( .A(n_502), .B(n_616), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_502), .Y(n_654) );
AND2x2_ASAP7_75t_L g666 ( .A(n_502), .B(n_512), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_502), .B(n_541), .Y(n_698) );
INVx4_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g563 ( .A(n_503), .B(n_512), .Y(n_563) );
BUFx3_ASAP7_75t_L g577 ( .A(n_503), .Y(n_577) );
AND3x2_ASAP7_75t_L g659 ( .A(n_503), .B(n_639), .C(n_660), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_512), .B(n_523), .C(n_524), .Y(n_522) );
INVx1_ASAP7_75t_SL g542 ( .A(n_512), .Y(n_542) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_512), .Y(n_644) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g638 ( .A(n_523), .B(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g645 ( .A(n_523), .Y(n_645) );
AND2x2_ASAP7_75t_L g683 ( .A(n_524), .B(n_661), .Y(n_683) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g564 ( .A(n_525), .Y(n_564) );
AND2x2_ASAP7_75t_L g639 ( .A(n_525), .B(n_542), .Y(n_639) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OR2x2_ASAP7_75t_L g583 ( .A(n_536), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g702 ( .A(n_536), .B(n_602), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_536), .B(n_538), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_537), .B(n_550), .Y(n_657) );
AND2x2_ASAP7_75t_L g704 ( .A(n_537), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g567 ( .A(n_538), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g584 ( .A(n_538), .B(n_550), .Y(n_584) );
INVx1_ASAP7_75t_L g594 ( .A(n_538), .Y(n_594) );
AND2x2_ASAP7_75t_L g625 ( .A(n_538), .B(n_550), .Y(n_625) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_540), .A2(n_668), .B1(n_672), .B2(n_674), .C(n_675), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x2_ASAP7_75t_L g571 ( .A(n_541), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_544), .B(n_578), .Y(n_721) );
AOI322xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_563), .A3(n_564), .B1(n_565), .B2(n_571), .C1(n_573), .C2(n_580), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_562), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_549), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_549), .B(n_612), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_549), .A2(n_562), .B(n_636), .C(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_549), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_549), .B(n_606), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_549), .B(n_688), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_549), .B(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_550), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_550), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g677 ( .A(n_550), .B(n_564), .Y(n_677) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_554), .B(n_561), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_552), .A2(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g569 ( .A(n_554), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_561), .Y(n_570) );
INVx1_ASAP7_75t_L g652 ( .A(n_562), .Y(n_652) );
OAI31xp33_ASAP7_75t_L g662 ( .A1(n_562), .A2(n_587), .A3(n_663), .B(n_665), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_562), .B(n_568), .Y(n_714) );
INVx1_ASAP7_75t_SL g575 ( .A(n_563), .Y(n_575) );
AND2x2_ASAP7_75t_L g608 ( .A(n_563), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g689 ( .A(n_563), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g574 ( .A(n_564), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g599 ( .A(n_564), .Y(n_599) );
AND2x2_ASAP7_75t_L g626 ( .A(n_564), .B(n_579), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_564), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g718 ( .A(n_564), .B(n_666), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_566), .B(n_636), .Y(n_709) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g605 ( .A(n_568), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g623 ( .A(n_568), .Y(n_623) );
NAND2xp33_ASAP7_75t_SL g573 ( .A(n_574), .B(n_576), .Y(n_573) );
OAI211xp5_ASAP7_75t_SL g617 ( .A1(n_575), .A2(n_618), .B(n_624), .C(n_640), .Y(n_617) );
OR2x2_ASAP7_75t_L g692 ( .A(n_575), .B(n_673), .Y(n_692) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
CKINVDCx16_ASAP7_75t_R g629 ( .A(n_577), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_577), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g598 ( .A(n_579), .B(n_599), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_588), .C(n_591), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g632 ( .A(n_584), .Y(n_632) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_587), .B(n_625), .Y(n_630) );
INVx1_ASAP7_75t_L g636 ( .A(n_587), .Y(n_636) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g595 ( .A(n_590), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g628 ( .A(n_590), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g690 ( .A(n_590), .Y(n_690) );
AOI21xp33_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B(n_595), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_593), .A2(n_604), .B(n_607), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_603), .C(n_610), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_598), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_601), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g614 ( .A(n_602), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_604), .A2(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_609), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g634 ( .A(n_609), .Y(n_634) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_614), .B(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g665 ( .A(n_616), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_622), .B(n_648), .Y(n_674) );
AND2x2_ASAP7_75t_L g687 ( .A(n_622), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g701 ( .A(n_622), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g711 ( .A(n_622), .B(n_649), .Y(n_711) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_627), .C(n_635), .Y(n_624) );
INVx1_ASAP7_75t_L g671 ( .A(n_625), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B1(n_631), .B2(n_633), .Y(n_627) );
OR2x2_ASAP7_75t_L g633 ( .A(n_629), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_629), .B(n_690), .Y(n_712) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g706 ( .A(n_639), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_646), .B1(n_649), .B2(n_650), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g724 ( .A(n_644), .Y(n_724) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g670 ( .A(n_648), .Y(n_670) );
OAI211xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_655), .C(n_662), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_670), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR5xp2_ASAP7_75t_L g680 ( .A(n_681), .B(n_699), .C(n_707), .D(n_713), .E(n_719), .Y(n_680) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_684), .B(n_686), .C(n_693), .Y(n_681) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_691), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_696), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B(n_706), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g722 ( .A(n_702), .Y(n_722) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
endmodule