module fake_jpeg_16948_n_294 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_15),
.Y(n_45)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_29),
.Y(n_82)
);

NAND2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_35),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_41),
.B1(n_26),
.B2(n_25),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_76)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_34),
.B1(n_36),
.B2(n_16),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_30),
.B1(n_24),
.B2(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_68),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_38),
.B1(n_37),
.B2(n_28),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_75),
.B1(n_83),
.B2(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_82),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_32),
.B1(n_38),
.B2(n_28),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_37),
.B1(n_15),
.B2(n_21),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_79),
.B(n_26),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_32),
.B1(n_18),
.B2(n_25),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_9),
.B1(n_14),
.B2(n_12),
.Y(n_86)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

XNOR2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_42),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_106),
.B(n_86),
.C(n_68),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_109),
.B1(n_89),
.B2(n_56),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_45),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_112),
.C(n_80),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_26),
.B(n_50),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_83),
.B(n_26),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_64),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_103),
.B1(n_89),
.B2(n_67),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_60),
.B(n_41),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_113),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_44),
.B1(n_49),
.B2(n_47),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_44),
.B1(n_55),
.B2(n_63),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_119),
.B1(n_90),
.B2(n_114),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_110),
.B1(n_113),
.B2(n_92),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_111),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_130),
.B1(n_135),
.B2(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_131),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_100),
.C(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_81),
.B1(n_44),
.B2(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_98),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_67),
.B1(n_87),
.B2(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_82),
.B1(n_56),
.B2(n_59),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_99),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_114),
.B1(n_90),
.B2(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_127),
.B1(n_130),
.B2(n_128),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_144),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_151),
.B1(n_161),
.B2(n_163),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_164),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_126),
.B1(n_123),
.B2(n_119),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_120),
.B(n_132),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_112),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_112),
.B(n_98),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_87),
.B1(n_63),
.B2(n_78),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_59),
.B1(n_62),
.B2(n_67),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_106),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

BUFx4f_ASAP7_75t_SL g206 ( 
.A(n_166),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_142),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_173),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_181),
.B(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_140),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_132),
.B(n_134),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_137),
.B(n_121),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_135),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_144),
.C(n_151),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_121),
.B1(n_138),
.B2(n_115),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_163),
.B1(n_142),
.B2(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_140),
.B(n_139),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_207),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_186),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_122),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_209),
.C(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_141),
.B(n_158),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_203),
.B(n_176),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_154),
.B(n_158),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_156),
.B(n_158),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_150),
.B(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_210),
.B1(n_184),
.B2(n_169),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_142),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_159),
.B(n_102),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_102),
.C(n_84),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_169),
.B1(n_178),
.B2(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_216),
.B1(n_205),
.B2(n_200),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_172),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_192),
.C(n_210),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_201),
.B1(n_203),
.B2(n_193),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_177),
.B1(n_180),
.B2(n_188),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_167),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_177),
.C(n_166),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_209),
.C(n_195),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_122),
.C(n_48),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_48),
.C(n_176),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_208),
.C(n_190),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_226),
.Y(n_248)
);

BUFx4f_ASAP7_75t_SL g234 ( 
.A(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_235),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_237),
.C(n_239),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_192),
.C(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_191),
.C(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_194),
.CI(n_196),
.CON(n_242),
.SN(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_196),
.C(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_206),
.C(n_194),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_71),
.C(n_2),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_248),
.B(n_251),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_220),
.B1(n_217),
.B2(n_206),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_3),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_217),
.B1(n_219),
.B2(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_225),
.B1(n_212),
.B2(n_43),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_1),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_260),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_1),
.C(n_3),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_245),
.B(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_256),
.C(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_239),
.B1(n_246),
.B2(n_242),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_12),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_269),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_7),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_271),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_7),
.B(n_10),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_248),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_267),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_279),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_256),
.C(n_258),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_270),
.B1(n_249),
.B2(n_269),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_273),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_280),
.A2(n_11),
.B(n_6),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_284),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_4),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C1(n_287),
.C2(n_291),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_10),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_4),
.Y(n_294)
);


endmodule