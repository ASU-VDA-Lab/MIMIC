module fake_netlist_6_4474_n_2044 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2044);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2044;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_873;
wire n_461;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1737;
wire n_236;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_80),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_33),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_115),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_78),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_0),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_91),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_23),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_32),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_102),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_10),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_52),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_78),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_28),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_124),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_60),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_37),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_172),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_167),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_51),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_38),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_89),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_17),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_30),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_26),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_93),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_100),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_112),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_104),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_210),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_73),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_189),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_86),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_181),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_157),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_205),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_208),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_54),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_158),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_68),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_119),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_10),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_106),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_25),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_34),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_55),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_79),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_168),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_50),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_92),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_175),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_171),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_117),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_120),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_107),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_37),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_26),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_137),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_190),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_94),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_56),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_101),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_150),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_194),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_4),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_122),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_191),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_35),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_87),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_56),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_32),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_183),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_17),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_73),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_69),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_64),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_67),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_138),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_77),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_63),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_133),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_13),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_83),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_201),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_193),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_67),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_27),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_7),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_19),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_31),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_109),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_47),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_188),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_42),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_72),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_209),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_86),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_114),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_125),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_127),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_166),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_121),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_173),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_12),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_108),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_6),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_33),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_77),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_90),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_39),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_47),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_64),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_57),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_51),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_75),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_58),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_55),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_58),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_60),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_98),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_99),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_20),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_68),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_155),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_144),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_159),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_28),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_57),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_80),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_162),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_96),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_118),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_6),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_126),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_149),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_195),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_76),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_143),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_146),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_165),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_12),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_70),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_178),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_36),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_81),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_1),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_35),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_185),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_25),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_4),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_123),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_179),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_52),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_74),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_197),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_82),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_48),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_11),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_132),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_11),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_59),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_131),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_186),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_202),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_142),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_177),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_53),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_164),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_38),
.Y(n_411)
);

CKINVDCx11_ASAP7_75t_R g412 ( 
.A(n_180),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_40),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_34),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_255),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_412),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_214),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_267),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_230),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_347),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_326),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_347),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_217),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_283),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_347),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_284),
.B(n_0),
.Y(n_429)
);

INVxp33_ASAP7_75t_SL g430 ( 
.A(n_320),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_220),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_374),
.B(n_2),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_320),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_411),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_318),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_222),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_260),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_329),
.B(n_270),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g444 ( 
.A(n_271),
.B(n_3),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_235),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_236),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_232),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_369),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_238),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_336),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_408),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_241),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_243),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_244),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_249),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_212),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_260),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_251),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_270),
.B(n_3),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_254),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_254),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_254),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_262),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_257),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_258),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_401),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_224),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_268),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_313),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_313),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_313),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_269),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_272),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_232),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_237),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_237),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_252),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_276),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_278),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_226),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_252),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_262),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_401),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_362),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_253),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_213),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_286),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_253),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_287),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_273),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_273),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_362),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_275),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_213),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_288),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_215),
.B(n_5),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_248),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_274),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_275),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_289),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_291),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_221),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_227),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_292),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_281),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_281),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_282),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_282),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_271),
.B(n_5),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_295),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_285),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_297),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_301),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_302),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_285),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_306),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_215),
.B(n_8),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_312),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_303),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_324),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_303),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_316),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_316),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_335),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_335),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_344),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_418),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_417),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_508),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_508),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_472),
.B(n_325),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_460),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_426),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_420),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_422),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_433),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_443),
.B(n_305),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_444),
.B(n_263),
.Y(n_548)
);

INVxp33_ASAP7_75t_SL g549 ( 
.A(n_416),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_427),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

AND3x2_ASAP7_75t_L g552 ( 
.A(n_464),
.B(n_311),
.C(n_263),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_425),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_492),
.B(n_263),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g557 ( 
.A1(n_428),
.A2(n_331),
.B(n_311),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_500),
.B(n_311),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_439),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_428),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_489),
.B(n_466),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_431),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_436),
.B(n_317),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_432),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_466),
.B(n_331),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_438),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_446),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_424),
.Y(n_570)
);

BUFx8_ASAP7_75t_L g571 ( 
.A(n_441),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_419),
.B(n_246),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_453),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_486),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_432),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_447),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_434),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_467),
.B(n_331),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_452),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_434),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_437),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_467),
.B(n_397),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_437),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_442),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_455),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_442),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_445),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_449),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_457),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_454),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_462),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_468),
.B(n_333),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_504),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_480),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_450),
.B(n_397),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_468),
.B(n_397),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_458),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_481),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_503),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_506),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_450),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_459),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_481),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_463),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_482),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_509),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_470),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_471),
.B(n_339),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_510),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_516),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_451),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_451),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_429),
.B(n_246),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_456),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_482),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_502),
.B(n_305),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_515),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_518),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_440),
.B(n_296),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_537),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_617),
.B(n_435),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_621),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_617),
.B(n_474),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_612),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_572),
.B(n_469),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_621),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_478),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_571),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_603),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_571),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_557),
.B(n_296),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_591),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_533),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_533),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_547),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_538),
.B(n_479),
.Y(n_641)
);

CKINVDCx6p67_ASAP7_75t_R g642 ( 
.A(n_603),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_556),
.B(n_441),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_604),
.Y(n_644)
);

INVx4_ASAP7_75t_SL g645 ( 
.A(n_547),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_612),
.B(n_498),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_613),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_597),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

INVxp33_ASAP7_75t_SL g651 ( 
.A(n_539),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_556),
.A2(n_558),
.B1(n_620),
.B2(n_548),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_536),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_538),
.B(n_484),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_547),
.B(n_485),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_623),
.A2(n_610),
.B1(n_526),
.B2(n_415),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_543),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_539),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_537),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_548),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_541),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_556),
.B(n_475),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_547),
.B(n_558),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_542),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_547),
.B(n_558),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_548),
.B(n_561),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_610),
.A2(n_564),
.B1(n_574),
.B2(n_569),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_542),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_566),
.B(n_475),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_545),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_493),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_602),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_620),
.B(n_305),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_548),
.B(n_317),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_547),
.B(n_495),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_547),
.B(n_501),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_566),
.B(n_476),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_571),
.Y(n_680)
);

INVx4_ASAP7_75t_SL g681 ( 
.A(n_547),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_566),
.B(n_476),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_578),
.B(n_477),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_569),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_620),
.A2(n_430),
.B1(n_523),
.B2(n_379),
.Y(n_685)
);

AO22x2_ASAP7_75t_L g686 ( 
.A1(n_578),
.A2(n_379),
.B1(n_259),
.B2(n_223),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_548),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_540),
.B(n_507),
.Y(n_688)
);

CKINVDCx16_ASAP7_75t_R g689 ( 
.A(n_550),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_544),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_602),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_578),
.B(n_477),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_594),
.B(n_519),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_574),
.A2(n_522),
.B1(n_524),
.B2(n_520),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_571),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_545),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_594),
.B(n_561),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_548),
.B(n_448),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_SL g699 ( 
.A(n_546),
.B(n_490),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_559),
.B(n_340),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_607),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_552),
.B(n_342),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_568),
.B(n_341),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_537),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_595),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_537),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_544),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_576),
.B(n_525),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_551),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_593),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_570),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_552),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_579),
.A2(n_342),
.B1(n_218),
.B2(n_343),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_585),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_590),
.B(n_601),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_609),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_606),
.B(n_345),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_608),
.B(n_349),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_537),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_609),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_551),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_619),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_537),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_571),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_611),
.B(n_229),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_619),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_570),
.B(n_223),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_537),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_582),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_588),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_588),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_549),
.B(n_366),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_582),
.B(n_234),
.C(n_231),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_600),
.B(n_598),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_553),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_553),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_620),
.B(n_368),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_553),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_593),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_599),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_599),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_620),
.B(n_373),
.Y(n_744)
);

BUFx8_ASAP7_75t_SL g745 ( 
.A(n_567),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_600),
.A2(n_259),
.B1(n_240),
.B2(n_247),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_555),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_555),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_555),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_600),
.B(n_376),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_563),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_598),
.B(n_456),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_562),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_535),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_563),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_598),
.B(n_250),
.C(n_239),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_575),
.B(n_261),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_575),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_577),
.B(n_264),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_620),
.B(n_380),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_588),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_577),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_598),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_SL g764 ( 
.A(n_614),
.B(n_277),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_588),
.Y(n_765)
);

AND3x2_ASAP7_75t_L g766 ( 
.A(n_598),
.B(n_219),
.C(n_216),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_588),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_557),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_580),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_580),
.B(n_381),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_562),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_730),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_736),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_712),
.B(n_216),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_625),
.A2(n_557),
.B1(n_225),
.B2(n_228),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_627),
.B(n_631),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_641),
.B(n_535),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_730),
.B(n_535),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_685),
.A2(n_402),
.B1(n_400),
.B2(n_398),
.C(n_360),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_SL g780 ( 
.A(n_640),
.B(n_305),
.Y(n_780)
);

BUFx4f_ASAP7_75t_L g781 ( 
.A(n_667),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_625),
.B(n_382),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_736),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_697),
.B(n_535),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_628),
.B(n_385),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_697),
.B(n_583),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_736),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_752),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_654),
.B(n_622),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_652),
.B(n_583),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_693),
.B(n_573),
.Y(n_791)
);

AND2x6_ASAP7_75t_L g792 ( 
.A(n_633),
.B(n_219),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_643),
.B(n_586),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_664),
.A2(n_557),
.B1(n_225),
.B2(n_233),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_708),
.B(n_592),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_628),
.B(n_393),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_643),
.B(n_586),
.Y(n_797)
);

AND2x2_ASAP7_75t_SL g798 ( 
.A(n_675),
.B(n_305),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_663),
.B(n_616),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_663),
.B(n_587),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_666),
.A2(n_557),
.B1(n_228),
.B2(n_242),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_634),
.A2(n_414),
.B1(n_395),
.B2(n_356),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_752),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_SL g804 ( 
.A(n_712),
.B(n_307),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_632),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_SL g806 ( 
.A1(n_657),
.A2(n_319),
.B1(n_310),
.B2(n_370),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_634),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_642),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_716),
.B(n_616),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_660),
.A2(n_290),
.B1(n_378),
.B2(n_377),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_670),
.B(n_587),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_735),
.B(n_630),
.C(n_626),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_660),
.A2(n_233),
.B(n_377),
.C(n_242),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_679),
.B(n_682),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_637),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_626),
.B(n_394),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_679),
.B(n_616),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_632),
.Y(n_818)
);

O2A1O1Ixp5_ASAP7_75t_L g819 ( 
.A1(n_739),
.A2(n_560),
.B(n_565),
.C(n_372),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_630),
.B(n_265),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_682),
.B(n_560),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_653),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_763),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_653),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_684),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_683),
.B(n_560),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_656),
.B(n_404),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_649),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_726),
.B(n_266),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_684),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_698),
.B(n_405),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_661),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_662),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_683),
.B(n_560),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_662),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_692),
.B(n_565),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_665),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_642),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_665),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_629),
.B(n_658),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_692),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_698),
.B(n_406),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_746),
.A2(n_398),
.B1(n_400),
.B2(n_402),
.C(n_371),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_669),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_711),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_728),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_669),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_651),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_694),
.B(n_407),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_702),
.B(n_410),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_676),
.B(n_245),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_651),
.B(n_279),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_742),
.Y(n_854)
);

AND2x6_ASAP7_75t_SL g855 ( 
.A(n_676),
.B(n_483),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_751),
.B(n_565),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_768),
.A2(n_565),
.B(n_256),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_671),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_688),
.B(n_280),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_768),
.B(n_588),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_650),
.B(n_290),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_674),
.B(n_299),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_691),
.B(n_300),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_687),
.A2(n_378),
.B1(n_367),
.B2(n_321),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_745),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_671),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_696),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_696),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_687),
.A2(n_338),
.B1(n_361),
.B2(n_305),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_701),
.B(n_361),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_700),
.B(n_293),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_717),
.B(n_562),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_713),
.B(n_390),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_721),
.B(n_581),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_733),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_723),
.B(n_581),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_733),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_703),
.B(n_294),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_727),
.B(n_581),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_728),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_742),
.B(n_304),
.C(n_298),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_755),
.B(n_584),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_769),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_640),
.B(n_390),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_763),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_308),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_758),
.B(n_618),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_769),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_638),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_762),
.B(n_618),
.Y(n_890)
);

AO22x1_ASAP7_75t_L g891 ( 
.A1(n_655),
.A2(n_390),
.B1(n_309),
.B2(n_314),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_640),
.B(n_390),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_719),
.B(n_315),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_638),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_754),
.B(n_618),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_754),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_710),
.B(n_483),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_639),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_686),
.B(n_487),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_754),
.B(n_589),
.Y(n_900)
);

NOR2x1p5_ASAP7_75t_L g901 ( 
.A(n_633),
.B(n_322),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_676),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_763),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_639),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_771),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_672),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_668),
.B(n_323),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_672),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_673),
.A2(n_596),
.B(n_589),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_770),
.B(n_589),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_636),
.B(n_615),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_667),
.A2(n_392),
.B1(n_327),
.B2(n_328),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_686),
.B(n_487),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_756),
.B(n_330),
.Y(n_914)
);

INVxp33_ASAP7_75t_L g915 ( 
.A(n_741),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_636),
.B(n_596),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_636),
.B(n_596),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_690),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_667),
.A2(n_221),
.B1(n_605),
.B2(n_615),
.Y(n_919)
);

INVx8_ASAP7_75t_L g920 ( 
.A(n_667),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_757),
.B(n_615),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_759),
.B(n_332),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_724),
.B(n_605),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_676),
.A2(n_221),
.B1(n_605),
.B2(n_389),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_686),
.B(n_491),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_707),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_724),
.B(n_221),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_724),
.B(n_624),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_857),
.A2(n_678),
.B(n_677),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_847),
.B(n_647),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_776),
.A2(n_675),
.B(n_750),
.C(n_744),
.Y(n_932)
);

CKINVDCx10_ASAP7_75t_R g933 ( 
.A(n_865),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_784),
.B(n_624),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_911),
.A2(n_706),
.B(n_659),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_854),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_916),
.A2(n_706),
.B(n_659),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_773),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_773),
.B(n_635),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_823),
.B(n_647),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_SL g941 ( 
.A1(n_813),
.A2(n_760),
.B(n_646),
.C(n_734),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_842),
.B(n_624),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_917),
.A2(n_860),
.B(n_777),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_847),
.B(n_699),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_910),
.A2(n_706),
.B(n_659),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_783),
.A2(n_764),
.B1(n_743),
.B2(n_647),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_823),
.B(n_635),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_783),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_880),
.B(n_644),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_775),
.A2(n_709),
.B(n_707),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_830),
.A2(n_725),
.B(n_680),
.C(n_695),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_790),
.A2(n_695),
.B1(n_725),
.B2(n_680),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_880),
.B(n_714),
.Y(n_953)
);

AOI22x1_ASAP7_75t_L g954 ( 
.A1(n_896),
.A2(n_686),
.B1(n_659),
.B2(n_704),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_772),
.B(n_624),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_846),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_787),
.Y(n_957)
);

OAI321xp33_ASAP7_75t_L g958 ( 
.A1(n_844),
.A2(n_711),
.A3(n_513),
.B1(n_494),
.B2(n_491),
.C(n_496),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_778),
.A2(n_704),
.B(n_720),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_787),
.A2(n_714),
.B1(n_704),
.B2(n_648),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_805),
.Y(n_961)
);

NOR2xp67_ASAP7_75t_L g962 ( 
.A(n_807),
.B(n_705),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_929),
.A2(n_704),
.B(n_720),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_854),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_786),
.B(n_704),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_823),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_819),
.A2(n_715),
.B(n_709),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_805),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_814),
.B(n_715),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_799),
.B(n_722),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_799),
.B(n_722),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_794),
.A2(n_738),
.B(n_737),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_846),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_809),
.B(n_737),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_828),
.Y(n_975)
);

AOI21x1_ASAP7_75t_L g976 ( 
.A1(n_909),
.A2(n_922),
.B(n_856),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_828),
.Y(n_977)
);

OA22x2_ASAP7_75t_L g978 ( 
.A1(n_899),
.A2(n_766),
.B1(n_705),
.B2(n_352),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_782),
.A2(n_714),
.B1(n_689),
.B2(n_748),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_818),
.B(n_738),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_834),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_853),
.B(n_657),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_834),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_818),
.B(n_740),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_841),
.B(n_334),
.Y(n_985)
);

NAND2x1p5_ASAP7_75t_L g986 ( 
.A(n_823),
.B(n_731),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_817),
.A2(n_729),
.B(n_720),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_821),
.A2(n_729),
.B(n_731),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_871),
.A2(n_740),
.B(n_753),
.C(n_749),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_826),
.A2(n_729),
.B(n_732),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_808),
.B(n_747),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_L g992 ( 
.A(n_820),
.B(n_354),
.C(n_337),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_822),
.B(n_747),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_L g994 ( 
.A(n_804),
.B(n_403),
.C(n_399),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_L g995 ( 
.A(n_802),
.B(n_357),
.C(n_346),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_835),
.A2(n_767),
.B(n_731),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_781),
.A2(n_748),
.B1(n_749),
.B2(n_753),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_801),
.A2(n_837),
.B(n_803),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_SL g999 ( 
.A1(n_873),
.A2(n_514),
.B(n_531),
.C(n_530),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_822),
.B(n_731),
.Y(n_1000)
);

CKINVDCx8_ASAP7_75t_R g1001 ( 
.A(n_865),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_824),
.B(n_732),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_903),
.A2(n_797),
.B(n_793),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_788),
.A2(n_765),
.B(n_645),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_781),
.A2(n_364),
.B1(n_348),
.B2(n_409),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_838),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_L g1007 ( 
.A(n_885),
.B(n_221),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_788),
.A2(n_645),
.B1(n_681),
.B2(n_761),
.Y(n_1008)
);

AOI22x1_ASAP7_75t_L g1009 ( 
.A1(n_896),
.A2(n_767),
.B1(n_732),
.B2(n_761),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_824),
.B(n_732),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_833),
.B(n_732),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_869),
.A2(n_465),
.B(n_461),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_781),
.A2(n_365),
.B1(n_350),
.B2(n_413),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_833),
.B(n_761),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_855),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_885),
.B(n_803),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_808),
.Y(n_1017)
);

AOI22x1_ASAP7_75t_L g1018 ( 
.A1(n_838),
.A2(n_353),
.B1(n_355),
.B2(n_358),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_849),
.B(n_745),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_878),
.A2(n_465),
.B(n_461),
.C(n_375),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_885),
.B(n_812),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_840),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_897),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_836),
.B(n_645),
.Y(n_1024)
);

BUFx4_ASAP7_75t_SL g1025 ( 
.A(n_897),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_836),
.B(n_645),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_779),
.A2(n_499),
.B(n_529),
.C(n_528),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_840),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_800),
.A2(n_765),
.B(n_532),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_858),
.B(n_221),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_858),
.B(n_221),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_901),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_866),
.B(n_351),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_845),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_811),
.A2(n_532),
.B(n_527),
.C(n_521),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_845),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_886),
.A2(n_359),
.B(n_363),
.C(n_383),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_866),
.A2(n_384),
.B1(n_386),
.B2(n_387),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_867),
.B(n_388),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_924),
.A2(n_527),
.B(n_521),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_920),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_895),
.A2(n_517),
.B(n_514),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_900),
.A2(n_890),
.B(n_887),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_848),
.Y(n_1044)
);

INVx6_ASAP7_75t_L g1045 ( 
.A(n_920),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_928),
.A2(n_874),
.B(n_872),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_876),
.A2(n_517),
.B(n_513),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_879),
.A2(n_512),
.B(n_511),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_795),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_806),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_868),
.B(n_396),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_882),
.A2(n_505),
.B(n_499),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_L g1053 ( 
.A(n_792),
.B(n_920),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_920),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_859),
.B(n_497),
.C(n_494),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_883),
.A2(n_211),
.B(n_207),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_888),
.A2(n_206),
.B(n_192),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_825),
.B(n_8),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_888),
.A2(n_176),
.B(n_170),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_839),
.B(n_169),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_867),
.B(n_9),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_852),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_832),
.A2(n_160),
.B(n_156),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_875),
.B(n_9),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_774),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_875),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_877),
.B(n_14),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_843),
.A2(n_152),
.B(n_151),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_877),
.B(n_147),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_905),
.A2(n_145),
.B(n_140),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_899),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_780),
.A2(n_136),
.B(n_134),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_902),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_913),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_815),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_913),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_893),
.B(n_116),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_831),
.B(n_21),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_919),
.B(n_902),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_852),
.B(n_22),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_791),
.A2(n_113),
.B1(n_105),
.B2(n_103),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_829),
.B(n_24),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_889),
.A2(n_97),
.B(n_95),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_864),
.B(n_798),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_889),
.A2(n_88),
.B(n_30),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_905),
.A2(n_29),
.B(n_36),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_789),
.B(n_29),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_798),
.B(n_40),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_918),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_894),
.A2(n_41),
.B(n_43),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_861),
.B(n_41),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_898),
.A2(n_43),
.B(n_44),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_923),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_915),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_862),
.B(n_45),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_904),
.A2(n_48),
.B(n_49),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_904),
.A2(n_49),
.B(n_50),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_906),
.A2(n_53),
.B(n_54),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_908),
.A2(n_59),
.B(n_61),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_918),
.A2(n_61),
.B(n_62),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_925),
.B(n_63),
.Y(n_1101)
);

AOI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_985),
.A2(n_915),
.B(n_827),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_956),
.B(n_852),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1049),
.B(n_796),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_930),
.A2(n_851),
.B(n_921),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_966),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_943),
.A2(n_921),
.B(n_927),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_966),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1003),
.A2(n_852),
.B(n_863),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_998),
.A2(n_870),
.B(n_816),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_937),
.A2(n_892),
.B(n_884),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_985),
.B(n_926),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_936),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_965),
.A2(n_914),
.B(n_891),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1066),
.B(n_1087),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_934),
.A2(n_891),
.B(n_785),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_997),
.A2(n_810),
.A3(n_912),
.B(n_926),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_932),
.A2(n_850),
.B(n_907),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_974),
.A2(n_774),
.B(n_804),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1087),
.B(n_774),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_958),
.A2(n_881),
.B(n_780),
.C(n_792),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_964),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1075),
.B(n_792),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_996),
.A2(n_792),
.B(n_66),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1041),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_967),
.A2(n_792),
.B(n_66),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1084),
.A2(n_792),
.B1(n_69),
.B2(n_70),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1023),
.B(n_65),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_973),
.B(n_65),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1023),
.B(n_71),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1046),
.A2(n_74),
.B(n_75),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_950),
.A2(n_1043),
.B(n_971),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_976),
.A2(n_76),
.B(n_79),
.C(n_81),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_948),
.B(n_84),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1009),
.A2(n_85),
.B(n_959),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_961),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_944),
.A2(n_982),
.B1(n_992),
.B2(n_1051),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_945),
.A2(n_969),
.B(n_970),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_949),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_988),
.A2(n_990),
.B(n_963),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1041),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1094),
.B(n_944),
.Y(n_1142)
);

AOI21xp33_ASAP7_75t_L g1143 ( 
.A1(n_995),
.A2(n_953),
.B(n_1051),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_953),
.B(n_1065),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1033),
.B(n_1039),
.Y(n_1145)
);

NOR2x1_ASAP7_75t_SL g1146 ( 
.A(n_966),
.B(n_1041),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_957),
.B(n_975),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_977),
.B(n_981),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_986),
.A2(n_987),
.B(n_1000),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_955),
.A2(n_972),
.B(n_1053),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1002),
.A2(n_1014),
.B(n_1011),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1079),
.A2(n_941),
.B(n_1021),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1086),
.A2(n_1100),
.B1(n_1080),
.B2(n_1088),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1079),
.A2(n_1010),
.B(n_1004),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_989),
.A2(n_993),
.B(n_980),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1101),
.A2(n_938),
.B(n_1037),
.C(n_1070),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1006),
.B(n_1022),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_984),
.A2(n_1026),
.B(n_1024),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1036),
.B(n_938),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1101),
.A2(n_1020),
.B(n_1082),
.C(n_1061),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1025),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_931),
.B(n_1078),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_968),
.B(n_983),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1025),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_994),
.A2(n_1065),
.B1(n_979),
.B2(n_978),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_966),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_1041),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1028),
.B(n_1034),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1064),
.A2(n_1067),
.B(n_1091),
.C(n_1095),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1030),
.A2(n_1031),
.B(n_942),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_951),
.A2(n_1069),
.B(n_1007),
.Y(n_1171)
);

AOI221x1_ASAP7_75t_L g1172 ( 
.A1(n_994),
.A2(n_1093),
.B1(n_1092),
.B2(n_1090),
.C(n_1099),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1017),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1069),
.A2(n_1077),
.B(n_1029),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_1012),
.A2(n_1072),
.B(n_1085),
.C(n_1044),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_940),
.A2(n_952),
.B(n_1016),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1096),
.A2(n_1098),
.A3(n_1097),
.B(n_1089),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_954),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_947),
.A2(n_1083),
.B(n_1056),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_962),
.B(n_946),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_978),
.A2(n_939),
.B1(n_960),
.B2(n_991),
.Y(n_1181)
);

AND2x6_ASAP7_75t_L g1182 ( 
.A(n_1054),
.B(n_1008),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_947),
.A2(n_1059),
.B(n_1057),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1073),
.B(n_939),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1042),
.A2(n_1040),
.B(n_1035),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1080),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1047),
.A2(n_1048),
.B(n_1052),
.Y(n_1187)
);

BUFx8_ASAP7_75t_L g1188 ( 
.A(n_1032),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1073),
.B(n_1055),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_999),
.Y(n_1190)
);

AND3x1_ASAP7_75t_SL g1191 ( 
.A(n_1050),
.B(n_1071),
.C(n_933),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1073),
.B(n_1058),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1073),
.B(n_1058),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1005),
.A2(n_1013),
.A3(n_1038),
.B(n_1074),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1071),
.B(n_1018),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1074),
.A2(n_1076),
.A3(n_1027),
.B(n_1081),
.Y(n_1196)
);

AND2x2_ASAP7_75t_SL g1197 ( 
.A(n_1019),
.B(n_1060),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1027),
.B(n_1054),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1076),
.A2(n_1045),
.B(n_1054),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1054),
.A2(n_1080),
.B(n_1045),
.C(n_1062),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1045),
.A2(n_1015),
.B(n_1001),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_930),
.A2(n_943),
.B(n_1003),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_956),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_985),
.B(n_776),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_935),
.A2(n_937),
.B(n_996),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_985),
.B(n_776),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1066),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_998),
.A2(n_776),
.B(n_932),
.Y(n_1208)
);

OAI222xp33_ASAP7_75t_L g1209 ( 
.A1(n_1071),
.A2(n_776),
.B1(n_1074),
.B2(n_1076),
.C1(n_1101),
.C2(n_779),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_985),
.B(n_776),
.Y(n_1210)
);

CKINVDCx11_ASAP7_75t_R g1211 ( 
.A(n_1001),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_992),
.B(n_807),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1094),
.B(n_634),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_SL g1214 ( 
.A1(n_1086),
.A2(n_1100),
.B(n_1070),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_930),
.A2(n_943),
.B(n_1003),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_985),
.B(n_776),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1066),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1087),
.A2(n_776),
.B(n_985),
.C(n_627),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_985),
.B(n_776),
.Y(n_1219)
);

OAI22x1_ASAP7_75t_L g1220 ( 
.A1(n_1087),
.A2(n_776),
.B1(n_634),
.B2(n_985),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_998),
.A2(n_776),
.B(n_932),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1023),
.B(n_634),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_1019),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1023),
.B(n_634),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1021),
.A2(n_1003),
.B(n_943),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_935),
.A2(n_937),
.B(n_996),
.Y(n_1226)
);

INVx6_ASAP7_75t_L g1227 ( 
.A(n_1041),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1084),
.A2(n_776),
.B1(n_998),
.B2(n_772),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1023),
.B(n_634),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1087),
.A2(n_776),
.B(n_985),
.C(n_627),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_933),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_930),
.A2(n_943),
.B(n_1003),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_958),
.A2(n_776),
.B1(n_1100),
.B2(n_1086),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_935),
.A2(n_937),
.B(n_996),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_966),
.B(n_1041),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_985),
.A2(n_776),
.B1(n_625),
.B2(n_1087),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_966),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_930),
.A2(n_943),
.B(n_1003),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_998),
.A2(n_776),
.B(n_932),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_935),
.A2(n_937),
.B(n_996),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_998),
.A2(n_776),
.B(n_932),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1021),
.A2(n_1003),
.B(n_943),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_935),
.A2(n_937),
.B(n_996),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1087),
.A2(n_776),
.B(n_985),
.C(n_627),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1049),
.B(n_776),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_985),
.B(n_776),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1087),
.A2(n_776),
.B(n_985),
.C(n_627),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_967),
.A2(n_930),
.B(n_943),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_956),
.Y(n_1249)
);

OAI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_985),
.A2(n_776),
.B(n_617),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_985),
.B(n_776),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1200),
.B(n_1103),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1207),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1217),
.Y(n_1254)
);

OR2x6_ASAP7_75t_L g1255 ( 
.A(n_1161),
.B(n_1164),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1136),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1236),
.A2(n_1216),
.B1(n_1246),
.B2(n_1210),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1148),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1213),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1137),
.B(n_1180),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1113),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1219),
.B(n_1251),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1103),
.B(n_1203),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1249),
.B(n_1201),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1157),
.Y(n_1266)
);

CKINVDCx8_ASAP7_75t_R g1267 ( 
.A(n_1231),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1139),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1152),
.A2(n_1215),
.B(n_1202),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1245),
.A2(n_1236),
.B1(n_1197),
.B2(n_1223),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_L g1271 ( 
.A(n_1125),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1167),
.B(n_1106),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1173),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1250),
.A2(n_1230),
.B1(n_1244),
.B2(n_1247),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1184),
.B(n_1162),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1222),
.B(n_1224),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1122),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1211),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1218),
.B(n_1112),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1125),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1129),
.Y(n_1281)
);

OR2x6_ASAP7_75t_SL g1282 ( 
.A(n_1145),
.B(n_1120),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1229),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1192),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1115),
.B(n_1208),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1125),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1220),
.A2(n_1165),
.B1(n_1233),
.B2(n_1142),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1147),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1221),
.A2(n_1239),
.B(n_1241),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1209),
.A2(n_1233),
.B(n_1153),
.C(n_1102),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1163),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1186),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1144),
.B(n_1212),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1228),
.B(n_1193),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1166),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1168),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1143),
.B(n_1181),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1128),
.B(n_1130),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1188),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_1159),
.Y(n_1301)
);

BUFx10_ASAP7_75t_L g1302 ( 
.A(n_1227),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1167),
.B(n_1141),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1141),
.Y(n_1304)
);

AOI21xp33_ASAP7_75t_L g1305 ( 
.A1(n_1153),
.A2(n_1214),
.B(n_1118),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1152),
.A2(n_1154),
.B(n_1110),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1209),
.A2(n_1160),
.B(n_1156),
.C(n_1127),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1188),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1166),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1141),
.B(n_1146),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1134),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1227),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1189),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1195),
.B(n_1119),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1235),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1191),
.A2(n_1198),
.B1(n_1235),
.B2(n_1227),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1232),
.A2(n_1132),
.B(n_1238),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1108),
.B(n_1199),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1237),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1237),
.B(n_1182),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1182),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1238),
.A2(n_1248),
.B(n_1138),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1182),
.B(n_1121),
.Y(n_1323)
);

BUFx2_ASAP7_75t_SL g1324 ( 
.A(n_1182),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1150),
.A2(n_1178),
.B(n_1109),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1131),
.A2(n_1123),
.B(n_1110),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1182),
.B(n_1172),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1109),
.A2(n_1178),
.B(n_1176),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1176),
.B(n_1126),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1116),
.B(n_1114),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1174),
.A2(n_1155),
.B(n_1105),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1194),
.B(n_1171),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1114),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1190),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1135),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1107),
.A2(n_1105),
.B(n_1170),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1124),
.B(n_1174),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1158),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1185),
.A2(n_1175),
.B(n_1151),
.C(n_1133),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1171),
.A2(n_1183),
.B1(n_1179),
.B2(n_1187),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_1242),
.B1(n_1225),
.B2(n_1194),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1149),
.B(n_1111),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1140),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1205),
.B(n_1243),
.Y(n_1345)
);

AND2x2_ASAP7_75t_SL g1346 ( 
.A(n_1196),
.B(n_1117),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1196),
.B(n_1117),
.C(n_1226),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1234),
.B(n_1240),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1211),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1200),
.B(n_1045),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1125),
.Y(n_1351)
);

AOI21xp33_ASAP7_75t_L g1352 ( 
.A1(n_1204),
.A2(n_1210),
.B(n_1206),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1207),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1207),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1204),
.A2(n_776),
.B1(n_764),
.B2(n_1206),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1207),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_L g1357 ( 
.A(n_1125),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1207),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1207),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1207),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1218),
.A2(n_1244),
.B(n_1247),
.C(n_1230),
.Y(n_1361)
);

BUFx4_ASAP7_75t_SL g1362 ( 
.A(n_1231),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1236),
.A2(n_1204),
.B1(n_1210),
.B2(n_1206),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1113),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1113),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1200),
.B(n_1103),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1204),
.B(n_776),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_SL g1371 ( 
.A1(n_1208),
.A2(n_776),
.B(n_1087),
.C(n_627),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1222),
.B(n_634),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1222),
.B(n_634),
.Y(n_1373)
);

AND2x4_ASAP7_75t_SL g1374 ( 
.A(n_1167),
.B(n_642),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1213),
.B(n_807),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_R g1376 ( 
.A(n_1211),
.B(n_657),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1204),
.A2(n_776),
.B1(n_1210),
.B2(n_1206),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1218),
.A2(n_1244),
.B(n_1247),
.C(n_1230),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1207),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1113),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1213),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1213),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1113),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1113),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1113),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1125),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1200),
.B(n_1103),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1207),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1207),
.Y(n_1390)
);

INVx3_ASAP7_75t_SL g1391 ( 
.A(n_1231),
.Y(n_1391)
);

INVx3_ASAP7_75t_SL g1392 ( 
.A(n_1231),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1113),
.Y(n_1393)
);

NOR2x1_ASAP7_75t_SL g1394 ( 
.A(n_1125),
.B(n_966),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1125),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1204),
.B(n_1206),
.Y(n_1396)
);

AO22x1_ASAP7_75t_L g1397 ( 
.A1(n_1245),
.A2(n_776),
.B1(n_1206),
.B2(n_1204),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1125),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1343),
.Y(n_1399)
);

BUFx2_ASAP7_75t_SL g1400 ( 
.A(n_1387),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1376),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1369),
.A2(n_1364),
.B1(n_1355),
.B2(n_1257),
.Y(n_1402)
);

BUFx8_ASAP7_75t_L g1403 ( 
.A(n_1300),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1387),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1314),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1356),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1333),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1296),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1333),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1349),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1263),
.B(n_1377),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1358),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1252),
.B(n_1368),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1321),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1267),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1259),
.B(n_1363),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1323),
.A2(n_1274),
.B1(n_1370),
.B2(n_1367),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1264),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1252),
.B(n_1368),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1359),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1360),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1364),
.A2(n_1261),
.B1(n_1287),
.B2(n_1270),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1320),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1284),
.B(n_1313),
.Y(n_1424)
);

CKINVDCx6p67_ASAP7_75t_R g1425 ( 
.A(n_1391),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1365),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1388),
.B(n_1320),
.Y(n_1428)
);

INVx11_ASAP7_75t_L g1429 ( 
.A(n_1362),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1323),
.A2(n_1338),
.B1(n_1299),
.B2(n_1324),
.Y(n_1430)
);

AO21x1_ASAP7_75t_L g1431 ( 
.A1(n_1290),
.A2(n_1378),
.B(n_1361),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1389),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1253),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1254),
.Y(n_1434)
);

CKINVDCx11_ASAP7_75t_R g1435 ( 
.A(n_1392),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1260),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1298),
.A2(n_1289),
.B1(n_1352),
.B2(n_1305),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1382),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1289),
.B(n_1285),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1353),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1352),
.A2(n_1305),
.B1(n_1370),
.B2(n_1367),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1308),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1259),
.A2(n_1396),
.B1(n_1363),
.B2(n_1379),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1382),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1284),
.B(n_1346),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1279),
.B(n_1275),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1309),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1339),
.A2(n_1322),
.B(n_1317),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1318),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1278),
.Y(n_1450)
);

BUFx10_ASAP7_75t_L g1451 ( 
.A(n_1374),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1383),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1379),
.A2(n_1396),
.B1(n_1294),
.B2(n_1327),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1334),
.A2(n_1282),
.B1(n_1383),
.B2(n_1311),
.Y(n_1454)
);

NOR2x1_ASAP7_75t_L g1455 ( 
.A(n_1375),
.B(n_1350),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1279),
.B(n_1275),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1390),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1397),
.A2(n_1316),
.B1(n_1293),
.B2(n_1388),
.Y(n_1458)
);

NAND2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1318),
.B(n_1327),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1372),
.B(n_1373),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1258),
.B(n_1266),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1256),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1387),
.Y(n_1463)
);

BUFx2_ASAP7_75t_SL g1464 ( 
.A(n_1387),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1291),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1297),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1330),
.A2(n_1276),
.B1(n_1273),
.B2(n_1283),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1288),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1350),
.B(n_1265),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1347),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1285),
.B(n_1295),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1307),
.B(n_1350),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1262),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1269),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1335),
.B(n_1332),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1366),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1335),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1385),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1292),
.A2(n_1384),
.B1(n_1381),
.B2(n_1386),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1295),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1265),
.A2(n_1281),
.B1(n_1393),
.B2(n_1306),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1335),
.B(n_1332),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1301),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1268),
.A2(n_1301),
.B1(n_1277),
.B2(n_1255),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1341),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1328),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1255),
.A2(n_1326),
.B1(n_1264),
.B2(n_1331),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1328),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1310),
.B(n_1303),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1255),
.A2(n_1329),
.B1(n_1306),
.B2(n_1337),
.Y(n_1490)
);

CKINVDCx9p33_ASAP7_75t_R g1491 ( 
.A(n_1342),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1302),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1348),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1329),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1302),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1329),
.A2(n_1337),
.B1(n_1319),
.B2(n_1344),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1271),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1312),
.A2(n_1315),
.B1(n_1272),
.B2(n_1310),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1271),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1337),
.A2(n_1319),
.B1(n_1303),
.B2(n_1336),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1336),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1280),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1319),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1340),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1371),
.A2(n_1345),
.B(n_1394),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1280),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1286),
.A2(n_1304),
.B1(n_1351),
.B2(n_1395),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1286),
.A2(n_1304),
.B1(n_1351),
.B2(n_1395),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1351),
.A2(n_1395),
.B1(n_1398),
.B2(n_1357),
.Y(n_1509)
);

BUFx12f_ASAP7_75t_L g1510 ( 
.A(n_1398),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1272),
.A2(n_1357),
.B(n_1398),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1339),
.A2(n_1325),
.B(n_1322),
.Y(n_1512)
);

CKINVDCx11_ASAP7_75t_R g1513 ( 
.A(n_1267),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1387),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1369),
.A2(n_776),
.B(n_1218),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1369),
.A2(n_776),
.B1(n_1236),
.B2(n_1206),
.Y(n_1516)
);

INVx6_ASAP7_75t_L g1517 ( 
.A(n_1387),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1321),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1354),
.Y(n_1519)
);

AOI21xp33_ASAP7_75t_L g1520 ( 
.A1(n_1371),
.A2(n_776),
.B(n_1204),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_SL g1521 ( 
.A(n_1308),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1369),
.B(n_1263),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1354),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1260),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1321),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1354),
.Y(n_1526)
);

CKINVDCx8_ASAP7_75t_R g1527 ( 
.A(n_1349),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1324),
.B(n_1290),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1377),
.A2(n_1206),
.B1(n_1210),
.B2(n_1204),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1264),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1270),
.A2(n_776),
.B1(n_1206),
.B2(n_1204),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1354),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1376),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1354),
.Y(n_1534)
);

NAND2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1318),
.B(n_1321),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1321),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1369),
.B(n_1263),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1387),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1369),
.A2(n_776),
.B1(n_1236),
.B2(n_1206),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1369),
.A2(n_776),
.B1(n_1245),
.B2(n_1206),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1369),
.B(n_1263),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1264),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1408),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1411),
.B(n_1443),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1475),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1399),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1445),
.B(n_1405),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1515),
.A2(n_1539),
.B(n_1516),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1436),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1459),
.B(n_1446),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1540),
.B(n_1522),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1492),
.Y(n_1552)
);

BUFx5_ASAP7_75t_L g1553 ( 
.A(n_1501),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_R g1554 ( 
.A(n_1513),
.B(n_1435),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1407),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1408),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1459),
.Y(n_1557)
);

OR2x6_ASAP7_75t_L g1558 ( 
.A(n_1494),
.B(n_1472),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_SL g1559 ( 
.A(n_1527),
.B(n_1415),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1433),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1459),
.B(n_1446),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1438),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1470),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1470),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1444),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1434),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1456),
.B(n_1471),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1452),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1429),
.Y(n_1569)
);

AO21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1422),
.A2(n_1485),
.B(n_1504),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1439),
.B(n_1501),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1524),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1493),
.B(n_1504),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1437),
.B(n_1472),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1531),
.A2(n_1520),
.B(n_1529),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1472),
.B(n_1480),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1472),
.B(n_1480),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1528),
.A2(n_1541),
.B1(n_1537),
.B2(n_1483),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1482),
.B(n_1528),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1447),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1424),
.B(n_1409),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1402),
.A2(n_1441),
.B(n_1487),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1447),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1528),
.B(n_1469),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1449),
.B(n_1469),
.Y(n_1585)
);

AO31x2_ASAP7_75t_L g1586 ( 
.A1(n_1486),
.A2(n_1488),
.A3(n_1431),
.B(n_1474),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1490),
.B(n_1440),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1460),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1462),
.B(n_1483),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1476),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1465),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1465),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1528),
.B(n_1461),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1477),
.B(n_1413),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1458),
.B(n_1473),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1457),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1517),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1453),
.B(n_1448),
.Y(n_1598)
);

BUFx4f_ASAP7_75t_SL g1599 ( 
.A(n_1415),
.Y(n_1599)
);

NAND2x1_ASAP7_75t_L g1600 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1448),
.B(n_1467),
.Y(n_1601)
);

BUFx2_ASAP7_75t_SL g1602 ( 
.A(n_1492),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1512),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1512),
.Y(n_1604)
);

AO21x2_ASAP7_75t_L g1605 ( 
.A1(n_1505),
.A2(n_1431),
.B(n_1417),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1512),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1406),
.B(n_1412),
.Y(n_1607)
);

AO21x2_ASAP7_75t_L g1608 ( 
.A1(n_1505),
.A2(n_1454),
.B(n_1466),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1412),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1420),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1535),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1416),
.B(n_1468),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1535),
.A2(n_1511),
.B(n_1423),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1421),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1426),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1432),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1432),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1519),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1519),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1523),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1523),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1413),
.B(n_1419),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1484),
.B(n_1526),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1532),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1546),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1558),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1599),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1567),
.B(n_1419),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1544),
.B(n_1430),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1579),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1580),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1583),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1558),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1601),
.B(n_1505),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1548),
.A2(n_1419),
.B1(n_1413),
.B2(n_1481),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1569),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1534),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1549),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1558),
.Y(n_1639)
);

INVx5_ASAP7_75t_L g1640 ( 
.A(n_1579),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1550),
.B(n_1428),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1581),
.B(n_1534),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1601),
.B(n_1598),
.Y(n_1643)
);

NAND2x1_ASAP7_75t_L g1644 ( 
.A(n_1584),
.B(n_1517),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1582),
.A2(n_1455),
.B1(n_1423),
.B2(n_1478),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1598),
.B(n_1479),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1602),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1551),
.B(n_1473),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1565),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1543),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1558),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1568),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1571),
.B(n_1536),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1561),
.B(n_1536),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1558),
.B(n_1584),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1602),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1586),
.B(n_1518),
.Y(n_1657)
);

NOR2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1414),
.Y(n_1658)
);

AND2x4_ASAP7_75t_SL g1659 ( 
.A(n_1622),
.B(n_1451),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1547),
.B(n_1576),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1584),
.B(n_1525),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1577),
.B(n_1525),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1572),
.B(n_1506),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_L g1665 ( 
.A(n_1611),
.B(n_1503),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1608),
.B(n_1400),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1556),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1563),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1563),
.Y(n_1669)
);

OA21x2_ASAP7_75t_L g1670 ( 
.A1(n_1603),
.A2(n_1511),
.B(n_1491),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1593),
.B(n_1489),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1575),
.A2(n_1498),
.B(n_1514),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1587),
.B(n_1489),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1587),
.B(n_1502),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1588),
.B(n_1478),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1564),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1584),
.B(n_1542),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1608),
.B(n_1400),
.Y(n_1678)
);

INVxp67_ASAP7_75t_SL g1679 ( 
.A(n_1555),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1595),
.A2(n_1509),
.B(n_1527),
.C(n_1442),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1586),
.B(n_1530),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1645),
.A2(n_1584),
.B1(n_1600),
.B2(n_1579),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1638),
.B(n_1562),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1625),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1660),
.B(n_1574),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1634),
.A2(n_1606),
.B(n_1604),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1634),
.A2(n_1606),
.B(n_1604),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1652),
.B(n_1556),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1649),
.B(n_1591),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1629),
.B(n_1578),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1672),
.B(n_1578),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1646),
.B(n_1623),
.C(n_1574),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1635),
.A2(n_1658),
.B1(n_1680),
.B2(n_1656),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1630),
.B(n_1622),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1646),
.B(n_1623),
.C(n_1612),
.Y(n_1695)
);

OR2x2_ASAP7_75t_SL g1696 ( 
.A(n_1631),
.B(n_1554),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1625),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1590),
.C(n_1573),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1666),
.B(n_1573),
.C(n_1614),
.Y(n_1700)
);

NOR3xp33_ASAP7_75t_L g1701 ( 
.A(n_1648),
.B(n_1554),
.C(n_1611),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1658),
.A2(n_1579),
.B1(n_1552),
.B2(n_1622),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1647),
.B(n_1674),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1664),
.B(n_1596),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1679),
.B(n_1596),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1628),
.B(n_1589),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1628),
.B(n_1589),
.Y(n_1707)
);

OAI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1644),
.A2(n_1579),
.B1(n_1559),
.B2(n_1552),
.Y(n_1708)
);

OA211x2_ASAP7_75t_L g1709 ( 
.A1(n_1644),
.A2(n_1608),
.B(n_1508),
.C(n_1507),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1667),
.B(n_1619),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1675),
.A2(n_1622),
.B1(n_1418),
.B2(n_1585),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1627),
.A2(n_1570),
.B1(n_1605),
.B2(n_1427),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1641),
.B(n_1585),
.Y(n_1713)
);

OAI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1678),
.A2(n_1495),
.B1(n_1450),
.B2(n_1611),
.C(n_1597),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1630),
.B(n_1585),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1643),
.B(n_1586),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1643),
.A2(n_1605),
.B1(n_1621),
.B2(n_1620),
.C(n_1618),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1673),
.A2(n_1605),
.B1(n_1621),
.B2(n_1620),
.C(n_1618),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1678),
.B(n_1624),
.C(n_1615),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1681),
.B(n_1624),
.C(n_1609),
.Y(n_1720)
);

OAI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1681),
.A2(n_1450),
.B1(n_1597),
.B2(n_1497),
.C(n_1499),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1665),
.A2(n_1613),
.B(n_1594),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_L g1723 ( 
.A(n_1670),
.B(n_1615),
.C(n_1609),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1673),
.B(n_1671),
.Y(n_1724)
);

OAI221xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1657),
.A2(n_1425),
.B1(n_1557),
.B2(n_1497),
.C(n_1499),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1671),
.B(n_1594),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1630),
.B(n_1553),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1670),
.B(n_1617),
.C(n_1616),
.Y(n_1728)
);

NAND4xp25_ASAP7_75t_L g1729 ( 
.A(n_1637),
.B(n_1607),
.C(n_1617),
.D(n_1616),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1642),
.B(n_1560),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1670),
.B(n_1610),
.C(n_1607),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1630),
.B(n_1640),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1655),
.A2(n_1403),
.B(n_1545),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1630),
.B(n_1553),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1653),
.B(n_1566),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_SL g1736 ( 
.A1(n_1655),
.A2(n_1659),
.B(n_1662),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1698),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1698),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1716),
.B(n_1657),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1686),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1684),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1705),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1686),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1685),
.B(n_1655),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1710),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1669),
.C(n_1668),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1735),
.Y(n_1747)
);

INVx4_ASAP7_75t_R g1748 ( 
.A(n_1696),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1697),
.B(n_1669),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1690),
.A2(n_1677),
.B1(n_1662),
.B2(n_1651),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1686),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1687),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1687),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1687),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1720),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1723),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1719),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1722),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1715),
.B(n_1662),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1688),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1683),
.B(n_1689),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1730),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1731),
.B(n_1676),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1704),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1728),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1662),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1732),
.B(n_1626),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1690),
.B(n_1654),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1700),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1732),
.B(n_1633),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1724),
.B(n_1633),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1727),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1724),
.B(n_1639),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1694),
.B(n_1651),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1694),
.B(n_1663),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1699),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1695),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1737),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1739),
.B(n_1692),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1737),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1706),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1740),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1748),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1763),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1775),
.B(n_1736),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1738),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1777),
.B(n_1707),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1775),
.B(n_1703),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1738),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1740),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1777),
.B(n_1703),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1769),
.B(n_1756),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1769),
.B(n_1729),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1744),
.B(n_1726),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1741),
.Y(n_1798)
);

OAI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1746),
.A2(n_1691),
.B(n_1712),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1776),
.B(n_1713),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1741),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1776),
.B(n_1718),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1760),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_SL g1804 ( 
.A(n_1758),
.B(n_1714),
.C(n_1701),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1744),
.B(n_1726),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1763),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1767),
.B(n_1759),
.Y(n_1807)
);

NOR2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1746),
.B(n_1425),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1756),
.B(n_1650),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1757),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1758),
.B(n_1708),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1756),
.B(n_1650),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1748),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1750),
.A2(n_1733),
.B(n_1693),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1745),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1751),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1751),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1742),
.B(n_1654),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1774),
.B(n_1727),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_1734),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1743),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1743),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1759),
.B(n_1734),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1742),
.B(n_1661),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1752),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1759),
.B(n_1702),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1764),
.B(n_1661),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1757),
.Y(n_1828)
);

NOR2xp67_ASAP7_75t_L g1829 ( 
.A(n_1765),
.B(n_1721),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1759),
.B(n_1677),
.Y(n_1830)
);

INVx3_ASAP7_75t_R g1831 ( 
.A(n_1765),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1798),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1799),
.A2(n_1682),
.B1(n_1709),
.B2(n_1755),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1798),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1802),
.B(n_1755),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1794),
.B(n_1765),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1803),
.B(n_1815),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1783),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1807),
.B(n_1767),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1799),
.A2(n_1770),
.B(n_1767),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1801),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1793),
.B(n_1768),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1810),
.B(n_1828),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1794),
.B(n_1772),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1807),
.B(n_1767),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1807),
.B(n_1770),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1795),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1795),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1783),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1784),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1807),
.B(n_1770),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1783),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1804),
.A2(n_1761),
.B1(n_1764),
.B2(n_1762),
.C(n_1747),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1784),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1801),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1829),
.B(n_1762),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1811),
.B(n_1712),
.C(n_1717),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1788),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1816),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1788),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1813),
.B(n_1725),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1813),
.B(n_1403),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1780),
.B(n_1772),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1779),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1778),
.B(n_1766),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1780),
.B(n_1772),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1788),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1806),
.B(n_1749),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1816),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1786),
.B(n_1766),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1817),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1806),
.B(n_1785),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_L g1874 ( 
.A(n_1808),
.B(n_1636),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1778),
.B(n_1766),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1789),
.B(n_1749),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1817),
.Y(n_1877)
);

INVxp67_ASAP7_75t_L g1878 ( 
.A(n_1809),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1825),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1792),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1808),
.B(n_1814),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1779),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1809),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1812),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1792),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1850),
.B(n_1823),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1835),
.B(n_1790),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1850),
.B(n_1854),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1861),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1866),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1866),
.B(n_1823),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1859),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1859),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1862),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1870),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1837),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1836),
.B(n_1789),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1883),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1870),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1881),
.B(n_1403),
.Y(n_1900)
);

NOR2x1_ASAP7_75t_L g1901 ( 
.A(n_1881),
.B(n_1812),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1871),
.B(n_1786),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1843),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1875),
.B(n_1819),
.Y(n_1904)
);

CKINVDCx16_ASAP7_75t_R g1905 ( 
.A(n_1881),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1884),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1881),
.A2(n_1814),
.B1(n_1826),
.B2(n_1766),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1836),
.B(n_1782),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1876),
.B(n_1782),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1863),
.B(n_1790),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1857),
.A2(n_1826),
.B1(n_1820),
.B2(n_1819),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1853),
.B(n_1820),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1872),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1874),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1876),
.B(n_1827),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1873),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1856),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1872),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1875),
.B(n_1830),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1864),
.B(n_1824),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1846),
.B(n_1830),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1877),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1846),
.B(n_1796),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1851),
.B(n_1796),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1838),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1905),
.B(n_1833),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1898),
.B(n_1847),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1889),
.A2(n_1840),
.B1(n_1848),
.B2(n_1878),
.Y(n_1928)
);

AOI322xp5_ASAP7_75t_SL g1929 ( 
.A1(n_1886),
.A2(n_1831),
.A3(n_1851),
.B1(n_1845),
.B2(n_1839),
.C1(n_1771),
.C2(n_1773),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1916),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1901),
.A2(n_1873),
.B(n_1867),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1888),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1912),
.A2(n_1842),
.B(n_1864),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1906),
.B(n_1867),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1892),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1888),
.B(n_1839),
.Y(n_1936)
);

AOI21xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1905),
.A2(n_1569),
.B(n_1831),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1892),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1914),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1890),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1893),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1923),
.B(n_1845),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1907),
.A2(n_1832),
.B1(n_1841),
.B2(n_1834),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1893),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1895),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1894),
.B(n_1844),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1902),
.A2(n_1855),
.B1(n_1869),
.B2(n_1865),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1894),
.B(n_1844),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1895),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1923),
.B(n_1869),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1917),
.B(n_1805),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1924),
.B(n_1882),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1896),
.B(n_1911),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1886),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1932),
.B(n_1887),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1939),
.B(n_1904),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1928),
.A2(n_1902),
.B1(n_1890),
.B2(n_1910),
.Y(n_1957)
);

OAI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1929),
.A2(n_1909),
.B1(n_1902),
.B2(n_1908),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1936),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_SL g1960 ( 
.A(n_1932),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1940),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1936),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1935),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1954),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1937),
.B(n_1900),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1942),
.B(n_1904),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1936),
.B(n_1897),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1954),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1926),
.A2(n_1903),
.B(n_1897),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_SL g1970 ( 
.A(n_1926),
.B(n_1401),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1952),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1938),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1930),
.B(n_1891),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1946),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1946),
.B(n_1891),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1934),
.B(n_1909),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_L g1977 ( 
.A(n_1953),
.B(n_1401),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1952),
.Y(n_1978)
);

O2A1O1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1958),
.A2(n_1931),
.B(n_1948),
.C(n_1927),
.Y(n_1979)
);

A2O1A1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1970),
.A2(n_1969),
.B(n_1974),
.C(n_1933),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_L g1981 ( 
.A(n_1970),
.B(n_1948),
.C(n_1943),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1956),
.B(n_1947),
.Y(n_1982)
);

NAND3xp33_ASAP7_75t_L g1983 ( 
.A(n_1977),
.B(n_1944),
.C(n_1941),
.Y(n_1983)
);

AOI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1957),
.A2(n_1945),
.B(n_1949),
.C(n_1951),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1956),
.A2(n_1942),
.B(n_1950),
.Y(n_1985)
);

NOR3xp33_ASAP7_75t_L g1986 ( 
.A(n_1977),
.B(n_1950),
.C(n_1913),
.Y(n_1986)
);

AOI222xp33_ASAP7_75t_L g1987 ( 
.A1(n_1967),
.A2(n_1922),
.B1(n_1913),
.B2(n_1918),
.C1(n_1899),
.C2(n_1919),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_SL g1988 ( 
.A(n_1959),
.B(n_1410),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1964),
.Y(n_1989)
);

OAI21xp33_ASAP7_75t_L g1990 ( 
.A1(n_1975),
.A2(n_1919),
.B(n_1921),
.Y(n_1990)
);

NAND5xp2_ASAP7_75t_L g1991 ( 
.A(n_1973),
.B(n_1966),
.C(n_1961),
.D(n_1963),
.E(n_1972),
.Y(n_1991)
);

AOI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1962),
.A2(n_1899),
.B1(n_1922),
.B2(n_1918),
.C(n_1925),
.Y(n_1992)
);

AOI21x1_ASAP7_75t_L g1993 ( 
.A1(n_1968),
.A2(n_1925),
.B(n_1879),
.Y(n_1993)
);

NAND4xp25_ASAP7_75t_L g1994 ( 
.A(n_1991),
.B(n_1965),
.C(n_1976),
.D(n_1968),
.Y(n_1994)
);

NOR3xp33_ASAP7_75t_L g1995 ( 
.A(n_1980),
.B(n_1976),
.C(n_1955),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1989),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1979),
.B(n_1955),
.C(n_1971),
.Y(n_1997)
);

NOR2x1_ASAP7_75t_L g1998 ( 
.A(n_1981),
.B(n_1533),
.Y(n_1998)
);

AOI211xp5_ASAP7_75t_L g1999 ( 
.A1(n_1982),
.A2(n_1978),
.B(n_1971),
.C(n_1966),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1983),
.B(n_1533),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1988),
.A2(n_1978),
.B1(n_1960),
.B2(n_1921),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_SL g2002 ( 
.A(n_1986),
.B(n_1908),
.C(n_1920),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1993),
.Y(n_2003)
);

NOR3x1_ASAP7_75t_L g2004 ( 
.A(n_1984),
.B(n_1920),
.C(n_1915),
.Y(n_2004)
);

AOI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_1985),
.A2(n_1924),
.B(n_1915),
.C(n_1877),
.Y(n_2005)
);

NOR2x1_ASAP7_75t_L g2006 ( 
.A(n_1990),
.B(n_1429),
.Y(n_2006)
);

OAI211xp5_ASAP7_75t_L g2007 ( 
.A1(n_1994),
.A2(n_1987),
.B(n_1992),
.C(n_1879),
.Y(n_2007)
);

NAND4xp25_ASAP7_75t_SL g2008 ( 
.A(n_2001),
.B(n_1885),
.C(n_1852),
.D(n_1838),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_2003),
.Y(n_2009)
);

NAND4xp25_ASAP7_75t_L g2010 ( 
.A(n_1998),
.B(n_1521),
.C(n_1849),
.D(n_1860),
.Y(n_2010)
);

AOI221x1_ASAP7_75t_L g2011 ( 
.A1(n_1997),
.A2(n_1996),
.B1(n_1995),
.B2(n_2002),
.C(n_1999),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_2000),
.B(n_2006),
.Y(n_2012)
);

NAND3xp33_ASAP7_75t_L g2013 ( 
.A(n_2005),
.B(n_1852),
.C(n_1849),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_2009),
.Y(n_2014)
);

NOR3xp33_ASAP7_75t_L g2015 ( 
.A(n_2012),
.B(n_2004),
.C(n_1410),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2013),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_2007),
.B(n_1858),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2011),
.Y(n_2018)
);

AO22x1_ASAP7_75t_L g2019 ( 
.A1(n_2008),
.A2(n_2010),
.B1(n_1521),
.B2(n_1880),
.Y(n_2019)
);

INVxp67_ASAP7_75t_L g2020 ( 
.A(n_2012),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_2011),
.A2(n_1860),
.B(n_1858),
.Y(n_2021)
);

OAI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_2018),
.A2(n_1885),
.B1(n_1880),
.B2(n_1868),
.C(n_1825),
.Y(n_2022)
);

AND4x1_ASAP7_75t_L g2023 ( 
.A(n_2015),
.B(n_1521),
.C(n_1451),
.D(n_1427),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2020),
.A2(n_1868),
.B1(n_1797),
.B2(n_1822),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2014),
.B(n_1818),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_SL g2026 ( 
.A(n_2016),
.B(n_1451),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_2021),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_2017),
.Y(n_2028)
);

OA22x2_ASAP7_75t_L g2029 ( 
.A1(n_2028),
.A2(n_2021),
.B1(n_2019),
.B2(n_1792),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_2023),
.Y(n_2030)
);

NOR3xp33_ASAP7_75t_L g2031 ( 
.A(n_2027),
.B(n_1514),
.C(n_1711),
.Y(n_2031)
);

AOI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_2026),
.A2(n_1822),
.B1(n_1797),
.B2(n_1821),
.Y(n_2032)
);

AO22x2_ASAP7_75t_L g2033 ( 
.A1(n_2030),
.A2(n_2025),
.B1(n_2022),
.B2(n_2024),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2029),
.Y(n_2034)
);

A2O1A1Ixp33_ASAP7_75t_L g2035 ( 
.A1(n_2034),
.A2(n_2031),
.B(n_2032),
.C(n_1822),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2035),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_2035),
.A2(n_2033),
.B1(n_1797),
.B2(n_1821),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_2036),
.A2(n_1821),
.B(n_1787),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2037),
.B(n_1781),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2039),
.A2(n_1787),
.B(n_1781),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_2040),
.A2(n_2038),
.B(n_1791),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_R g2042 ( 
.A1(n_2041),
.A2(n_1791),
.B1(n_1753),
.B2(n_1752),
.Y(n_2042)
);

OAI221xp5_ASAP7_75t_R g2043 ( 
.A1(n_2042),
.A2(n_1510),
.B1(n_1464),
.B2(n_1753),
.C(n_1754),
.Y(n_2043)
);

AOI211xp5_ASAP7_75t_L g2044 ( 
.A1(n_2043),
.A2(n_1463),
.B(n_1404),
.C(n_1538),
.Y(n_2044)
);


endmodule