module fake_jpeg_4995_n_16 (n_3, n_2, n_1, n_0, n_4, n_16);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_16;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_0),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_2),
.B(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_2),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_0),
.Y(n_9)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_11),
.B(n_7),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g10 ( 
.A1(n_6),
.A2(n_1),
.B(n_2),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_12),
.C(n_5),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

AOI322xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_14),
.A3(n_5),
.B1(n_4),
.B2(n_3),
.C1(n_1),
.C2(n_8),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_8),
.B1(n_4),
.B2(n_3),
.Y(n_16)
);


endmodule