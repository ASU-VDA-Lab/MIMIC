module fake_netlist_6_1_n_1848 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1848);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1848;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_100),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_35),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_60),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_15),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_99),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_51),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_66),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_147),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_81),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_6),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_23),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_86),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_164),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_26),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_105),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_155),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_19),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_36),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_98),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_124),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_9),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_82),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_109),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_50),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_102),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_55),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_36),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_120),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_110),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_3),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_13),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_143),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_41),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_42),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_76),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_152),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_72),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_114),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_145),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_56),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_23),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_106),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_61),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_113),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_107),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_103),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_131),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_51),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_62),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_166),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_77),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_168),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_169),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_156),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_45),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_58),
.Y(n_273)
);

BUFx2_ASAP7_75t_R g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_29),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_96),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_157),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_12),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_95),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_118),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_180),
.Y(n_283)
);

BUFx2_ASAP7_75t_SL g284 ( 
.A(n_150),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_93),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_126),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_75),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_160),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_18),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_44),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_174),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_141),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_178),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_116),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_78),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_14),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_123),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_38),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_64),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_63),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_133),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_183),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_35),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_173),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_52),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_88),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_30),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_13),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_5),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_44),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_71),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_162),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_39),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_16),
.Y(n_317)
);

BUFx2_ASAP7_75t_SL g318 ( 
.A(n_1),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_8),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_53),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_129),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_54),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_4),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_153),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_127),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_84),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_40),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_20),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_22),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_90),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_53),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_41),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_0),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_20),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_37),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_31),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_33),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_119),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_137),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_80),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_144),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_167),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_111),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_135),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_56),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_28),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_67),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_104),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_159),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_50),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_4),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_108),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_140),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_70),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_179),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_32),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_151),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_33),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_18),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_55),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_10),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_59),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_122),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_15),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_207),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_212),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_203),
.B(n_0),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_245),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_249),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_272),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_216),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_194),
.B(n_2),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_258),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_213),
.B(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_249),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_277),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_249),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_325),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_343),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_213),
.B(n_7),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_249),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_249),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_249),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_249),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_249),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_365),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_217),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_259),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_210),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_220),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_360),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_211),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_214),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_226),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_218),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_269),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_219),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_259),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_269),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_227),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_215),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_230),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_239),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_242),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_243),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_254),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_259),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_259),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_222),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_223),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_261),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_283),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_267),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_259),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_208),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_275),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_197),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_231),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_224),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_279),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_294),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_233),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_298),
.Y(n_429)
);

BUFx2_ASAP7_75t_SL g430 ( 
.A(n_283),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_238),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_197),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_260),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_228),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_271),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_308),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_360),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_276),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_237),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_289),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_311),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_319),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_248),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_320),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_253),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_300),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_255),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_306),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_323),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_310),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_316),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_354),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_328),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_329),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_336),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_338),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_354),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_188),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_196),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_199),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_204),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_395),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_423),
.B(n_274),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_370),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_378),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_398),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_399),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_418),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_376),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_388),
.A2(n_252),
.B(n_250),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_401),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_265),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_403),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_397),
.B(n_265),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_421),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_415),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_R g491 ( 
.A(n_416),
.B(n_425),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_434),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_432),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_459),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_460),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_431),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_433),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_439),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_457),
.B(n_302),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_371),
.A2(n_317),
.B1(n_313),
.B2(n_358),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_402),
.B(n_194),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_446),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_405),
.B(n_302),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_377),
.B(n_185),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_379),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_448),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_443),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_445),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_452),
.B(n_192),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_447),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_367),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_390),
.B(n_290),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_393),
.B(n_430),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_454),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_384),
.B(n_341),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_367),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_368),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_375),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_382),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_368),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_374),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_373),
.B(n_290),
.Y(n_531)
);

AND2x4_ASAP7_75t_SL g532 ( 
.A(n_383),
.B(n_221),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_374),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_392),
.B(n_256),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_391),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_392),
.B(n_185),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_396),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_396),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_400),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_400),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_494),
.B(n_407),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_509),
.B(n_406),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_491),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_465),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_481),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_523),
.B(n_423),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_510),
.B(n_221),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_534),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_523),
.A2(n_426),
.B1(n_449),
.B2(n_444),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_530),
.B(n_192),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_517),
.B(n_437),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_509),
.B(n_406),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_487),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_530),
.B(n_232),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_481),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_465),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_469),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_530),
.B(n_232),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_468),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_462),
.B(n_408),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_472),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_474),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_470),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_475),
.B(n_206),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_536),
.B(n_408),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_488),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_494),
.Y(n_577)
);

INVxp33_ASAP7_75t_L g578 ( 
.A(n_527),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_509),
.B(n_409),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_530),
.B(n_234),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_477),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_470),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_511),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_470),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_530),
.B(n_234),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_486),
.A2(n_453),
.B1(n_449),
.B2(n_444),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_509),
.B(n_409),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_521),
.B(n_410),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_529),
.B(n_184),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_482),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_481),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_530),
.B(n_235),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_SL g597 ( 
.A(n_510),
.B(n_201),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_479),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_528),
.B(n_410),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_504),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_535),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_411),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_475),
.B(n_411),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_412),
.Y(n_607)
);

INVx4_ASAP7_75t_SL g608 ( 
.A(n_478),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_492),
.B(n_412),
.Y(n_610)
);

BUFx6f_ASAP7_75t_SL g611 ( 
.A(n_492),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_478),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_517),
.B(n_235),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_531),
.B(n_201),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_478),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_526),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_481),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_508),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_519),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_532),
.B(n_246),
.Y(n_622)
);

BUFx4f_ASAP7_75t_L g623 ( 
.A(n_479),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_467),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_515),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_532),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_479),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_467),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_515),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_503),
.A2(n_312),
.B1(n_266),
.B2(n_369),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_478),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_479),
.A2(n_252),
.B1(n_305),
.B2(n_250),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_471),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_476),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_517),
.B(n_417),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_533),
.B(n_240),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_473),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_532),
.Y(n_639)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_501),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_476),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_501),
.B(n_225),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_480),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_531),
.B(n_417),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_478),
.B(n_501),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_520),
.B(n_419),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_537),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_538),
.B(n_419),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_524),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_480),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

INVx4_ASAP7_75t_SL g653 ( 
.A(n_496),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_520),
.B(n_422),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_540),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_497),
.B(n_229),
.Y(n_657)
);

BUFx4f_ASAP7_75t_L g658 ( 
.A(n_496),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_496),
.B(n_426),
.Y(n_660)
);

AND2x6_ASAP7_75t_L g661 ( 
.A(n_502),
.B(n_251),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_502),
.B(n_251),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_539),
.B(n_427),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_498),
.Y(n_664)
);

BUFx4f_ASAP7_75t_L g665 ( 
.A(n_496),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_498),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_502),
.B(n_280),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_507),
.B(n_429),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_498),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_507),
.B(n_429),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_507),
.B(n_436),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_503),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_498),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_490),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_484),
.B(n_381),
.C(n_436),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_498),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_490),
.B(n_441),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_495),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_495),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_622),
.B(n_221),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_622),
.B(n_221),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_595),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_557),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_595),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_553),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_671),
.B(n_442),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_546),
.B(n_603),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_670),
.B(n_442),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_640),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_670),
.B(n_453),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_598),
.B(n_221),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_578),
.B(n_244),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_575),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_598),
.B(n_236),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_612),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_598),
.B(n_236),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_677),
.B(n_495),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_543),
.B(n_483),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_660),
.B(n_484),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_627),
.A2(n_305),
.B1(n_318),
.B2(n_364),
.Y(n_701)
);

INVx8_ASAP7_75t_L g702 ( 
.A(n_640),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_612),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_606),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_562),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_564),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_576),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_627),
.B(n_209),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_672),
.A2(n_466),
.B1(n_353),
.B2(n_361),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_564),
.Y(n_710)
);

NOR2x1p5_ASAP7_75t_L g711 ( 
.A(n_543),
.B(n_485),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_565),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_583),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_565),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_569),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_623),
.A2(n_499),
.B(n_497),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_623),
.B(n_236),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_601),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_605),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_620),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_619),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_569),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_578),
.B(n_186),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_625),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_645),
.B(n_241),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_630),
.B(n_262),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_648),
.B(n_489),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_619),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_649),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_650),
.B(n_263),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_600),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_570),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_668),
.B(n_542),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_SL g735 ( 
.A1(n_633),
.A2(n_281),
.B(n_355),
.C(n_350),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_556),
.A2(n_513),
.B(n_512),
.C(n_506),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_614),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_570),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_672),
.A2(n_268),
.B(n_321),
.C(n_327),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_579),
.B(n_278),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_573),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_591),
.B(n_186),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_636),
.B(n_187),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_640),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_541),
.B(n_617),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_644),
.B(n_493),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_590),
.B(n_285),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_628),
.A2(n_304),
.B1(n_236),
.B2(n_247),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_646),
.B(n_500),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_550),
.B(n_187),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_654),
.B(n_189),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_551),
.B(n_296),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_592),
.B(n_514),
.Y(n_753)
);

NOR3xp33_ASAP7_75t_L g754 ( 
.A(n_631),
.B(n_516),
.C(n_518),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_604),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_639),
.B(n_497),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_574),
.A2(n_301),
.B1(n_264),
.B2(n_270),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_658),
.A2(n_522),
.B(n_513),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_604),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_593),
.B(n_247),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_552),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_614),
.B(n_282),
.Y(n_762)
);

AND2x2_ASAP7_75t_SL g763 ( 
.A(n_548),
.B(n_466),
.Y(n_763)
);

O2A1O1Ixp5_ASAP7_75t_L g764 ( 
.A1(n_559),
.A2(n_346),
.B(n_513),
.C(n_512),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_597),
.A2(n_303),
.B1(n_292),
.B2(n_287),
.Y(n_765)
);

AND2x4_ASAP7_75t_SL g766 ( 
.A(n_656),
.B(n_247),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_640),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_609),
.Y(n_768)
);

BUFx6f_ASAP7_75t_SL g769 ( 
.A(n_656),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_609),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_573),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_597),
.A2(n_307),
.B1(n_295),
.B2(n_288),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_618),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_637),
.A2(n_314),
.B1(n_299),
.B2(n_291),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_639),
.B(n_247),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_559),
.B(n_499),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_607),
.B(n_190),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_610),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_589),
.B(n_190),
.Y(n_779)
);

NOR2x1p5_ASAP7_75t_L g780 ( 
.A(n_554),
.B(n_353),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_618),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_563),
.B(n_499),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_554),
.B(n_257),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_614),
.A2(n_324),
.B1(n_315),
.B2(n_293),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_563),
.B(n_506),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_624),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_547),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_545),
.B(n_257),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_549),
.B(n_191),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_580),
.B(n_257),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_547),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_585),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_652),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_577),
.B(n_506),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_585),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_580),
.B(n_588),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_634),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_588),
.B(n_257),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_663),
.B(n_337),
.C(n_339),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_629),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_596),
.B(n_512),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_596),
.B(n_522),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_577),
.B(n_191),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_635),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_626),
.B(n_522),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_652),
.B(n_257),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_545),
.B(n_273),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_664),
.B(n_297),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_584),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_642),
.B(n_309),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_584),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_642),
.B(n_326),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_647),
.B(n_330),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_635),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_615),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_560),
.B(n_273),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_614),
.B(n_332),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_615),
.A2(n_642),
.B(n_548),
.C(n_675),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_560),
.B(n_340),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_641),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_641),
.B(n_342),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_572),
.B(n_611),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_674),
.B(n_273),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_586),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_643),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_658),
.A2(n_344),
.B(n_349),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_651),
.B(n_351),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_651),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_586),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_594),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_547),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_674),
.B(n_273),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_614),
.A2(n_284),
.B1(n_198),
.B2(n_195),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_678),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_572),
.B(n_366),
.C(n_331),
.Y(n_835)
);

NAND2x1_ASAP7_75t_L g836 ( 
.A(n_614),
.B(n_273),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_737),
.A2(n_658),
.B(n_665),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_687),
.B(n_567),
.C(n_581),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_800),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_687),
.B(n_656),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_737),
.A2(n_665),
.B(n_561),
.Y(n_841)
);

AOI22x1_ASAP7_75t_L g842 ( 
.A1(n_716),
.A2(n_691),
.B1(n_694),
.B2(n_685),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_737),
.A2(n_544),
.B(n_566),
.Y(n_843)
);

BUFx12f_ASAP7_75t_L g844 ( 
.A(n_797),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_682),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_800),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_700),
.B(n_679),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_734),
.B(n_594),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_731),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_761),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_794),
.B(n_621),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_698),
.B(n_657),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_748),
.A2(n_362),
.B1(n_363),
.B2(n_657),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_745),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_793),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_748),
.B(n_743),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_779),
.B(n_634),
.C(n_638),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_743),
.B(n_555),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_693),
.B(n_621),
.Y(n_859)
);

INVx11_ASAP7_75t_L g860 ( 
.A(n_769),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_732),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_686),
.B(n_555),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_793),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_803),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_688),
.B(n_638),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_742),
.B(n_571),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_693),
.B(n_599),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_779),
.B(n_335),
.C(n_333),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_697),
.A2(n_582),
.B(n_571),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_717),
.A2(n_676),
.B(n_669),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_750),
.A2(n_667),
.B1(n_662),
.B2(n_661),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_796),
.A2(n_782),
.B(n_776),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_742),
.B(n_571),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_701),
.B(n_582),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_739),
.A2(n_681),
.B(n_680),
.C(n_818),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_582),
.Y(n_876)
);

AND2x2_ASAP7_75t_SL g877 ( 
.A(n_763),
.B(n_621),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_750),
.A2(n_613),
.B(n_659),
.C(n_666),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_R g879 ( 
.A(n_769),
.B(n_602),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_805),
.B(n_655),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_690),
.A2(n_611),
.B1(n_667),
.B2(n_662),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_815),
.B(n_602),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_682),
.Y(n_883)
);

INVx11_ASAP7_75t_L g884 ( 
.A(n_809),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_684),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_818),
.A2(n_666),
.B(n_357),
.C(n_356),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_778),
.B(n_568),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_680),
.A2(n_611),
.B1(n_667),
.B2(n_662),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_740),
.B(n_547),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_684),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_747),
.B(n_707),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_SL g892 ( 
.A(n_799),
.B(n_352),
.C(n_334),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_763),
.A2(n_661),
.B1(n_667),
.B2(n_662),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_811),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_739),
.A2(n_667),
.B(n_662),
.C(n_661),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_751),
.B(n_655),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_713),
.B(n_587),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_708),
.A2(n_566),
.B(n_632),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_755),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_718),
.B(n_587),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_719),
.B(n_587),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_789),
.B(n_193),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_704),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_681),
.A2(n_667),
.B(n_662),
.C(n_661),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_703),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_720),
.A2(n_347),
.B1(n_348),
.B2(n_193),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_728),
.A2(n_673),
.B(n_587),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_789),
.B(n_655),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_780),
.Y(n_909)
);

BUFx8_ASAP7_75t_L g910 ( 
.A(n_749),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_683),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_724),
.A2(n_200),
.B1(n_202),
.B2(n_205),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_783),
.A2(n_616),
.B1(n_357),
.B2(n_356),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_728),
.A2(n_616),
.B(n_608),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_L g915 ( 
.A(n_723),
.B(n_803),
.C(n_777),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_783),
.A2(n_616),
.B1(n_359),
.B2(n_202),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_796),
.A2(n_359),
.B(n_205),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_729),
.A2(n_364),
.B1(n_304),
.B2(n_286),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_760),
.A2(n_608),
.B(n_10),
.C(n_11),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_759),
.B(n_768),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_753),
.B(n_8),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_822),
.A2(n_608),
.B1(n_364),
.B2(n_304),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_703),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_770),
.B(n_653),
.Y(n_924)
);

OA22x2_ASAP7_75t_L g925 ( 
.A1(n_746),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_736),
.A2(n_286),
.B(n_304),
.C(n_364),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_696),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_813),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_835),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_767),
.B(n_727),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_773),
.B(n_364),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_709),
.B(n_17),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_822),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_781),
.B(n_304),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_744),
.B(n_286),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_767),
.B(n_286),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_786),
.B(n_286),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_787),
.A2(n_181),
.B(n_177),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_764),
.A2(n_172),
.B(n_163),
.Y(n_939)
);

INVx3_ASAP7_75t_SL g940 ( 
.A(n_766),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_699),
.B(n_149),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_696),
.Y(n_942)
);

AO22x1_ASAP7_75t_L g943 ( 
.A1(n_754),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_775),
.A2(n_730),
.B(n_726),
.C(n_752),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_709),
.B(n_21),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_810),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_757),
.B(n_24),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_774),
.B(n_25),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_787),
.A2(n_142),
.B(n_138),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_785),
.A2(n_801),
.B(n_802),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_711),
.B(n_132),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_756),
.A2(n_820),
.B1(n_825),
.B2(n_804),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_831),
.A2(n_128),
.B(n_121),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_766),
.B(n_25),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_831),
.A2(n_115),
.B(n_112),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_812),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_765),
.B(n_26),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_814),
.B(n_27),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_828),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_834),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_772),
.B(n_31),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_696),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_808),
.B(n_94),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_791),
.A2(n_87),
.B(n_85),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_821),
.A2(n_83),
.B1(n_74),
.B2(n_69),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_833),
.A2(n_32),
.B(n_34),
.C(n_37),
.Y(n_966)
);

AO21x2_ASAP7_75t_L g967 ( 
.A1(n_775),
.A2(n_65),
.B(n_38),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_725),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_762),
.A2(n_34),
.B(n_40),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_784),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_817),
.A2(n_46),
.B(n_48),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_696),
.Y(n_972)
);

OA22x2_ASAP7_75t_L g973 ( 
.A1(n_790),
.A2(n_798),
.B1(n_826),
.B2(n_827),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_721),
.B(n_49),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_819),
.A2(n_52),
.B(n_54),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_689),
.A2(n_702),
.B(n_721),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_689),
.A2(n_702),
.B(n_721),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_705),
.A2(n_722),
.B(n_830),
.C(n_706),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_710),
.A2(n_771),
.B1(n_829),
.B2(n_712),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_714),
.A2(n_738),
.B(n_795),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_689),
.A2(n_702),
.B(n_721),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_836),
.A2(n_758),
.B(n_733),
.C(n_824),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_715),
.A2(n_741),
.B(n_792),
.C(n_735),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_806),
.A2(n_823),
.B(n_832),
.C(n_816),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_832),
.A2(n_823),
.B(n_807),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_816),
.A2(n_687),
.B(n_546),
.C(n_779),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_788),
.A2(n_623),
.B(n_598),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_788),
.B(n_807),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_793),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_687),
.B(n_700),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_687),
.B(n_700),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_737),
.A2(n_623),
.B(n_598),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_687),
.B(n_700),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_687),
.B(n_546),
.C(n_779),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_737),
.A2(n_623),
.B(n_598),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_737),
.A2(n_623),
.B(n_598),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_L g997 ( 
.A1(n_687),
.A2(n_546),
.B(n_750),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_850),
.Y(n_998)
);

OAI21x1_ASAP7_75t_SL g999 ( 
.A1(n_875),
.A2(n_971),
.B(n_969),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_997),
.A2(n_994),
.B1(n_915),
.B2(n_947),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_888),
.B(n_881),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_990),
.A2(n_991),
.B1(n_993),
.B2(n_856),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_R g1003 ( 
.A(n_894),
.B(n_892),
.Y(n_1003)
);

NOR2x1_ASAP7_75t_L g1004 ( 
.A(n_880),
.B(n_857),
.Y(n_1004)
);

OAI22x1_ASAP7_75t_L g1005 ( 
.A1(n_945),
.A2(n_908),
.B1(n_921),
.B2(n_932),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_927),
.B(n_972),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_854),
.B(n_990),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_991),
.B(n_968),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_968),
.B(n_864),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_986),
.A2(n_877),
.B1(n_848),
.B2(n_957),
.Y(n_1010)
);

NAND2xp33_ASAP7_75t_L g1011 ( 
.A(n_896),
.B(n_946),
.Y(n_1011)
);

AO31x2_ASAP7_75t_L g1012 ( 
.A1(n_878),
.A2(n_886),
.A3(n_926),
.B(n_983),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_948),
.A2(n_917),
.B(n_956),
.C(n_868),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_917),
.A2(n_865),
.B(n_944),
.C(n_929),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_848),
.A2(n_893),
.B1(n_847),
.B2(n_871),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_891),
.B(n_852),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_987),
.A2(n_995),
.B(n_992),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_982),
.A2(n_872),
.B(n_870),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_SL g1019 ( 
.A1(n_904),
.A2(n_895),
.B(n_976),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_851),
.B(n_859),
.Y(n_1020)
);

OA22x2_ASAP7_75t_L g1021 ( 
.A1(n_928),
.A2(n_961),
.B1(n_970),
.B2(n_909),
.Y(n_1021)
);

NAND2x1_ASAP7_75t_L g1022 ( 
.A(n_927),
.B(n_972),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_902),
.B(n_890),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_996),
.A2(n_837),
.B(n_898),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_890),
.B(n_849),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_950),
.A2(n_973),
.B(n_876),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_861),
.B(n_899),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_903),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_874),
.A2(n_925),
.B1(n_853),
.B2(n_973),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_959),
.B(n_862),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_866),
.A2(n_873),
.B(n_858),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_840),
.B(n_845),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_910),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_984),
.A2(n_966),
.A3(n_918),
.B(n_934),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_863),
.B(n_989),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_907),
.A2(n_842),
.B(n_841),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_SL g1037 ( 
.A(n_927),
.B(n_972),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_869),
.A2(n_975),
.B(n_919),
.C(n_867),
.Y(n_1038)
);

AOI211x1_ASAP7_75t_L g1039 ( 
.A1(n_943),
.A2(n_970),
.B(n_853),
.C(n_912),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_843),
.A2(n_980),
.B(n_914),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_942),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_980),
.A2(n_950),
.B(n_977),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_978),
.A2(n_939),
.B(n_985),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_918),
.A2(n_931),
.A3(n_937),
.B(n_960),
.Y(n_1044)
);

BUFx5_ASAP7_75t_L g1045 ( 
.A(n_839),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_889),
.B(n_911),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_981),
.A2(n_979),
.B(n_924),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_939),
.A2(n_952),
.B(n_838),
.C(n_974),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_845),
.B(n_923),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_884),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_979),
.A2(n_963),
.B(n_922),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_844),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_935),
.A2(n_897),
.B(n_900),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_901),
.A2(n_942),
.B(n_962),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_846),
.A2(n_949),
.B(n_955),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_910),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_882),
.B(n_933),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_941),
.A2(n_958),
.B(n_965),
.C(n_916),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_936),
.A2(n_913),
.B(n_964),
.Y(n_1059)
);

OA22x2_ASAP7_75t_L g1060 ( 
.A1(n_887),
.A2(n_954),
.B1(n_925),
.B2(n_940),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_845),
.B(n_923),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_938),
.A2(n_953),
.B(n_930),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_883),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_883),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_935),
.A2(n_988),
.B(n_905),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_883),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_885),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_879),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_951),
.A2(n_912),
.B(n_906),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_885),
.B(n_905),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_885),
.A2(n_905),
.B(n_923),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_906),
.A2(n_878),
.A3(n_886),
.B(n_926),
.Y(n_1072)
);

O2A1O1Ixp5_ASAP7_75t_L g1073 ( 
.A1(n_967),
.A2(n_856),
.B(n_986),
.C(n_915),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_967),
.A2(n_860),
.B(n_997),
.C(n_994),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_850),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_920),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_878),
.A2(n_886),
.A3(n_926),
.B(n_983),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_870),
.A2(n_695),
.B(n_692),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_845),
.B(n_883),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_990),
.A2(n_748),
.B1(n_991),
.B2(n_993),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_844),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_856),
.A2(n_875),
.B(n_994),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_850),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_880),
.B(n_687),
.Y(n_1087)
);

OA22x2_ASAP7_75t_L g1088 ( 
.A1(n_997),
.A2(n_503),
.B1(n_550),
.B2(n_815),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_SL g1089 ( 
.A1(n_875),
.A2(n_971),
.B(n_969),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_870),
.A2(n_695),
.B(n_692),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_994),
.B(n_745),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_997),
.B(n_994),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_856),
.A2(n_875),
.B(n_994),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_993),
.B(n_990),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_993),
.B(n_990),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_856),
.A2(n_875),
.B(n_994),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_993),
.B(n_990),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_993),
.B(n_990),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_L g1101 ( 
.A(n_844),
.B(n_797),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_994),
.B(n_997),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_870),
.A2(n_695),
.B(n_692),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_994),
.B(n_745),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_990),
.A2(n_748),
.B1(n_991),
.B2(n_993),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_SL g1108 ( 
.A1(n_875),
.A2(n_971),
.B(n_969),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_855),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_993),
.B(n_990),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_845),
.B(n_883),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_878),
.A2(n_886),
.A3(n_926),
.B(n_983),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_920),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_880),
.B(n_687),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_855),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_920),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_870),
.A2(n_695),
.B(n_692),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_993),
.B(n_990),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_997),
.B(n_994),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_856),
.A2(n_875),
.B(n_994),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_880),
.B(n_687),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_855),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_993),
.B(n_990),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_994),
.B(n_997),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_850),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_982),
.A2(n_872),
.B(n_987),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_994),
.B(n_997),
.C(n_750),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_997),
.A2(n_994),
.B(n_915),
.C(n_856),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_927),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_870),
.A2(n_695),
.B(n_692),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1127),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1027),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1075),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_998),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1063),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1043),
.A2(n_1016),
.B(n_1019),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1008),
.B(n_1101),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1129),
.A2(n_1121),
.B(n_1092),
.C(n_1013),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1061),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1075),
.Y(n_1143)
);

AOI211xp5_ASAP7_75t_L g1144 ( 
.A1(n_1010),
.A2(n_1126),
.B(n_1102),
.C(n_1014),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1073),
.A2(n_1094),
.B(n_1084),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_R g1147 ( 
.A(n_1068),
.B(n_1052),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1005),
.A2(n_1088),
.B1(n_1000),
.B2(n_1010),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1070),
.B(n_1080),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1086),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_1028),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1061),
.B(n_1071),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1061),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1067),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1111),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1123),
.B(n_1020),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1009),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1098),
.B(n_1100),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1111),
.B(n_1064),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1098),
.B(n_1100),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1043),
.A2(n_1026),
.B(n_1018),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_SL g1163 ( 
.A(n_1050),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1007),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1165)
);

OR2x6_ASAP7_75t_SL g1166 ( 
.A(n_1083),
.B(n_1105),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1066),
.B(n_1004),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1120),
.B(n_1125),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1022),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1049),
.Y(n_1170)
);

OR2x6_ASAP7_75t_L g1171 ( 
.A(n_1033),
.B(n_1056),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1006),
.Y(n_1172)
);

BUFx8_ASAP7_75t_SL g1173 ( 
.A(n_1131),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1110),
.B(n_1120),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1109),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1125),
.A2(n_1106),
.B1(n_1081),
.B2(n_1002),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1002),
.B(n_1081),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1106),
.B(n_1076),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1041),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1011),
.Y(n_1180)
);

OAI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_1088),
.A2(n_1130),
.B(n_1084),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1115),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1006),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1032),
.B(n_1037),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1003),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1058),
.A2(n_1122),
.B(n_1094),
.C(n_1097),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1041),
.Y(n_1188)
);

CKINVDCx6p67_ASAP7_75t_R g1189 ( 
.A(n_1023),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1021),
.B(n_1060),
.Y(n_1190)
);

NAND2x1_ASAP7_75t_L g1191 ( 
.A(n_1124),
.B(n_999),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1021),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1035),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1025),
.B(n_1065),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1060),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1045),
.Y(n_1196)
);

BUFx4f_ASAP7_75t_SL g1197 ( 
.A(n_1045),
.Y(n_1197)
);

BUFx12f_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1097),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1036),
.A2(n_1024),
.B(n_1128),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_1001),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1074),
.B(n_1069),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1122),
.B(n_1048),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1030),
.B(n_1046),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1046),
.B(n_1015),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1045),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1038),
.B(n_1026),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1015),
.B(n_1039),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1029),
.A2(n_1051),
.B1(n_1059),
.B2(n_1053),
.Y(n_1209)
);

INVx3_ASAP7_75t_SL g1210 ( 
.A(n_1045),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1045),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1047),
.B(n_1054),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_1029),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1042),
.Y(n_1214)
);

AO21x2_ASAP7_75t_L g1215 ( 
.A1(n_1089),
.A2(n_1108),
.B(n_1031),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1062),
.B(n_1055),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1072),
.B(n_1001),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1040),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1001),
.A2(n_1034),
.B1(n_1044),
.B2(n_1012),
.C(n_1112),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_SL g1220 ( 
.A(n_1034),
.B(n_1132),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1078),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1078),
.B(n_1112),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1077),
.A2(n_1099),
.B(n_1118),
.C(n_1117),
.Y(n_1223)
);

AO21x1_ASAP7_75t_L g1224 ( 
.A1(n_1079),
.A2(n_1119),
.B(n_1104),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1112),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1090),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1082),
.B(n_1107),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1085),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1093),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1044),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1103),
.B(n_993),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1052),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1068),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1020),
.B(n_951),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1087),
.B(n_997),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1129),
.A2(n_997),
.B1(n_994),
.B2(n_687),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1127),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1061),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1068),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1027),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1095),
.B(n_993),
.Y(n_1243)
);

INVx8_ASAP7_75t_L g1244 ( 
.A(n_1063),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1095),
.B(n_993),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1013),
.A2(n_997),
.B(n_994),
.C(n_986),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1110),
.B(n_993),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_998),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1033),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1095),
.B(n_993),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1061),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1052),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1027),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1087),
.B(n_880),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1258)
);

OR2x2_ASAP7_75t_SL g1259 ( 
.A(n_1129),
.B(n_994),
.Y(n_1259)
);

INVxp67_ASAP7_75t_SL g1260 ( 
.A(n_998),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1095),
.B(n_993),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1027),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1027),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_998),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1063),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1075),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1127),
.Y(n_1271)
);

BUFx2_ASAP7_75t_R g1272 ( 
.A(n_1166),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1199),
.B(n_1174),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1184),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1148),
.A2(n_1181),
.B1(n_1203),
.B2(n_1213),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1239),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1136),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1195),
.A2(n_1198),
.B1(n_1201),
.B2(n_1180),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1236),
.A2(n_1247),
.B1(n_1180),
.B2(n_1245),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1197),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1181),
.A2(n_1236),
.B1(n_1235),
.B2(n_1145),
.Y(n_1281)
);

BUFx2_ASAP7_75t_R g1282 ( 
.A(n_1173),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1239),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1145),
.A2(n_1192),
.B1(n_1165),
.B2(n_1209),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1239),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1149),
.B(n_1167),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1233),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1175),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1151),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1252),
.B(n_1201),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1135),
.B(n_1237),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1252),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1182),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1190),
.B(n_1146),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1209),
.A2(n_1177),
.B1(n_1207),
.B2(n_1176),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1255),
.B(n_1258),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1243),
.A2(n_1245),
.B1(n_1251),
.B2(n_1261),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1146),
.B(n_1154),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1252),
.Y(n_1300)
);

AO21x1_ASAP7_75t_L g1301 ( 
.A1(n_1144),
.A2(n_1246),
.B(n_1176),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1243),
.A2(n_1251),
.B1(n_1261),
.B2(n_1159),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1269),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1151),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1227),
.A2(n_1216),
.B(n_1229),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1172),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1232),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1141),
.B(n_1144),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1134),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1242),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1227),
.A2(n_1216),
.B(n_1229),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1256),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1262),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1264),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1238),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1158),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1271),
.Y(n_1317)
);

BUFx2_ASAP7_75t_R g1318 ( 
.A(n_1186),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1164),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1254),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1263),
.B(n_1265),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1164),
.Y(n_1322)
);

INVx8_ASAP7_75t_L g1323 ( 
.A(n_1244),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1250),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1154),
.B(n_1161),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1241),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1249),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1253),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1177),
.A2(n_1157),
.B1(n_1168),
.B2(n_1139),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1149),
.B(n_1167),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1257),
.A2(n_1234),
.B1(n_1208),
.B2(n_1178),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1133),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1137),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1259),
.B(n_1268),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1225),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1234),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1172),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1260),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1270),
.Y(n_1339)
);

BUFx12f_ASAP7_75t_L g1340 ( 
.A(n_1267),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1234),
.A2(n_1202),
.B1(n_1208),
.B2(n_1244),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1162),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1156),
.B(n_1160),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1187),
.B(n_1204),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1172),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1140),
.B(n_1178),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_1150),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1183),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1170),
.Y(n_1349)
);

BUFx2_ASAP7_75t_R g1350 ( 
.A(n_1240),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1214),
.A2(n_1191),
.B(n_1231),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1221),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_SL g1353 ( 
.A(n_1138),
.Y(n_1353)
);

INVx6_ASAP7_75t_SL g1354 ( 
.A(n_1171),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1147),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1179),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1155),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1214),
.A2(n_1224),
.B(n_1217),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1234),
.A2(n_1205),
.B1(n_1202),
.B2(n_1219),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1188),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1248),
.B(n_1266),
.Y(n_1361)
);

AO21x2_ASAP7_75t_L g1362 ( 
.A1(n_1223),
.A2(n_1215),
.B(n_1205),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1162),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1215),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1222),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1206),
.A2(n_1211),
.B(n_1152),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1230),
.A2(n_1222),
.B(n_1212),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1189),
.A2(n_1226),
.B1(n_1142),
.B2(n_1153),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1196),
.A2(n_1220),
.B(n_1228),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1185),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1194),
.A2(n_1171),
.B1(n_1185),
.B2(n_1142),
.Y(n_1371)
);

BUFx2_ASAP7_75t_R g1372 ( 
.A(n_1210),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1152),
.B(n_1220),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1244),
.A2(n_1267),
.B1(n_1171),
.B2(n_1163),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1152),
.A2(n_1163),
.B1(n_1183),
.B2(n_1169),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1267),
.B(n_1169),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1218),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1184),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1239),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1174),
.B(n_993),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1149),
.B(n_1167),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1184),
.Y(n_1382)
);

BUFx8_ASAP7_75t_SL g1383 ( 
.A(n_1232),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1199),
.A2(n_994),
.B1(n_997),
.B2(n_993),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1184),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1238),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1135),
.B(n_1237),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1239),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1173),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1190),
.B(n_1148),
.Y(n_1390)
);

BUFx2_ASAP7_75t_SL g1391 ( 
.A(n_1163),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1173),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1184),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1200),
.A2(n_1036),
.B(n_1017),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1193),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1250),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1184),
.Y(n_1397)
);

CKINVDCx6p67_ASAP7_75t_R g1398 ( 
.A(n_1287),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1308),
.A2(n_1301),
.B1(n_1275),
.B2(n_1384),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1319),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1364),
.A2(n_1363),
.A3(n_1342),
.B(n_1335),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1367),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1336),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1322),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1367),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1344),
.B(n_1294),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1367),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1299),
.B(n_1325),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1366),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1299),
.B(n_1325),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1377),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1308),
.A2(n_1290),
.B(n_1302),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1352),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1273),
.B(n_1380),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1287),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1369),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1273),
.A2(n_1275),
.B1(n_1278),
.B2(n_1281),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1390),
.B(n_1296),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1390),
.B(n_1296),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1394),
.A2(n_1311),
.B(n_1305),
.Y(n_1421)
);

INVx11_ASAP7_75t_L g1422 ( 
.A(n_1340),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1323),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1365),
.B(n_1373),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1338),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1277),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1291),
.B(n_1297),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1304),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1284),
.B(n_1281),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1284),
.B(n_1359),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1351),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1346),
.B(n_1329),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1329),
.B(n_1359),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1377),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1358),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1362),
.A2(n_1351),
.B(n_1358),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1362),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1331),
.A2(n_1371),
.B(n_1314),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1334),
.B(n_1395),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1309),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1310),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1312),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1326),
.B(n_1327),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1313),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1334),
.B(n_1331),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1336),
.B(n_1370),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1336),
.B(n_1286),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1321),
.B(n_1387),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1288),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1328),
.B(n_1339),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1290),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1298),
.A2(n_1279),
.B(n_1356),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1293),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1316),
.B(n_1274),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1292),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1378),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1303),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1382),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1385),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1393),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1397),
.B(n_1286),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1333),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1303),
.B(n_1289),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1354),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1292),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1354),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1292),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1315),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1341),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1285),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1295),
.B(n_1317),
.Y(n_1471)
);

INVx8_ASAP7_75t_L g1472 ( 
.A(n_1323),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1276),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1357),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1386),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1286),
.B(n_1330),
.Y(n_1476)
);

OR2x6_ASAP7_75t_L g1477 ( 
.A(n_1323),
.B(n_1368),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1330),
.B(n_1381),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1276),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1283),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1355),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1283),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1349),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1361),
.B(n_1381),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1417),
.A2(n_1381),
.B1(n_1330),
.B2(n_1343),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1406),
.B(n_1360),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1406),
.B(n_1360),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1402),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1402),
.B(n_1332),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1432),
.B(n_1375),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1432),
.B(n_1300),
.Y(n_1491)
);

AOI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1437),
.A2(n_1376),
.B(n_1348),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1405),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1401),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1403),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1410),
.B(n_1408),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1410),
.B(n_1388),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1457),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1416),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1407),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1440),
.B(n_1388),
.Y(n_1501)
);

NAND2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1403),
.B(n_1379),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1446),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1399),
.A2(n_1354),
.B1(n_1396),
.B2(n_1324),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1407),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1398),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1425),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1413),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1437),
.A2(n_1345),
.B(n_1348),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1434),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1424),
.B(n_1337),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1414),
.B(n_1318),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1439),
.B(n_1337),
.Y(n_1513)
);

BUFx2_ASAP7_75t_SL g1514 ( 
.A(n_1411),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1439),
.B(n_1337),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1445),
.B(n_1337),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1445),
.B(n_1306),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1409),
.B(n_1391),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1440),
.B(n_1306),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1463),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1434),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1442),
.B(n_1306),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1442),
.B(n_1300),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1400),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1444),
.B(n_1306),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1444),
.B(n_1345),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1520),
.B(n_1404),
.Y(n_1527)
);

NOR3xp33_ASAP7_75t_L g1528 ( 
.A(n_1490),
.B(n_1469),
.C(n_1374),
.Y(n_1528)
);

OAI21xp33_ASAP7_75t_L g1529 ( 
.A1(n_1490),
.A2(n_1412),
.B(n_1430),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1504),
.A2(n_1429),
.B1(n_1430),
.B2(n_1469),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1520),
.B(n_1426),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1504),
.A2(n_1433),
.B1(n_1462),
.B2(n_1412),
.C(n_1466),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1485),
.A2(n_1272),
.B1(n_1433),
.B2(n_1429),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1516),
.B(n_1409),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1516),
.B(n_1435),
.Y(n_1536)
);

OAI21xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1485),
.A2(n_1420),
.B(n_1419),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1494),
.A2(n_1421),
.B(n_1431),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1524),
.B(n_1468),
.Y(n_1539)
);

NAND2xp33_ASAP7_75t_L g1540 ( 
.A(n_1518),
.B(n_1285),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1518),
.B(n_1467),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1496),
.B(n_1458),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1496),
.B(n_1458),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1514),
.A2(n_1420),
.B1(n_1419),
.B2(n_1438),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1459),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1507),
.B(n_1459),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1498),
.B(n_1460),
.Y(n_1547)
);

NAND4xp25_ASAP7_75t_L g1548 ( 
.A(n_1491),
.B(n_1463),
.C(n_1483),
.D(n_1471),
.Y(n_1548)
);

NAND4xp25_ASAP7_75t_L g1549 ( 
.A(n_1491),
.B(n_1483),
.C(n_1443),
.D(n_1454),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1512),
.A2(n_1466),
.B(n_1464),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1517),
.B(n_1438),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1513),
.B(n_1438),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1501),
.B(n_1473),
.C(n_1482),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1510),
.A2(n_1477),
.B1(n_1447),
.B2(n_1452),
.Y(n_1554)
);

NAND4xp25_ASAP7_75t_L g1555 ( 
.A(n_1489),
.B(n_1443),
.C(n_1454),
.D(n_1450),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1494),
.A2(n_1421),
.B(n_1431),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1473),
.C(n_1479),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_L g1558 ( 
.A1(n_1498),
.A2(n_1464),
.B1(n_1474),
.B2(n_1484),
.C(n_1411),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1497),
.B(n_1460),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1513),
.B(n_1438),
.Y(n_1560)
);

AND2x2_ASAP7_75t_SL g1561 ( 
.A(n_1509),
.B(n_1447),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1497),
.B(n_1456),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1503),
.B(n_1467),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1515),
.B(n_1418),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1489),
.B(n_1456),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1510),
.A2(n_1477),
.B1(n_1447),
.B2(n_1452),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1495),
.B(n_1470),
.C(n_1455),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1519),
.B(n_1450),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_1418),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1511),
.B(n_1461),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1510),
.A2(n_1477),
.B1(n_1447),
.B2(n_1452),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1486),
.B(n_1461),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1523),
.B(n_1482),
.C(n_1480),
.Y(n_1573)
);

NOR2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1521),
.B(n_1398),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1514),
.A2(n_1477),
.B1(n_1427),
.B2(n_1372),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1486),
.B(n_1431),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1487),
.B(n_1436),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1519),
.B(n_1522),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1522),
.B(n_1475),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1525),
.B(n_1441),
.Y(n_1580)
);

NOR2xp67_ASAP7_75t_L g1581 ( 
.A(n_1499),
.B(n_1479),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1525),
.B(n_1441),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1523),
.A2(n_1484),
.B1(n_1477),
.B2(n_1347),
.C(n_1448),
.Y(n_1583)
);

NAND4xp25_ASAP7_75t_L g1584 ( 
.A(n_1526),
.B(n_1448),
.C(n_1453),
.D(n_1449),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1521),
.A2(n_1478),
.B1(n_1476),
.B2(n_1451),
.Y(n_1585)
);

AOI21xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1506),
.A2(n_1415),
.B(n_1323),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1581),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1581),
.B(n_1499),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1488),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1543),
.B(n_1565),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1561),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1562),
.B(n_1488),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1509),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1561),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1547),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1569),
.B(n_1499),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1538),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1577),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1577),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1560),
.B(n_1509),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1576),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1545),
.B(n_1493),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1546),
.B(n_1493),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1538),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1556),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1527),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1556),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1531),
.B(n_1500),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1555),
.B(n_1500),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1536),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1556),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1564),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1559),
.B(n_1505),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1534),
.B(n_1505),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1558),
.B(n_1521),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1574),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1536),
.B(n_1508),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1553),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1608),
.B(n_1572),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1603),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1591),
.B(n_1570),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1615),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1620),
.A2(n_1529),
.B1(n_1533),
.B2(n_1528),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1623),
.B(n_1612),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1608),
.B(n_1572),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1591),
.B(n_1570),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1549),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1615),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1591),
.B(n_1544),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1621),
.B(n_1574),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1588),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1623),
.B(n_1535),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1595),
.B(n_1619),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1603),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1595),
.B(n_1579),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1590),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1595),
.B(n_1539),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1503),
.Y(n_1644)
);

INVx3_ASAP7_75t_R g1645 ( 
.A(n_1612),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1601),
.B(n_1503),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1601),
.B(n_1503),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1598),
.B(n_1503),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1612),
.B(n_1548),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1598),
.B(n_1503),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1587),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1621),
.B(n_1567),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1620),
.A2(n_1537),
.B1(n_1575),
.B2(n_1550),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1603),
.Y(n_1656)
);

AOI32xp33_ASAP7_75t_L g1657 ( 
.A1(n_1594),
.A2(n_1537),
.A3(n_1540),
.B1(n_1530),
.B2(n_1585),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1622),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1598),
.B(n_1554),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1621),
.A2(n_1571),
.B1(n_1566),
.B2(n_1532),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1619),
.B(n_1557),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1590),
.Y(n_1662)
);

NAND2x1_ASAP7_75t_L g1663 ( 
.A(n_1594),
.B(n_1573),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1587),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1625),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1636),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1629),
.B(n_1617),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1638),
.Y(n_1671)
);

NAND4xp25_ASAP7_75t_L g1672 ( 
.A(n_1628),
.B(n_1583),
.C(n_1586),
.D(n_1611),
.Y(n_1672)
);

BUFx8_ASAP7_75t_SL g1673 ( 
.A(n_1636),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1661),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1627),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1640),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1662),
.B(n_1618),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1640),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1635),
.B(n_1598),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1654),
.A2(n_1621),
.B1(n_1540),
.B2(n_1541),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1656),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1656),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1627),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1639),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1634),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1636),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1626),
.B(n_1593),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1634),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1626),
.B(n_1593),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1645),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1638),
.B(n_1324),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1631),
.B(n_1593),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1655),
.B(n_1618),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1588),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1631),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1659),
.B(n_1599),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1644),
.Y(n_1701)
);

CKINVDCx14_ASAP7_75t_R g1702 ( 
.A(n_1659),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1643),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1655),
.B(n_1605),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1652),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1653),
.B(n_1599),
.Y(n_1706)
);

OAI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1657),
.A2(n_1611),
.B(n_1605),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1705),
.B(n_1650),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1686),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1694),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1705),
.B(n_1650),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1706),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1687),
.B(n_1653),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1670),
.B(n_1689),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1695),
.B(n_1663),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1674),
.B(n_1633),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1665),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1687),
.B(n_1663),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1702),
.B(n_1633),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1706),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1665),
.Y(n_1721)
);

AND3x2_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1664),
.C(n_1651),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1669),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1688),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1707),
.B(n_1660),
.C(n_1641),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1687),
.B(n_1637),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1676),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1688),
.Y(n_1729)
);

AO21x2_ASAP7_75t_L g1730 ( 
.A1(n_1676),
.A2(n_1645),
.B(n_1610),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_SL g1731 ( 
.A1(n_1679),
.A2(n_1651),
.B1(n_1649),
.B2(n_1647),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1673),
.B(n_1396),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1670),
.B(n_1624),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1678),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1680),
.B(n_1586),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1667),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1667),
.A2(n_1630),
.B1(n_1600),
.B2(n_1648),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1679),
.B(n_1637),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1698),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1678),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1672),
.A2(n_1649),
.B1(n_1647),
.B2(n_1644),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1703),
.B(n_1618),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_1622),
.Y(n_1743)
);

AOI21xp33_ASAP7_75t_SL g1744 ( 
.A1(n_1735),
.A2(n_1355),
.B(n_1692),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1721),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1726),
.B(n_1736),
.C(n_1719),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1739),
.Y(n_1747)
);

NAND4xp75_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1666),
.C(n_1700),
.D(n_1697),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1710),
.B(n_1692),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1710),
.B(n_1666),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1739),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1732),
.A2(n_1389),
.B1(n_1392),
.B2(n_1481),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1727),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1741),
.B(n_1701),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1722),
.A2(n_1698),
.B1(n_1701),
.B2(n_1693),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1709),
.B(n_1693),
.Y(n_1756)
);

NOR3x1_ASAP7_75t_L g1757 ( 
.A(n_1708),
.B(n_1704),
.C(n_1677),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1721),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1708),
.B(n_1383),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_SL g1760 ( 
.A(n_1711),
.B(n_1704),
.C(n_1700),
.Y(n_1760)
);

AOI211xp5_ASAP7_75t_L g1761 ( 
.A1(n_1711),
.A2(n_1698),
.B(n_1684),
.C(n_1699),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1731),
.A2(n_1699),
.B1(n_1668),
.B2(n_1600),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_SL g1763 ( 
.A(n_1718),
.B(n_1684),
.C(n_1691),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1717),
.B(n_1681),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1724),
.Y(n_1765)
);

OAI322xp33_ASAP7_75t_L g1766 ( 
.A1(n_1714),
.A2(n_1682),
.A3(n_1681),
.B1(n_1685),
.B2(n_1690),
.C1(n_1683),
.C2(n_1675),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1712),
.A2(n_1646),
.B1(n_1691),
.B2(n_1696),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1724),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1713),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1759),
.B(n_1714),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1747),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1745),
.Y(n_1772)
);

NAND2x1_ASAP7_75t_SL g1773 ( 
.A(n_1755),
.B(n_1718),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1769),
.B(n_1712),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1748),
.A2(n_1720),
.B1(n_1716),
.B2(n_1733),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1751),
.B(n_1720),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1758),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1750),
.B(n_1733),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1749),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1753),
.B(n_1713),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1757),
.B(n_1738),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1752),
.B(n_1389),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1746),
.A2(n_1737),
.B1(n_1743),
.B2(n_1738),
.C(n_1725),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1761),
.B(n_1727),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1760),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1765),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1754),
.B(n_1725),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1744),
.A2(n_1743),
.B1(n_1729),
.B2(n_1742),
.C(n_1734),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1763),
.B(n_1392),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1785),
.A2(n_1762),
.B1(n_1767),
.B2(n_1756),
.C(n_1764),
.Y(n_1790)
);

AOI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1789),
.A2(n_1762),
.B(n_1766),
.C(n_1756),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1783),
.A2(n_1729),
.B1(n_1764),
.B2(n_1727),
.Y(n_1792)
);

NAND4xp25_ASAP7_75t_L g1793 ( 
.A(n_1770),
.B(n_1768),
.C(n_1740),
.D(n_1728),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1781),
.A2(n_1723),
.B1(n_1740),
.B2(n_1728),
.C(n_1730),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1771),
.B(n_1730),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1773),
.A2(n_1730),
.B(n_1614),
.C(n_1682),
.Y(n_1796)
);

OAI321xp33_ASAP7_75t_L g1797 ( 
.A1(n_1775),
.A2(n_1685),
.A3(n_1696),
.B1(n_1690),
.B2(n_1683),
.C(n_1675),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1779),
.A2(n_1614),
.B(n_1606),
.C(n_1646),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1781),
.B(n_1599),
.Y(n_1799)
);

OA22x2_ASAP7_75t_L g1800 ( 
.A1(n_1784),
.A2(n_1588),
.B1(n_1613),
.B2(n_1614),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1789),
.A2(n_1606),
.B(n_1607),
.C(n_1597),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1784),
.A2(n_1563),
.B1(n_1340),
.B2(n_1307),
.Y(n_1802)
);

OAI211xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1770),
.A2(n_1320),
.B(n_1616),
.C(n_1592),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1795),
.Y(n_1804)
);

OAI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1790),
.A2(n_1797),
.B1(n_1792),
.B2(n_1800),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1791),
.B(n_1780),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1802),
.B(n_1782),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1796),
.A2(n_1782),
.B(n_1787),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1799),
.Y(n_1809)
);

XNOR2xp5_ASAP7_75t_L g1810 ( 
.A(n_1793),
.B(n_1774),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1794),
.B(n_1776),
.C(n_1772),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_SL g1812 ( 
.A(n_1798),
.B(n_1788),
.C(n_1778),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1803),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1786),
.C(n_1777),
.Y(n_1814)
);

NOR3x1_ASAP7_75t_SL g1815 ( 
.A(n_1813),
.B(n_1383),
.C(n_1320),
.Y(n_1815)
);

AOI211x1_ASAP7_75t_L g1816 ( 
.A1(n_1805),
.A2(n_1602),
.B(n_1592),
.C(n_1616),
.Y(n_1816)
);

OAI211xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1806),
.A2(n_1307),
.B(n_1353),
.C(n_1282),
.Y(n_1817)
);

AOI222xp33_ASAP7_75t_L g1818 ( 
.A1(n_1812),
.A2(n_1606),
.B1(n_1610),
.B2(n_1609),
.C1(n_1602),
.C2(n_1607),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1811),
.B(n_1280),
.C(n_1300),
.Y(n_1819)
);

NAND3x1_ASAP7_75t_L g1820 ( 
.A(n_1808),
.B(n_1422),
.C(n_1350),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1819),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1820),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1815),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1816),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1818),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1817),
.A2(n_1810),
.B1(n_1804),
.B2(n_1809),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1820),
.A2(n_1807),
.B1(n_1814),
.B2(n_1602),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1821),
.Y(n_1828)
);

NAND5xp2_ASAP7_75t_L g1829 ( 
.A(n_1823),
.B(n_1827),
.C(n_1824),
.D(n_1826),
.E(n_1822),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1825),
.B(n_1422),
.C(n_1280),
.Y(n_1830)
);

NAND2x1_ASAP7_75t_L g1831 ( 
.A(n_1823),
.B(n_1280),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1823),
.A2(n_1589),
.B(n_1465),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1821),
.Y(n_1833)
);

NOR3xp33_ASAP7_75t_L g1834 ( 
.A(n_1829),
.B(n_1465),
.C(n_1455),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1828),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1833),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1837),
.A2(n_1830),
.B1(n_1834),
.B2(n_1831),
.C(n_1832),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1836),
.B1(n_1300),
.B2(n_1379),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1423),
.B1(n_1588),
.B2(n_1613),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1589),
.B(n_1588),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1840),
.A2(n_1606),
.B(n_1492),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1841),
.A2(n_1480),
.B(n_1502),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1842),
.A2(n_1423),
.B1(n_1588),
.B2(n_1596),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1843),
.B(n_1467),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1845),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_R g1847 ( 
.A1(n_1846),
.A2(n_1844),
.B1(n_1472),
.B2(n_1423),
.C(n_1606),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1847),
.A2(n_1423),
.B1(n_1379),
.B2(n_1606),
.Y(n_1848)
);


endmodule