module fake_netlist_1_5345_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_16), .B(n_15), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_16), .B(n_14), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_13), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_18), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_14), .B1(n_12), .B2(n_11), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_20), .B(n_12), .Y(n_27) );
OAI22xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_11), .B1(n_3), .B2(n_4), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_11), .Y(n_29) );
OR4x1_ASAP7_75t_L g30 ( .A(n_28), .B(n_11), .C(n_5), .D(n_6), .Y(n_30) );
NAND4xp75_ASAP7_75t_L g31 ( .A(n_29), .B(n_1), .C(n_6), .D(n_7), .Y(n_31) );
OA22x2_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_29), .B1(n_7), .B2(n_11), .Y(n_32) );
NAND3xp33_ASAP7_75t_L g33 ( .A(n_31), .B(n_11), .C(n_8), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AOI221xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_10), .B1(n_11), .B2(n_33), .C(n_30), .Y(n_35) );
endmodule