module fake_jpeg_28975_n_264 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_45),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_34),
.B1(n_22),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_63),
.B1(n_77),
.B2(n_47),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_86),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_22),
.B1(n_37),
.B2(n_21),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_22),
.B1(n_26),
.B2(n_32),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_81),
.B1(n_53),
.B2(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_40),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_38),
.C(n_37),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_38),
.B1(n_20),
.B2(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_31),
.Y(n_81)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_1),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_29),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_42),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_56),
.B(n_28),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_92),
.B(n_85),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_53),
.B(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_95),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_50),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_49),
.B1(n_57),
.B2(n_42),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_85),
.B1(n_87),
.B2(n_70),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_23),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_23),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_114),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_42),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_19),
.C(n_17),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_120),
.Y(n_129)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_47),
.B1(n_65),
.B2(n_74),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_2),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_137),
.B(n_96),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_60),
.B1(n_61),
.B2(n_83),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_132),
.B1(n_138),
.B2(n_92),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_87),
.B1(n_104),
.B2(n_65),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_57),
.B1(n_44),
.B2(n_49),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_59),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_97),
.Y(n_170)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_97),
.Y(n_143)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_96),
.B1(n_107),
.B2(n_98),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_154),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_99),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_143),
.A3(n_144),
.B1(n_148),
.B2(n_127),
.C1(n_130),
.C2(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_174),
.B1(n_129),
.B2(n_146),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_99),
.C(n_94),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_167),
.C(n_74),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_163),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_122),
.B(n_116),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_103),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_102),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_17),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_147),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_103),
.C(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_138),
.B1(n_131),
.B2(n_132),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_148),
.B1(n_143),
.B2(n_117),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_3),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_195),
.B1(n_164),
.B2(n_171),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_187),
.B1(n_151),
.B2(n_173),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_169),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_155),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_196),
.C(n_167),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_130),
.B(n_127),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_188),
.B(n_187),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_126),
.B1(n_148),
.B2(n_121),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_3),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_126),
.B1(n_86),
.B2(n_143),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_86),
.C(n_4),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_207),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_177),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_152),
.B1(n_165),
.B2(n_158),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_214),
.C(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_164),
.B1(n_168),
.B2(n_160),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_211),
.B(n_186),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_180),
.B1(n_181),
.B2(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_163),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_173),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_3),
.Y(n_213)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_201),
.B1(n_205),
.B2(n_208),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_191),
.C(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_222),
.B1(n_208),
.B2(n_198),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_214),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_213),
.B(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_197),
.C(n_185),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_R g228 ( 
.A(n_207),
.B(n_178),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_228),
.B(n_190),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_215),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_227),
.B1(n_218),
.B2(n_219),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_237),
.C(n_223),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_206),
.B(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_216),
.B1(n_215),
.B2(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_238),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_190),
.C(n_204),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_227),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_247),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_219),
.C(n_189),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_234),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_237),
.C(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_251),
.C(n_247),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_230),
.B(n_6),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_253),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_5),
.C(n_7),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_257),
.A2(n_252),
.B(n_9),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_8),
.Y(n_261)
);

AOI31xp33_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_262),
.A3(n_9),
.B(n_12),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_250),
.C2(n_259),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_12),
.Y(n_264)
);


endmodule