module fake_jpeg_30431_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_13),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_47),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_29),
.B1(n_23),
.B2(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_48),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_20),
.B1(n_25),
.B2(n_35),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_77),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_84),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_82),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_43),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_86),
.B(n_91),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_116),
.B1(n_36),
.B2(n_33),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_25),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_35),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_97),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_47),
.C(n_42),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_101),
.C(n_102),
.Y(n_130)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_51),
.B1(n_45),
.B2(n_27),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_36),
.B(n_33),
.C(n_31),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_16),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_28),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_110),
.B1(n_36),
.B2(n_31),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_32),
.B1(n_19),
.B2(n_27),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_44),
.B1(n_19),
.B2(n_33),
.Y(n_123)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_18),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_51),
.B1(n_45),
.B2(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_44),
.B1(n_30),
.B2(n_34),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_51),
.B1(n_30),
.B2(n_34),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_28),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_57),
.B(n_32),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_44),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_120),
.B1(n_134),
.B2(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_133),
.B1(n_149),
.B2(n_102),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_100),
.B1(n_74),
.B2(n_75),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_30),
.B1(n_18),
.B2(n_19),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_44),
.B1(n_18),
.B2(n_22),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_44),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_116),
.B(n_99),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_22),
.B1(n_15),
.B2(n_2),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_80),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_88),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_76),
.B1(n_86),
.B2(n_84),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_157),
.B1(n_162),
.B2(n_167),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_76),
.B(n_118),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_177),
.B(n_141),
.Y(n_204)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_164),
.Y(n_186)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_94),
.B1(n_96),
.B2(n_77),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_97),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_115),
.B1(n_75),
.B2(n_89),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_174),
.B(n_175),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_100),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_173),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_89),
.C(n_109),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_178),
.C(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_125),
.B(n_100),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_100),
.B1(n_137),
.B2(n_145),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_124),
.A2(n_110),
.B(n_105),
.C(n_106),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_109),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_127),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_134),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_108),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_113),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_182),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_136),
.C(n_138),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_188),
.C(n_195),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_138),
.B1(n_136),
.B2(n_120),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_206),
.B1(n_106),
.B2(n_105),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_165),
.B1(n_121),
.B2(n_156),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_153),
.B1(n_168),
.B2(n_175),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_138),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_138),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_197),
.C(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_133),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_140),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_4),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_135),
.B1(n_140),
.B2(n_151),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_203),
.B1(n_163),
.B2(n_159),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_140),
.B1(n_74),
.B2(n_132),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_199),
.B(n_187),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_79),
.C(n_108),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_162),
.B1(n_157),
.B2(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_210),
.B1(n_213),
.B2(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_179),
.B1(n_172),
.B2(n_166),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_224),
.B1(n_225),
.B2(n_191),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_92),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_226),
.C(n_183),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_197),
.B1(n_193),
.B2(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_217),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_222),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_119),
.B1(n_132),
.B2(n_141),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_139),
.B(n_150),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_198),
.A2(n_150),
.B(n_95),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_132),
.B1(n_79),
.B2(n_92),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_98),
.C(n_1),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_227),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_98),
.B1(n_1),
.B2(n_3),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_228),
.A2(n_201),
.B1(n_200),
.B2(n_205),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_231),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_5),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_4),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_4),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_5),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_233),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_238),
.B1(n_246),
.B2(n_221),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_248),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_199),
.B1(n_188),
.B2(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_182),
.C(n_201),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_254),
.C(n_255),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_208),
.B1(n_218),
.B2(n_228),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_5),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_232),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_230),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_6),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_212),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_7),
.C(n_8),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_8),
.C(n_9),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_271),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_234),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_265),
.Y(n_289)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_225),
.B1(n_222),
.B2(n_223),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_226),
.C(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_214),
.B(n_219),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_217),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_252),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_274),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_227),
.C(n_10),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_243),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_266),
.B1(n_256),
.B2(n_255),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_282),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_239),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_258),
.Y(n_293)
);

BUFx12_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_287),
.Y(n_297)
);

AO22x1_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_247),
.B1(n_253),
.B2(n_250),
.Y(n_287)
);

AO221x1_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_250),
.B1(n_233),
.B2(n_251),
.C(n_11),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_265),
.B(n_274),
.C(n_263),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_12),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_299),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_265),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_290),
.C(n_278),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_262),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_257),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_283),
.C(n_276),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_267),
.B(n_11),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_285),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_286),
.B1(n_280),
.B2(n_283),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_267),
.C(n_9),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_292),
.C(n_12),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_309),
.A2(n_292),
.B(n_295),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_306),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_322),
.A2(n_324),
.B(n_317),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_312),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_322),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_310),
.B(n_323),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_318),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_304),
.Y(n_329)
);


endmodule