module fake_jpeg_12630_n_414 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_414);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_414;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_58),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_56),
.Y(n_134)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_22),
.B(n_0),
.CON(n_68),
.SN(n_68)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_22),
.CON(n_100),
.SN(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_72),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_78),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_42),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_79),
.Y(n_138)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_89),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_44),
.B1(n_32),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_132),
.B1(n_21),
.B2(n_17),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_22),
.B1(n_32),
.B2(n_39),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_105),
.B1(n_133),
.B2(n_137),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_101),
.B(n_125),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_45),
.B(n_39),
.C(n_30),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_21),
.C(n_17),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_46),
.A2(n_28),
.B1(n_30),
.B2(n_39),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_51),
.A2(n_42),
.B1(n_37),
.B2(n_34),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_17),
.B1(n_88),
.B2(n_5),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_118),
.A2(n_92),
.B1(n_116),
.B2(n_102),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_47),
.B(n_26),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_26),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_129),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_SL g128 ( 
.A(n_64),
.B(n_25),
.C(n_23),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_62),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_80),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_55),
.A2(n_28),
.B1(n_19),
.B2(n_16),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_67),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_136),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_2),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_88),
.A2(n_89),
.B1(n_85),
.B2(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_143),
.B(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_156),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_113),
.B(n_101),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_121),
.B(n_130),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_91),
.A2(n_53),
.B1(n_76),
.B2(n_73),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_149),
.A2(n_161),
.B1(n_169),
.B2(n_171),
.Y(n_222)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_70),
.B1(n_49),
.B2(n_21),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_174),
.B1(n_176),
.B2(n_181),
.Y(n_225)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_154),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_120),
.C(n_96),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_2),
.Y(n_168)
);

AO22x1_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_178),
.B1(n_11),
.B2(n_155),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_12),
.B1(n_4),
.B2(n_7),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_116),
.B1(n_140),
.B2(n_115),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_108),
.B1(n_139),
.B2(n_104),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_182),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_97),
.A2(n_3),
.B1(n_7),
.B2(n_9),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_142),
.B1(n_127),
.B2(n_102),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_164),
.C(n_175),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_115),
.A2(n_3),
.B1(n_7),
.B2(n_9),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_109),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_112),
.Y(n_218)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_122),
.A2(n_10),
.A3(n_11),
.B1(n_116),
.B2(n_121),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_102),
.B(n_123),
.C(n_139),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_92),
.B1(n_108),
.B2(n_130),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_221),
.B(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_195),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_209),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_110),
.B1(n_129),
.B2(n_94),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_120),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_203),
.C(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_219),
.Y(n_234)
);

OAI22x1_ASAP7_75t_SL g209 ( 
.A1(n_144),
.A2(n_96),
.B1(n_102),
.B2(n_114),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_224),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_155),
.A2(n_141),
.B1(n_98),
.B2(n_112),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_173),
.B1(n_159),
.B2(n_153),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_110),
.C(n_98),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_156),
.B(n_90),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_146),
.A2(n_104),
.B(n_90),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_177),
.B(n_150),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_164),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_185),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_160),
.B(n_182),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_246),
.B(n_253),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_143),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_238),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_165),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_245),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_161),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_251),
.C(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_170),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_214),
.B(n_200),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_247),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_178),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_248),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_167),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_158),
.C(n_184),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_178),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_178),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_196),
.A2(n_170),
.B(n_171),
.Y(n_254)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_201),
.B1(n_191),
.B2(n_205),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_170),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_222),
.B1(n_221),
.B2(n_209),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_271),
.B1(n_249),
.B2(n_241),
.Y(n_296)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_222),
.B1(n_221),
.B2(n_225),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_278),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_204),
.C(n_205),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_281),
.C(n_251),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_201),
.C(n_192),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_233),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_287),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_234),
.A2(n_253),
.B1(n_257),
.B2(n_244),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_235),
.B1(n_234),
.B2(n_232),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_233),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_240),
.B1(n_279),
.B2(n_270),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_291),
.B1(n_292),
.B2(n_304),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_256),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_248),
.B1(n_249),
.B2(n_254),
.Y(n_291)
);

A2O1A1O1Ixp25_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_226),
.B(n_246),
.C(n_231),
.D(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_293),
.B(n_307),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_265),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_309),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_260),
.A2(n_245),
.B1(n_242),
.B2(n_250),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_296),
.B1(n_314),
.B2(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_297),
.B(n_300),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_305),
.C(n_313),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_248),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_273),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_239),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_248),
.B1(n_227),
.B2(n_197),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_239),
.C(n_229),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_261),
.B(n_272),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_282),
.A2(n_275),
.B(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_308),
.B(n_293),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_265),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_228),
.B1(n_243),
.B2(n_247),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_273),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_217),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_191),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_275),
.A2(n_217),
.B1(n_211),
.B2(n_183),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_276),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_318),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_267),
.C(n_283),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_324),
.C(n_329),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_326),
.B1(n_330),
.B2(n_316),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_313),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_327),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_269),
.C(n_262),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_288),
.B1(n_266),
.B2(n_262),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_266),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_328),
.B(n_335),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_288),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_290),
.B1(n_314),
.B2(n_301),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_336),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_189),
.C(n_207),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_328),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_291),
.B1(n_289),
.B2(n_304),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_338),
.A2(n_340),
.B1(n_348),
.B2(n_353),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_290),
.B1(n_294),
.B2(n_309),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_342),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_306),
.B1(n_303),
.B2(n_302),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_322),
.A2(n_303),
.B(n_306),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_344),
.B(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_346),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_320),
.A2(n_274),
.B1(n_263),
.B2(n_278),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_329),
.A2(n_274),
.B1(n_263),
.B2(n_211),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_325),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_274),
.B(n_264),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_356),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_215),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_317),
.C(n_319),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_364),
.C(n_365),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_317),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_343),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_362),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_343),
.B(n_324),
.CI(n_334),
.CON(n_363),
.SN(n_363)
);

OAI321xp33_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_350),
.A3(n_341),
.B1(n_352),
.B2(n_351),
.C(n_353),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_323),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_327),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_337),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_367),
.C(n_370),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_326),
.Y(n_367)
);

XOR2x2_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_332),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_369),
.A2(n_354),
.B(n_342),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_336),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_349),
.C(n_338),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_369),
.Y(n_377)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_344),
.C(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_379),
.B(n_380),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_361),
.A2(n_341),
.B1(n_350),
.B2(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_381),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_368),
.A2(n_351),
.B1(n_352),
.B2(n_356),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_382),
.B(n_360),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_383),
.A2(n_189),
.B(n_264),
.Y(n_393)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_375),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_393),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_364),
.C(n_358),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_390),
.B(n_391),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_374),
.A2(n_363),
.B(n_360),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_375),
.C(n_372),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_372),
.C(n_202),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_395),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_153),
.C(n_159),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_393),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_400),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_255),
.C(n_163),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_373),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_401),
.A2(n_390),
.B(n_391),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_405),
.B(n_406),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_397),
.A2(n_389),
.B(n_387),
.Y(n_405)
);

AOI31xp67_ASAP7_75t_L g406 ( 
.A1(n_399),
.A2(n_385),
.A3(n_255),
.B(n_152),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_403),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_409),
.C(n_400),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_404),
.A2(n_394),
.B(n_398),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_407),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_410),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_411),
.B1(n_395),
.B2(n_166),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_148),
.Y(n_414)
);


endmodule