module fake_aes_6773_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AND2x4_ASAP7_75t_L g3 ( .A(n_1), .B(n_2), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_1), .B(n_2), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
AND2x4_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_5), .B(n_3), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
INVxp67_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
OAI21x1_ASAP7_75t_SL g11 ( .A1(n_9), .A2(n_6), .B(n_3), .Y(n_11) );
AOI211xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_4), .B(n_6), .C(n_3), .Y(n_12) );
NAND4xp75_ASAP7_75t_L g13 ( .A(n_12), .B(n_4), .C(n_1), .D(n_0), .Y(n_13) );
AOI222xp33_ASAP7_75t_SL g14 ( .A1(n_13), .A2(n_0), .B1(n_3), .B2(n_4), .C1(n_11), .C2(n_1), .Y(n_14) );
endmodule