module fake_jpeg_3378_n_89 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_28),
.B1(n_36),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_49),
.B1(n_0),
.B2(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_32),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_28),
.B1(n_34),
.B2(n_27),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_5),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_47),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_47),
.C(n_21),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_78),
.C(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_6),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_75),
.Y(n_81)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_47),
.B1(n_18),
.B2(n_13),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_7),
.B(n_8),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_76),
.A2(n_69),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_7),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_80),
.C(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_74),
.C(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_71),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_75),
.B(n_81),
.C(n_77),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_8),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_9),
.B(n_10),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_9),
.C(n_11),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_11),
.Y(n_89)
);


endmodule