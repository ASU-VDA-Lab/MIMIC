module fake_jpeg_25206_n_237 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_40),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_28),
.B1(n_19),
.B2(n_33),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_59),
.B1(n_22),
.B2(n_26),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_60),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_34),
.B1(n_17),
.B2(n_24),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_38),
.B1(n_37),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_76),
.B1(n_57),
.B2(n_61),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_71),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_40),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_92),
.B(n_25),
.C(n_32),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_38),
.B(n_37),
.C(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_42),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_44),
.B(n_43),
.C(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_90),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_43),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_43),
.B(n_2),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_77),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_96),
.A2(n_73),
.B(n_77),
.Y(n_142)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_21),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_29),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_76),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_89),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_83),
.B(n_92),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_128),
.B1(n_118),
.B2(n_114),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_83),
.B(n_65),
.C(n_71),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_126),
.B(n_132),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_113),
.C(n_99),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_141),
.C(n_96),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_124),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_66),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_67),
.B1(n_80),
.B2(n_68),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_66),
.C(n_15),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_74),
.B(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_134),
.Y(n_162)
);

CKINVDCx12_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_32),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_82),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_91),
.B1(n_77),
.B2(n_89),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_142),
.B(n_118),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_85),
.C(n_61),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_147),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_97),
.C(n_101),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_152),
.C(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_153),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_101),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_102),
.C(n_98),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_102),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_1),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_120),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_126),
.B(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_126),
.B1(n_125),
.B2(n_121),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_114),
.C(n_107),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_107),
.C(n_95),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_166),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_139),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_120),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_169),
.B(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_178),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_181),
.B1(n_182),
.B2(n_29),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_121),
.B1(n_143),
.B2(n_139),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_161),
.B1(n_156),
.B2(n_54),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_155),
.B(n_163),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_25),
.B(n_54),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_121),
.B1(n_136),
.B2(n_127),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_136),
.B1(n_129),
.B2(n_58),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_1),
.B(n_2),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_3),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_2),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_187),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_10),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_158),
.CI(n_145),
.CON(n_188),
.SN(n_188)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_196),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_146),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_200),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_194),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_162),
.C(n_156),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_199),
.C(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_152),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_158),
.B(n_165),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_191),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_11),
.C(n_10),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_185),
.C(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_208),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_177),
.C(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_174),
.C(n_184),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_195),
.C(n_200),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_168),
.B1(n_186),
.B2(n_20),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_196),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_192),
.B(n_195),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_220),
.B(n_3),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_168),
.B1(n_188),
.B2(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_222),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_204),
.B(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_203),
.B(n_4),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_20),
.Y(n_222)
);

NAND4xp25_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_211),
.C(n_4),
.D(n_6),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_6),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_9),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_222),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_8),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_235),
.A2(n_9),
.B1(n_234),
.B2(n_229),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g237 ( 
.A(n_236),
.Y(n_237)
);


endmodule