module fake_jpeg_32149_n_75 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_71;
wire n_52;
wire n_68;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_3),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_17),
.B1(n_15),
.B2(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_17),
.B1(n_11),
.B2(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_26),
.B(n_24),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_18),
.B1(n_12),
.B2(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_45),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_27),
.B(n_13),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_48),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_20),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_35),
.B(n_36),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_21),
.C(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_45),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_48),
.B1(n_40),
.B2(n_37),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_52),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_43),
.B1(n_38),
.B2(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_25),
.C(n_18),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_50),
.C(n_25),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_61),
.B1(n_55),
.B2(n_50),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_67),
.B(n_59),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_54),
.B(n_11),
.C(n_12),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_70),
.C(n_68),
.Y(n_73)
);

AOI221xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_9),
.B1(n_67),
.B2(n_65),
.C(n_72),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);


endmodule