module real_aes_7982_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_0), .A2(n_74), .B1(n_148), .B2(n_152), .Y(n_147) );
INVx1_ASAP7_75t_L g275 ( .A(n_1), .Y(n_275) );
AOI21xp33_ASAP7_75t_L g244 ( .A1(n_2), .A2(n_219), .B(n_245), .Y(n_244) );
AOI22xp5_ASAP7_75t_SL g529 ( .A1(n_2), .A2(n_81), .B1(n_174), .B2(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_2), .Y(n_530) );
INVx1_ASAP7_75t_L g202 ( .A(n_3), .Y(n_202) );
AND2x6_ASAP7_75t_L g224 ( .A(n_3), .B(n_200), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_3), .B(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_4), .A2(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g251 ( .A(n_5), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_6), .B(n_317), .Y(n_316) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_7), .A2(n_26), .B1(n_89), .B2(n_94), .Y(n_97) );
INVx1_ASAP7_75t_L g217 ( .A(n_8), .Y(n_217) );
INVx1_ASAP7_75t_L g331 ( .A(n_9), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_10), .A2(n_49), .B1(n_188), .B2(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_10), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_11), .B(n_232), .Y(n_304) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_12), .A2(n_27), .B1(n_89), .B2(n_90), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_13), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_14), .B(n_219), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_15), .A2(n_33), .B1(n_181), .B2(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_15), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_16), .B(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_17), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_18), .A2(n_329), .B(n_330), .C(n_332), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_19), .A2(n_81), .B1(n_173), .B2(n_174), .Y(n_80) );
INVx1_ASAP7_75t_L g173 ( .A(n_19), .Y(n_173) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_20), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_21), .B(n_249), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_22), .A2(n_53), .B1(n_131), .B2(n_134), .Y(n_130) );
INVx1_ASAP7_75t_L g265 ( .A(n_23), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_24), .A2(n_36), .B1(n_108), .B2(n_113), .Y(n_107) );
INVx2_ASAP7_75t_L g222 ( .A(n_25), .Y(n_222) );
OAI221xp5_ASAP7_75t_L g193 ( .A1(n_27), .A2(n_40), .B1(n_50), .B2(n_194), .C(n_195), .Y(n_193) );
INVxp67_ASAP7_75t_L g196 ( .A(n_27), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_28), .Y(n_100) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_29), .A2(n_224), .B(n_227), .C(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g263 ( .A(n_30), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_31), .B(n_249), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_32), .A2(n_48), .B1(n_118), .B2(n_126), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_33), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_34), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_35), .B(n_219), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_37), .A2(n_227), .B1(n_259), .B2(n_261), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_38), .Y(n_297) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_39), .Y(n_272) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_40), .A2(n_60), .B1(n_89), .B2(n_90), .Y(n_88) );
INVxp67_ASAP7_75t_L g197 ( .A(n_40), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_41), .A2(n_236), .B(n_248), .C(n_250), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_42), .Y(n_307) );
INVx1_ASAP7_75t_L g246 ( .A(n_43), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_44), .A2(n_81), .B1(n_174), .B2(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_44), .Y(n_539) );
INVx1_ASAP7_75t_L g200 ( .A(n_45), .Y(n_200) );
INVx1_ASAP7_75t_L g216 ( .A(n_46), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_47), .Y(n_194) );
INVx1_ASAP7_75t_L g188 ( .A(n_49), .Y(n_188) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_50), .A2(n_66), .B1(n_89), .B2(n_94), .Y(n_93) );
A2O1A1Ixp33_ASAP7_75t_SL g231 ( .A1(n_51), .A2(n_232), .B(n_233), .C(n_236), .Y(n_231) );
INVxp67_ASAP7_75t_L g234 ( .A(n_52), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_54), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_55), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_56), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_57), .A2(n_180), .B1(n_183), .B2(n_184), .Y(n_179) );
INVx1_ASAP7_75t_L g183 ( .A(n_57), .Y(n_183) );
INVx1_ASAP7_75t_L g300 ( .A(n_57), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_58), .A2(n_224), .B(n_227), .C(n_302), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_59), .A2(n_178), .B1(n_179), .B2(n_185), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_59), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_61), .B(n_276), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_62), .Y(n_106) );
INVx2_ASAP7_75t_L g214 ( .A(n_63), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_64), .B(n_232), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_65), .A2(n_224), .B(n_227), .C(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_67), .B(n_253), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_68), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g313 ( .A1(n_69), .A2(n_224), .B(n_227), .C(n_314), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_70), .Y(n_321) );
INVx1_ASAP7_75t_L g230 ( .A(n_71), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_72), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_73), .B(n_276), .Y(n_315) );
INVx1_ASAP7_75t_L g89 ( .A(n_75), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_76), .B(n_212), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_77), .A2(n_219), .B(n_225), .Y(n_218) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_190), .B1(n_203), .B2(n_526), .C(n_528), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_175), .Y(n_79) );
INVx1_ASAP7_75t_L g174 ( .A(n_81), .Y(n_174) );
AND2x2_ASAP7_75t_SL g81 ( .A(n_82), .B(n_136), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_116), .Y(n_82) );
OAI221xp5_ASAP7_75t_SL g83 ( .A1(n_84), .A2(n_100), .B1(n_101), .B2(n_106), .C(n_107), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x2_ASAP7_75t_L g111 ( .A(n_87), .B(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_88), .B(n_93), .Y(n_105) );
INVx2_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
AND2x2_ASAP7_75t_L g151 ( .A(n_88), .B(n_97), .Y(n_151) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
INVx1_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
AND2x2_ASAP7_75t_L g129 ( .A(n_93), .B(n_124), .Y(n_129) );
INVx1_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
AND2x4_ASAP7_75t_L g103 ( .A(n_95), .B(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g128 ( .A(n_95), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g133 ( .A(n_95), .B(n_123), .Y(n_133) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g112 ( .A(n_96), .B(n_99), .Y(n_112) );
OR2x2_ASAP7_75t_L g122 ( .A(n_96), .B(n_99), .Y(n_122) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g155 ( .A(n_97), .B(n_99), .Y(n_155) );
AND2x2_ASAP7_75t_L g160 ( .A(n_98), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g115 ( .A(n_99), .Y(n_115) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x6_ASAP7_75t_L g114 ( .A(n_105), .B(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx8_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g135 ( .A(n_112), .B(n_123), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_112), .B(n_129), .Y(n_145) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_130), .Y(n_116) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx11_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g139 ( .A(n_122), .B(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g165 ( .A(n_123), .B(n_155), .Y(n_165) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
BUFx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_156), .Y(n_136) );
OAI221xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_141), .B1(n_142), .B2(n_146), .C(n_147), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x4_ASAP7_75t_L g159 ( .A(n_151), .B(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g170 ( .A(n_151), .B(n_171), .Y(n_170) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
OAI222xp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_162), .B1(n_163), .B2(n_166), .C1(n_167), .C2(n_172), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g171 ( .A(n_161), .Y(n_171) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVxp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B1(n_186), .B2(n_187), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_179), .Y(n_185) );
INVx1_ASAP7_75t_L g184 ( .A(n_180), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_182), .A2(n_238), .B1(n_258), .B2(n_266), .Y(n_257) );
CKINVDCx14_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
AND3x1_ASAP7_75t_SL g192 ( .A(n_193), .B(n_198), .C(n_201), .Y(n_192) );
INVxp67_ASAP7_75t_L g534 ( .A(n_193), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_198), .A2(n_227), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g543 ( .A(n_198), .Y(n_543) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OAI322xp33_ASAP7_75t_L g528 ( .A1(n_199), .A2(n_246), .A3(n_529), .B1(n_531), .B2(n_535), .C1(n_538), .C2(n_540), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_199), .B(n_202), .Y(n_537) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OR2x2_ASAP7_75t_SL g542 ( .A(n_201), .B(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND4x1_ASAP7_75t_L g204 ( .A(n_205), .B(n_444), .C(n_491), .D(n_511), .Y(n_204) );
NOR3xp33_ASAP7_75t_SL g205 ( .A(n_206), .B(n_374), .C(n_399), .Y(n_205) );
OAI211xp5_ASAP7_75t_SL g206 ( .A1(n_207), .A2(n_282), .B(n_334), .C(n_364), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_254), .Y(n_208) );
INVx3_ASAP7_75t_SL g416 ( .A(n_209), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_209), .B(n_347), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_209), .B(n_269), .Y(n_497) );
AND2x2_ASAP7_75t_L g520 ( .A(n_209), .B(n_386), .Y(n_520) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_242), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g338 ( .A(n_211), .B(n_243), .Y(n_338) );
INVx3_ASAP7_75t_L g351 ( .A(n_211), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_211), .B(n_242), .Y(n_356) );
OR2x2_ASAP7_75t_L g407 ( .A(n_211), .B(n_348), .Y(n_407) );
BUFx2_ASAP7_75t_L g427 ( .A(n_211), .Y(n_427) );
AND2x2_ASAP7_75t_L g437 ( .A(n_211), .B(n_348), .Y(n_437) );
AND2x2_ASAP7_75t_L g443 ( .A(n_211), .B(n_255), .Y(n_443) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_239), .Y(n_211) );
INVx4_ASAP7_75t_L g241 ( .A(n_212), .Y(n_241) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g256 ( .A(n_213), .Y(n_256) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_214), .B(n_215), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
BUFx2_ASAP7_75t_L g325 ( .A(n_219), .Y(n_325) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_220), .B(n_224), .Y(n_266) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g228 ( .A(n_222), .Y(n_228) );
INVx1_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
INVx1_ASAP7_75t_L g229 ( .A(n_223), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_223), .Y(n_232) );
INVx3_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
INVx4_ASAP7_75t_SL g238 ( .A(n_224), .Y(n_238) );
BUFx3_ASAP7_75t_L g527 ( .A(n_224), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_230), .B(n_231), .C(n_238), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_226), .A2(n_238), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_226), .A2(n_238), .B(n_327), .C(n_328), .Y(n_326) );
INVx5_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g526 ( .A(n_227), .B(n_527), .Y(n_526) );
AND2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_228), .Y(n_237) );
BUFx3_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_235), .B(n_251), .Y(n_250) );
INVx5_ASAP7_75t_L g276 ( .A(n_235), .Y(n_276) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_237), .Y(n_318) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_240), .A2(n_244), .B(n_252), .Y(n_243) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_241), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_243), .B(n_348), .Y(n_362) );
INVx2_ASAP7_75t_L g372 ( .A(n_243), .Y(n_372) );
AND2x2_ASAP7_75t_L g385 ( .A(n_243), .B(n_351), .Y(n_385) );
OR2x2_ASAP7_75t_L g396 ( .A(n_243), .B(n_348), .Y(n_396) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_243), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g454 ( .A(n_243), .Y(n_454) );
AND2x2_ASAP7_75t_L g500 ( .A(n_243), .B(n_255), .Y(n_500) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx4_ASAP7_75t_L g317 ( .A(n_249), .Y(n_317) );
INVx1_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
INVx2_ASAP7_75t_L g311 ( .A(n_253), .Y(n_311) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_253), .A2(n_324), .B(n_333), .Y(n_323) );
INVx3_ASAP7_75t_SL g373 ( .A(n_254), .Y(n_373) );
OR2x2_ASAP7_75t_L g426 ( .A(n_254), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_269), .Y(n_254) );
INVx3_ASAP7_75t_L g348 ( .A(n_255), .Y(n_348) );
AND2x2_ASAP7_75t_L g415 ( .A(n_255), .B(n_270), .Y(n_415) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_255), .Y(n_483) );
AOI33xp33_ASAP7_75t_L g487 ( .A1(n_255), .A2(n_416), .A3(n_423), .B1(n_432), .B2(n_488), .B3(n_489), .Y(n_487) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_267), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_256), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_256), .A2(n_271), .B(n_279), .Y(n_270) );
INVx2_ASAP7_75t_L g295 ( .A(n_256), .Y(n_295) );
INVx2_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_263), .B1(n_264), .B2(n_265), .Y(n_261) );
INVx2_ASAP7_75t_L g264 ( .A(n_262), .Y(n_264) );
INVx4_ASAP7_75t_L g329 ( .A(n_262), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_266), .A2(n_272), .B(n_273), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_266), .A2(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_269), .B(n_351), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_269), .B(n_411), .C(n_413), .Y(n_410) );
AND2x2_ASAP7_75t_L g436 ( .A(n_269), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_269), .B(n_443), .Y(n_446) );
AND2x2_ASAP7_75t_L g499 ( .A(n_269), .B(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g355 ( .A(n_270), .Y(n_355) );
OR2x2_ASAP7_75t_L g449 ( .A(n_270), .B(n_348), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_277), .C(n_278), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_281), .B(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_281), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_308), .Y(n_282) );
AOI32xp33_ASAP7_75t_L g400 ( .A1(n_283), .A2(n_401), .A3(n_403), .B1(n_405), .B2(n_408), .Y(n_400) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_283), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g503 ( .A(n_283), .Y(n_503) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g435 ( .A(n_284), .B(n_419), .Y(n_435) );
AND2x2_ASAP7_75t_L g455 ( .A(n_284), .B(n_381), .Y(n_455) );
AND2x2_ASAP7_75t_L g523 ( .A(n_284), .B(n_441), .Y(n_523) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_298), .Y(n_284) );
INVx3_ASAP7_75t_L g344 ( .A(n_285), .Y(n_344) );
AND2x2_ASAP7_75t_L g358 ( .A(n_285), .B(n_342), .Y(n_358) );
OR2x2_ASAP7_75t_L g363 ( .A(n_285), .B(n_341), .Y(n_363) );
INVx1_ASAP7_75t_L g370 ( .A(n_285), .Y(n_370) );
AND2x2_ASAP7_75t_L g378 ( .A(n_285), .B(n_352), .Y(n_378) );
AND2x2_ASAP7_75t_L g380 ( .A(n_285), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_285), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g433 ( .A(n_285), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_285), .B(n_518), .Y(n_517) );
OR2x6_ASAP7_75t_L g285 ( .A(n_286), .B(n_296), .Y(n_285) );
AOI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_288), .B(n_295), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_292), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_292), .A2(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
INVx1_ASAP7_75t_L g305 ( .A(n_295), .Y(n_305) );
INVx2_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
AND2x2_ASAP7_75t_L g388 ( .A(n_298), .B(n_309), .Y(n_388) );
AND2x2_ASAP7_75t_L g398 ( .A(n_298), .B(n_323), .Y(n_398) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_305), .B(n_306), .Y(n_298) );
INVx2_ASAP7_75t_L g518 ( .A(n_308), .Y(n_518) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_322), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_309), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g359 ( .A(n_309), .Y(n_359) );
AND2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g419 ( .A(n_309), .B(n_382), .Y(n_419) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
AND2x2_ASAP7_75t_L g381 ( .A(n_310), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g432 ( .A(n_310), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_310), .B(n_342), .Y(n_464) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_320), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_319), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B(n_318), .Y(n_314) );
AND2x2_ASAP7_75t_L g343 ( .A(n_322), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g404 ( .A(n_322), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_322), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g441 ( .A(n_322), .Y(n_441) );
INVx1_ASAP7_75t_L g474 ( .A(n_322), .Y(n_474) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g352 ( .A(n_323), .B(n_342), .Y(n_352) );
INVx1_ASAP7_75t_L g382 ( .A(n_323), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_329), .B(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_339), .B1(n_345), .B2(n_352), .C(n_353), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_336), .B(n_356), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_336), .B(n_419), .Y(n_496) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_338), .B(n_386), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_338), .B(n_347), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_338), .B(n_361), .Y(n_490) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g412 ( .A(n_342), .Y(n_412) );
AND2x2_ASAP7_75t_L g387 ( .A(n_343), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g465 ( .A(n_343), .Y(n_465) );
AND2x2_ASAP7_75t_L g397 ( .A(n_344), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_344), .B(n_367), .Y(n_413) );
AND2x2_ASAP7_75t_L g477 ( .A(n_344), .B(n_403), .Y(n_477) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g386 ( .A(n_348), .B(n_355), .Y(n_386) );
AND2x2_ASAP7_75t_L g482 ( .A(n_349), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_351), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_352), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_352), .B(n_359), .Y(n_447) );
AND2x2_ASAP7_75t_L g467 ( .A(n_352), .B(n_367), .Y(n_467) );
AND2x2_ASAP7_75t_L g488 ( .A(n_352), .B(n_432), .Y(n_488) );
OAI32xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .A3(n_359), .B1(n_360), .B2(n_363), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_SL g361 ( .A(n_355), .Y(n_361) );
NAND2x1_ASAP7_75t_L g402 ( .A(n_355), .B(n_385), .Y(n_402) );
OR2x2_ASAP7_75t_L g406 ( .A(n_355), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_355), .B(n_454), .Y(n_507) );
INVx1_ASAP7_75t_L g375 ( .A(n_356), .Y(n_375) );
OAI221xp5_ASAP7_75t_SL g493 ( .A1(n_357), .A2(n_448), .B1(n_494), .B2(n_497), .C(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g365 ( .A(n_358), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g408 ( .A(n_358), .B(n_381), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_358), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g486 ( .A(n_358), .B(n_419), .Y(n_486) );
INVxp67_ASAP7_75t_L g422 ( .A(n_359), .Y(n_422) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g492 ( .A(n_361), .B(n_479), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_361), .B(n_442), .Y(n_515) );
INVx1_ASAP7_75t_L g390 ( .A(n_363), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_363), .B(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g508 ( .A(n_363), .B(n_509), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_368), .B(n_371), .Y(n_364) );
AND2x2_ASAP7_75t_L g377 ( .A(n_366), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g461 ( .A(n_370), .B(n_381), .Y(n_461) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AND2x2_ASAP7_75t_L g479 ( .A(n_372), .B(n_437), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_372), .B(n_436), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_373), .B(n_385), .Y(n_459) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_379), .C(n_389), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_410), .B1(n_414), .B2(n_417), .C(n_420), .Y(n_409) );
AOI31xp33_ASAP7_75t_L g504 ( .A1(n_375), .A2(n_505), .A3(n_506), .B(n_508), .Y(n_504) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_385), .B2(n_387), .Y(n_379) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g505 ( .A(n_385), .Y(n_505) );
INVx1_ASAP7_75t_L g468 ( .A(n_386), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_388), .A2(n_512), .B(n_514), .C(n_516), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_393), .B2(n_397), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_394), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_396), .A2(n_430), .B1(n_449), .B2(n_485), .C(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g480 ( .A(n_397), .Y(n_480) );
INVx1_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
NAND3xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_409), .C(n_424), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g450 ( .A1(n_401), .A2(n_451), .B(n_455), .Y(n_450) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_403), .B(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g510 ( .A(n_404), .Y(n_510) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g448 ( .A(n_411), .B(n_431), .Y(n_448) );
INVx1_ASAP7_75t_L g423 ( .A(n_412), .Y(n_423) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g421 ( .A(n_415), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_415), .B(n_453), .Y(n_452) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_416), .B(n_421), .C(n_422), .D(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_429), .B1(n_435), .B2(n_436), .C1(n_438), .C2(n_442), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g522 ( .A(n_426), .Y(n_522) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_438), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g498 ( .A1(n_443), .A2(n_499), .B(n_501), .Y(n_498) );
NOR4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_456), .C(n_469), .D(n_484), .Y(n_444) );
OAI221xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_447), .B1(n_448), .B2(n_449), .C(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_453), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
OAI222xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B1(n_462), .B2(n_463), .C1(n_466), .C2(n_468), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g491 ( .A1(n_461), .A2(n_492), .B(n_493), .C(n_504), .Y(n_491) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
OAI222xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_475), .B1(n_476), .B2(n_478), .C1(n_480), .C2(n_481), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_486), .A2(n_489), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI211xp5_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_519), .B(n_521), .C(n_524), .Y(n_516) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
endmodule