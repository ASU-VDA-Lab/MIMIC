module fake_jpeg_27336_n_70 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_67;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_38),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_44),
.B1(n_17),
.B2(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_7),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_15),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_16),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_61),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_60),
.C(n_57),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OAI221xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_55),
.B1(n_58),
.B2(n_56),
.C(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_24),
.Y(n_70)
);


endmodule