module fake_jpeg_27351_n_84 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

BUFx3_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx2_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_52),
.Y(n_53)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp67_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_0),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_59),
.B(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

FAx1_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_0),
.CI(n_37),
.CON(n_66),
.SN(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_58),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_75),
.A3(n_60),
.B1(n_12),
.B2(n_14),
.C(n_15),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_9),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_10),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_20),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_22),
.C(n_23),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_25),
.B(n_28),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_30),
.Y(n_84)
);


endmodule