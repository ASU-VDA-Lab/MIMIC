module fake_jpeg_11040_n_426 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_50),
.Y(n_95)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_49),
.Y(n_120)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_53),
.B(n_54),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_59),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_60),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_78),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_0),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_84),
.Y(n_130)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_0),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_61),
.C(n_59),
.Y(n_112)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_36),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_42),
.B1(n_37),
.B2(n_41),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_41),
.B1(n_42),
.B2(n_37),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_42),
.B1(n_37),
.B2(n_24),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_24),
.B1(n_34),
.B2(n_33),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_107),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_101),
.A2(n_102),
.B1(n_117),
.B2(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_29),
.B1(n_38),
.B2(n_36),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_36),
.B1(n_16),
.B2(n_38),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_46),
.B1(n_48),
.B2(n_68),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_36),
.B1(n_16),
.B2(n_3),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_62),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_57),
.B1(n_45),
.B2(n_83),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_74),
.B1(n_77),
.B2(n_66),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_136),
.B1(n_86),
.B2(n_82),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_76),
.A2(n_70),
.B1(n_73),
.B2(n_71),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_84),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_141),
.A2(n_137),
.B1(n_131),
.B2(n_115),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_142),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_112),
.B(n_135),
.C(n_133),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_146),
.B(n_150),
.C(n_154),
.Y(n_197)
);

BUFx4f_ASAP7_75t_SL g144 ( 
.A(n_103),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_69),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_79),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_149),
.B(n_164),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_1),
.Y(n_150)
);

BUFx4f_ASAP7_75t_SL g153 ( 
.A(n_103),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_156),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_157),
.A2(n_152),
.B1(n_155),
.B2(n_191),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_167),
.Y(n_213)
);

NAND2x1_ASAP7_75t_SL g162 ( 
.A(n_126),
.B(n_76),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_175),
.B(n_184),
.Y(n_201)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_124),
.B(n_80),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_175),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_5),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_5),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_100),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_176),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_65),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_62),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_179),
.Y(n_229)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_110),
.A2(n_52),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_6),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_8),
.B(n_10),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_185),
.B(n_129),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_110),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_119),
.A2(n_8),
.B(n_10),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_11),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_106),
.Y(n_187)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_188),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_140),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_11),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_12),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_127),
.A2(n_12),
.B1(n_139),
.B2(n_118),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_101),
.B1(n_139),
.B2(n_129),
.Y(n_194)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_217),
.B1(n_222),
.B2(n_236),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_195),
.B(n_205),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_219),
.C(n_153),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_148),
.B(n_177),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_200),
.A2(n_204),
.B(n_208),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_148),
.A2(n_119),
.B(n_121),
.Y(n_204)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_161),
.B(n_121),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_151),
.A2(n_108),
.B(n_140),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_209),
.A2(n_227),
.B1(n_226),
.B2(n_194),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_151),
.A2(n_108),
.B(n_140),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_237),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_215),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_170),
.A2(n_137),
.B1(n_131),
.B2(n_132),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_143),
.B(n_98),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_170),
.A2(n_132),
.B1(n_97),
.B2(n_111),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_111),
.Y(n_228)
);

NOR2x1_ASAP7_75t_R g233 ( 
.A(n_175),
.B(n_171),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_182),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_184),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_239),
.B(n_247),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_206),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_241),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_198),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_196),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_258),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_221),
.C(n_200),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_246),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_181),
.B1(n_172),
.B2(n_184),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_252),
.B1(n_261),
.B2(n_273),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_144),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_144),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_250),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_179),
.B1(n_185),
.B2(n_193),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_191),
.B1(n_160),
.B2(n_178),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_165),
.C(n_163),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_248),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_153),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_254),
.Y(n_309)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_214),
.B(n_173),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_257),
.B(n_266),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_196),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_229),
.A2(n_191),
.B1(n_145),
.B2(n_158),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_195),
.A2(n_159),
.B1(n_142),
.B2(n_183),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_189),
.B1(n_192),
.B2(n_162),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_209),
.A2(n_142),
.B1(n_188),
.B2(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_188),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_212),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_202),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_201),
.B(n_204),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_199),
.B(n_212),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_194),
.A2(n_202),
.B1(n_197),
.B2(n_210),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_233),
.A2(n_213),
.B1(n_205),
.B2(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_246),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_205),
.A2(n_213),
.B1(n_211),
.B2(n_234),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_230),
.B1(n_223),
.B2(n_235),
.Y(n_286)
);

AO22x2_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_216),
.B1(n_220),
.B2(n_199),
.Y(n_278)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_216),
.B1(n_220),
.B2(n_232),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_305),
.B1(n_242),
.B2(n_293),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_255),
.A2(n_235),
.B(n_230),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_286),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_225),
.B(n_223),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_299),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_299),
.B(n_301),
.C(n_280),
.D(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_238),
.A2(n_245),
.B1(n_249),
.B2(n_252),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_301),
.B1(n_295),
.B2(n_291),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_225),
.B(n_271),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_297),
.A2(n_304),
.B(n_282),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_271),
.B(n_244),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_307),
.C(n_292),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_249),
.A2(n_276),
.B1(n_261),
.B2(n_269),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_243),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_304),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_258),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_259),
.A2(n_271),
.B1(n_275),
.B2(n_248),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_241),
.B(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_270),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_265),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_317),
.C(n_320),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_312),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_288),
.B(n_256),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_314),
.B(n_315),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_318),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_303),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_280),
.A2(n_274),
.B1(n_268),
.B2(n_242),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_319),
.A2(n_324),
.B1(n_336),
.B2(n_278),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_274),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_321),
.A2(n_306),
.B1(n_326),
.B2(n_322),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_281),
.B(n_307),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_295),
.A2(n_289),
.B1(n_285),
.B2(n_305),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_298),
.B(n_294),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_309),
.C(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_334),
.Y(n_339)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_283),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_278),
.A2(n_284),
.B1(n_290),
.B2(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_297),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_355),
.C(n_356),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_278),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_278),
.B(n_287),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_357),
.Y(n_368)
);

OA22x2_ASAP7_75t_L g353 ( 
.A1(n_326),
.A2(n_306),
.B1(n_331),
.B2(n_323),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_306),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_310),
.B(n_313),
.C(n_315),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_324),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_322),
.C(n_311),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_311),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_364),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_354),
.B(n_316),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_361),
.B(n_369),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_311),
.C(n_332),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_373),
.C(n_377),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_338),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_327),
.C(n_328),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_374),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_346),
.B(n_329),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_375),
.B(n_337),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_335),
.C(n_319),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_341),
.C(n_358),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_348),
.C(n_353),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_376),
.A2(n_339),
.B(n_349),
.C(n_351),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_383),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_337),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_364),
.B(n_359),
.CI(n_346),
.CON(n_384),
.SN(n_384)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_362),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_386),
.B(n_390),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_368),
.A2(n_343),
.B1(n_348),
.B2(n_353),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_393),
.B1(n_363),
.B2(n_350),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_392),
.B(n_381),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_368),
.A2(n_353),
.B1(n_357),
.B2(n_347),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_365),
.C(n_362),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_403),
.C(n_391),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_385),
.A2(n_363),
.B1(n_366),
.B2(n_376),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_395),
.A2(n_391),
.B1(n_382),
.B2(n_393),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_396),
.A2(n_399),
.B(n_384),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_392),
.A2(n_378),
.B(n_377),
.Y(n_399)
);

NOR2x1p5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_380),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_401),
.B(n_387),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_402),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_360),
.C(n_352),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_404),
.B(n_408),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g406 ( 
.A1(n_398),
.A2(n_382),
.B(n_384),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_406),
.A2(n_407),
.B(n_397),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_403),
.B(n_389),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_411),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_411),
.B(n_394),
.C(n_400),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_415),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_414),
.B(n_404),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_418),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_408),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_419),
.B(n_412),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_SL g422 ( 
.A1(n_421),
.A2(n_405),
.B(n_416),
.C(n_409),
.Y(n_422)
);

OAI321xp33_ASAP7_75t_L g423 ( 
.A1(n_422),
.A2(n_388),
.A3(n_420),
.B1(n_350),
.B2(n_347),
.C(n_352),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_379),
.B(n_388),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_379),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_379),
.Y(n_426)
);


endmodule