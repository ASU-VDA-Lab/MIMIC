module fake_jpeg_19596_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_31),
.B1(n_21),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_54),
.B1(n_62),
.B2(n_41),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_21),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_38),
.C(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_31),
.B1(n_24),
.B2(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_28),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_0),
.B(n_1),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_31),
.B1(n_37),
.B2(n_36),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_47),
.B1(n_44),
.B2(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_30),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_70),
.Y(n_98)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_75),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_18),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_22),
.B1(n_32),
.B2(n_23),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_29),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_35),
.B(n_33),
.C(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_38),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_52),
.B1(n_49),
.B2(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_33),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_32),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_69),
.B1(n_90),
.B2(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_122),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_48),
.B1(n_54),
.B2(n_42),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_42),
.B1(n_41),
.B2(n_49),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_41),
.B1(n_38),
.B2(n_26),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_73),
.A2(n_38),
.B1(n_26),
.B2(n_27),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_126),
.Y(n_158)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_68),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_136),
.B(n_139),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_90),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_131),
.C(n_137),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_138),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_84),
.B(n_78),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_69),
.Y(n_137)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_84),
.B(n_74),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_79),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_147),
.Y(n_160)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_94),
.C(n_67),
.Y(n_149)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_156),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_163),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_112),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_173),
.B(n_0),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_97),
.B1(n_119),
.B2(n_99),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_179),
.B1(n_133),
.B2(n_1),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_118),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_177),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_65),
.B1(n_83),
.B2(n_86),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_172),
.B1(n_108),
.B2(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_83),
.B1(n_108),
.B2(n_110),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_138),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_16),
.C(n_13),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_140),
.B1(n_145),
.B2(n_150),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_165),
.B1(n_164),
.B2(n_179),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_130),
.C(n_137),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_184),
.C(n_191),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_131),
.C(n_134),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_134),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_190),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_171),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_145),
.C(n_89),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_178),
.B1(n_160),
.B2(n_155),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_SL g197 ( 
.A(n_162),
.B(n_27),
.C(n_26),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_155),
.B(n_159),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_27),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_2),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_13),
.C(n_3),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_167),
.C(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_214),
.B1(n_215),
.B2(n_174),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_164),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_216),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_176),
.C(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_194),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_220),
.Y(n_232)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_227),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_204),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_191),
.B(n_176),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_200),
.C(n_195),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_231),
.C(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_211),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_161),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_181),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_201),
.C(n_3),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_9),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_212),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_204),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_245),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_203),
.B(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_213),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_237),
.B(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_209),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_225),
.B(n_220),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_239),
.B(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_240),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_258),
.B(n_246),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_2),
.B(n_4),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_4),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_8),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_265),
.B(n_5),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_6),
.C(n_8),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_5),
.B(n_6),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_266),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_8),
.B(n_267),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.Y(n_271)
);


endmodule