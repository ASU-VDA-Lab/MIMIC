module fake_jpeg_1355_n_502 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_19),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_59),
.B(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_15),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_76),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_78),
.Y(n_143)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_0),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_81),
.B(n_85),
.Y(n_187)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_87),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_21),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_88),
.B(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_92),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_12),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_40),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_96),
.B(n_114),
.Y(n_170)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_37),
.Y(n_153)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_44),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_45),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_113),
.B(n_18),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_40),
.B(n_1),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_119),
.B1(n_108),
.B2(n_58),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_130),
.A2(n_156),
.B1(n_176),
.B2(n_153),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_54),
.B1(n_35),
.B2(n_48),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_131),
.A2(n_147),
.B1(n_158),
.B2(n_162),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_139),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_91),
.B(n_54),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_140),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_57),
.A2(n_54),
.B1(n_48),
.B2(n_47),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_153),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_60),
.A2(n_24),
.B1(n_41),
.B2(n_34),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_64),
.A2(n_47),
.B1(n_37),
.B2(n_55),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_157),
.A2(n_167),
.B1(n_152),
.B2(n_146),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_98),
.A2(n_49),
.B1(n_41),
.B2(n_55),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_99),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_161),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_61),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_79),
.A2(n_49),
.B1(n_18),
.B2(n_34),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_164),
.B(n_134),
.Y(n_239)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_62),
.A2(n_33),
.B(n_24),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_168),
.B(n_140),
.CI(n_158),
.CON(n_225),
.SN(n_225)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_83),
.A2(n_49),
.B1(n_33),
.B2(n_51),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_169),
.A2(n_182),
.B1(n_184),
.B2(n_188),
.Y(n_211)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_2),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_195),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_83),
.A2(n_51),
.B1(n_50),
.B2(n_22),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_84),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_84),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_69),
.B(n_2),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_116),
.A2(n_77),
.B1(n_87),
.B2(n_68),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_196),
.A2(n_101),
.B1(n_7),
.B2(n_11),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_68),
.B(n_3),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_6),
.Y(n_212)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_107),
.B1(n_63),
.B2(n_87),
.Y(n_203)
);

AOI22x1_ASAP7_75t_L g311 ( 
.A1(n_203),
.A2(n_268),
.B1(n_264),
.B2(n_240),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_143),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_217),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_223),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_218),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_212),
.B(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_101),
.B1(n_7),
.B2(n_11),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_216),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_6),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_166),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_201),
.B1(n_194),
.B2(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_230),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_226),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_142),
.B(n_170),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_148),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_228),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_144),
.B(n_195),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_145),
.A2(n_163),
.B1(n_182),
.B2(n_178),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_229),
.A2(n_234),
.B1(n_237),
.B2(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_132),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_122),
.B(n_127),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_193),
.A2(n_149),
.B1(n_180),
.B2(n_136),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_193),
.A2(n_138),
.B1(n_132),
.B2(n_155),
.Y(n_237)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_177),
.Y(n_240)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_128),
.B(n_137),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_241),
.B(n_258),
.Y(n_300)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_150),
.Y(n_242)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_177),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_243),
.B(n_256),
.Y(n_292)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_135),
.A2(n_129),
.A3(n_154),
.B1(n_131),
.B2(n_184),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_244),
.A2(n_245),
.B(n_252),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_162),
.A2(n_169),
.B(n_147),
.C(n_188),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_245),
.A2(n_212),
.B(n_244),
.C(n_207),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_246),
.A2(n_247),
.B1(n_263),
.B2(n_250),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_125),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_121),
.B(n_191),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_249),
.C(n_266),
.Y(n_299)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_138),
.B(n_197),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_124),
.Y(n_251)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_174),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_246),
.B1(n_251),
.B2(n_247),
.Y(n_297)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_179),
.A2(n_126),
.B1(n_174),
.B2(n_141),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_146),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_257),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_198),
.B(n_190),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_167),
.B(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_265),
.Y(n_307)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_141),
.Y(n_260)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_181),
.A2(n_175),
.B1(n_157),
.B2(n_140),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_261),
.A2(n_264),
.B1(n_240),
.B2(n_219),
.Y(n_317)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_139),
.Y(n_262)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_193),
.Y(n_264)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_139),
.Y(n_265)
);

INVx6_ASAP7_75t_SL g266 ( 
.A(n_176),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_175),
.B(n_199),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_248),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_157),
.A2(n_162),
.B1(n_168),
.B2(n_182),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_206),
.A2(n_211),
.B1(n_208),
.B2(n_225),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_298),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_215),
.A2(n_225),
.B1(n_267),
.B2(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_272),
.A2(n_280),
.B1(n_310),
.B2(n_314),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_204),
.A2(n_228),
.B1(n_239),
.B2(n_221),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_255),
.A2(n_221),
.B1(n_257),
.B2(n_256),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_282),
.A2(n_297),
.B1(n_303),
.B2(n_316),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_294),
.A2(n_286),
.B(n_301),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_222),
.A2(n_217),
.B1(n_212),
.B2(n_227),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_SL g305 ( 
.A(n_222),
.B(n_249),
.C(n_232),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_308),
.C(n_210),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_241),
.B(n_232),
.C(n_218),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_248),
.B(n_243),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_210),
.B(n_213),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_312),
.B(n_273),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_250),
.A2(n_254),
.B1(n_263),
.B2(n_231),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_260),
.A2(n_254),
.B1(n_219),
.B2(n_224),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_233),
.B1(n_236),
.B2(n_202),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_265),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_321),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_355),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_275),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_331),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_324),
.B(n_326),
.Y(n_370)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_220),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_325),
.A2(n_302),
.B1(n_310),
.B2(n_285),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_253),
.B(n_242),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_238),
.C(n_272),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_339),
.C(n_271),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_343),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_269),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_269),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_334),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_287),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_287),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_341),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_292),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_342),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_344),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_280),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_286),
.B(n_288),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_283),
.A2(n_298),
.B(n_301),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_299),
.B(n_281),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_314),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_351),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_281),
.B(n_276),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_347),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_276),
.B(n_313),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_301),
.A2(n_311),
.B(n_283),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_349),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_306),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_293),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_353),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_296),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_354),
.A2(n_302),
.B1(n_285),
.B2(n_271),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_296),
.B(n_317),
.Y(n_355)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_271),
.B1(n_311),
.B2(n_279),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_363),
.A2(n_364),
.B1(n_368),
.B2(n_373),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_372),
.C(n_376),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_338),
.A2(n_315),
.B1(n_278),
.B2(n_277),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_367),
.A2(n_323),
.B1(n_326),
.B2(n_345),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_350),
.A2(n_315),
.B1(n_278),
.B2(n_290),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_277),
.C(n_289),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_350),
.A2(n_290),
.B1(n_289),
.B2(n_291),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_354),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_380),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_320),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_319),
.A2(n_332),
.B1(n_341),
.B2(n_321),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_378),
.A2(n_323),
.B(n_343),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_346),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_352),
.A2(n_350),
.B1(n_336),
.B2(n_348),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_334),
.B1(n_319),
.B2(n_322),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_352),
.A2(n_326),
.B1(n_331),
.B2(n_333),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_329),
.B1(n_318),
.B2(n_337),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_389),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_L g388 ( 
.A1(n_359),
.A2(n_324),
.B(n_344),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_388),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_362),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_377),
.Y(n_390)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_392),
.A2(n_393),
.B(n_396),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_370),
.A2(n_330),
.B(n_319),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_356),
.A2(n_319),
.B(n_343),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_320),
.C(n_339),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_374),
.C(n_365),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_357),
.B(n_335),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_357),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_356),
.Y(n_401)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_358),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_402),
.Y(n_419)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_358),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_404),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_405),
.A2(n_407),
.B1(n_380),
.B2(n_360),
.Y(n_429)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_378),
.A2(n_324),
.B(n_329),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_408),
.B(n_410),
.Y(n_412)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_379),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_409),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_385),
.A2(n_355),
.B(n_351),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_369),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_411),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_417),
.C(n_422),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_374),
.C(n_372),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_400),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_356),
.C(n_382),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_369),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_424),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_384),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_399),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_381),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_393),
.Y(n_447)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_434),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_433),
.A2(n_405),
.B1(n_394),
.B2(n_411),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_439),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_449),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_428),
.A2(n_389),
.B1(n_402),
.B2(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_399),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_441),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_433),
.A2(n_394),
.B1(n_387),
.B2(n_395),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_427),
.A2(n_386),
.B1(n_363),
.B2(n_387),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_442),
.A2(n_448),
.B1(n_450),
.B2(n_421),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_415),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_412),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_447),
.B(n_430),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_432),
.A2(n_418),
.B1(n_381),
.B2(n_421),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_396),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_418),
.A2(n_410),
.B1(n_360),
.B2(n_401),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_450),
.A2(n_415),
.B(n_396),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_454),
.A2(n_442),
.B(n_396),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_449),
.Y(n_473)
);

AOI322xp5_ASAP7_75t_L g459 ( 
.A1(n_439),
.A2(n_392),
.A3(n_375),
.B1(n_429),
.B2(n_424),
.C1(n_385),
.C2(n_431),
.Y(n_459)
);

OAI221xp5_ASAP7_75t_L g471 ( 
.A1(n_459),
.A2(n_440),
.B1(n_444),
.B2(n_413),
.C(n_425),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_417),
.C(n_414),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_446),
.C(n_422),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_SL g468 ( 
.A1(n_463),
.A2(n_412),
.B(n_437),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_462),
.A2(n_435),
.B1(n_441),
.B2(n_448),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_464),
.A2(n_472),
.B1(n_460),
.B2(n_452),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_465),
.B(n_473),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_455),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_468),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_460),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_474),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_470),
.B(n_471),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_453),
.A2(n_373),
.B1(n_368),
.B2(n_425),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_453),
.A2(n_371),
.B1(n_367),
.B2(n_391),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_466),
.A2(n_456),
.B1(n_455),
.B2(n_457),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g484 ( 
.A1(n_475),
.A2(n_466),
.B(n_471),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_461),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_436),
.Y(n_488)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_482),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_465),
.A2(n_454),
.B(n_457),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_483),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_486),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_436),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_485),
.B(n_488),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_473),
.Y(n_489)
);

NAND4xp25_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_480),
.C(n_479),
.D(n_481),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_491),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_475),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_486),
.C(n_469),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_496),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_451),
.C(n_458),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_491),
.B(n_490),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_499),
.A2(n_497),
.B(n_451),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_500),
.A2(n_416),
.B(n_406),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_416),
.B1(n_409),
.B2(n_403),
.Y(n_502)
);


endmodule