module real_jpeg_32651_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_0),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_0),
.B(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_2),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_98),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_6),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_7),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_7),
.B(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_12),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_12),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_12),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_13),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_13),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_13),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_13),
.B(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_140),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_93),
.B(n_139),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_60),
.Y(n_17)
);

NAND2xp33_ASAP7_75t_L g139 ( 
.A(n_18),
.B(n_60),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.C(n_50),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_19),
.A2(n_20),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_33),
.C(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_27),
.Y(n_179)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_32),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_35),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_41),
.A2(n_50),
.B1(n_51),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_45),
.Y(n_151)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_53),
.B(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_54),
.Y(n_184)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_78),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_R g144 ( 
.A(n_64),
.B(n_68),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_64),
.B(n_188),
.C(n_189),
.Y(n_187)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_69),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_143),
.C(n_144),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_79),
.B(n_81),
.C(n_88),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

AOI21x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_110),
.B(n_138),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.C(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_131),
.B(n_137),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_126),
.B(n_130),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_117),
.Y(n_130)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_123),
.Y(n_132)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_190),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_145),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_167),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_166),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_165),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_158),
.B1(n_159),
.B2(n_164),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_180),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_176),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);


endmodule