module fake_jpeg_2811_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_3),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_60),
.Y(n_174)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_61),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_104),
.Y(n_136)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_17),
.B(n_16),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_66),
.A2(n_115),
.B(n_30),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_67),
.B(n_92),
.Y(n_157)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_68),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_69),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_73),
.Y(n_178)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_75),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_79),
.Y(n_183)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_36),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_84),
.B(n_111),
.Y(n_139)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

CKINVDCx10_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_25),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_94),
.Y(n_186)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_32),
.B(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_106),
.Y(n_130)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_103),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_20),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_32),
.B(n_13),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_113),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_12),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_112),
.Y(n_195)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_117),
.Y(n_143)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_20),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_120),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_37),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_121),
.Y(n_172)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_125),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_92),
.A2(n_26),
.B1(n_53),
.B2(n_47),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_131),
.A2(n_141),
.B1(n_148),
.B2(n_164),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_135),
.B(n_161),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_58),
.A2(n_26),
.B1(n_39),
.B2(n_47),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_109),
.B1(n_118),
.B2(n_64),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_144),
.A2(n_155),
.B1(n_197),
.B2(n_182),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_88),
.B(n_54),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_147),
.B(n_181),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_62),
.A2(n_42),
.B1(n_39),
.B2(n_34),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_72),
.A2(n_38),
.B1(n_51),
.B2(n_27),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_149),
.A2(n_173),
.B1(n_189),
.B2(n_205),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_96),
.A2(n_38),
.B1(n_42),
.B2(n_34),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_151),
.A2(n_194),
.B1(n_195),
.B2(n_204),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_59),
.B(n_51),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_171),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_70),
.B(n_29),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_162),
.A2(n_175),
.B(n_214),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_105),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_77),
.A2(n_50),
.B1(n_33),
.B2(n_31),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_166),
.A2(n_180),
.B1(n_149),
.B2(n_144),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_61),
.B(n_50),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_81),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_90),
.A2(n_23),
.B(n_43),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_87),
.A2(n_94),
.B1(n_89),
.B2(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_121),
.B(n_0),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_79),
.B(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_188),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_76),
.B(n_1),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_9),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_101),
.B(n_2),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_125),
.B(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_193),
.B(n_209),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_122),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_194)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_93),
.B(n_6),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_206),
.B(n_214),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_11),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_100),
.B(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_213),
.B(n_165),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_63),
.B(n_7),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_136),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_215),
.A2(n_244),
.B1(n_256),
.B2(n_258),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_216),
.A2(n_222),
.B(n_227),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_10),
.B1(n_157),
.B2(n_161),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_217),
.A2(n_224),
.B1(n_252),
.B2(n_274),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_218),
.Y(n_326)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

INVx3_ASAP7_75t_SL g221 ( 
.A(n_177),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_221),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_128),
.A2(n_151),
.B1(n_170),
.B2(n_186),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_144),
.A2(n_140),
.B1(n_199),
.B2(n_135),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_226),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_174),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_150),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_230),
.Y(n_294)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_229),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_146),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_140),
.A2(n_146),
.B1(n_143),
.B2(n_156),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_231),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_292)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_145),
.B(n_154),
.C(n_168),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_264),
.Y(n_291)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_236),
.Y(n_334)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_174),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_239),
.Y(n_317)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_138),
.Y(n_240)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_157),
.A2(n_139),
.B1(n_193),
.B2(n_130),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_245),
.B(n_254),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_134),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_271),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_137),
.A2(n_169),
.B(n_208),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_249),
.A2(n_265),
.B(n_276),
.C(n_269),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_194),
.A2(n_186),
.B1(n_152),
.B2(n_201),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_250),
.A2(n_257),
.B1(n_279),
.B2(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_251),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_200),
.B(n_179),
.Y(n_254)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_142),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_129),
.A2(n_158),
.B1(n_191),
.B2(n_133),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_152),
.A2(n_172),
.B1(n_158),
.B2(n_129),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_132),
.A2(n_182),
.B1(n_197),
.B2(n_155),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_133),
.A2(n_191),
.B1(n_207),
.B2(n_202),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_259),
.A2(n_261),
.B1(n_272),
.B2(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_190),
.A2(n_210),
.B1(n_203),
.B2(n_192),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_142),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_192),
.C(n_210),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_177),
.A2(n_178),
.B(n_203),
.C(n_190),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_137),
.A2(n_126),
.B1(n_178),
.B2(n_211),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_126),
.A2(n_211),
.B1(n_198),
.B2(n_204),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_176),
.A2(n_167),
.B1(n_127),
.B2(n_196),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_183),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_269),
.B(n_273),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_127),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_196),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_165),
.A2(n_167),
.B1(n_159),
.B2(n_187),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_159),
.A2(n_206),
.B1(n_157),
.B2(n_161),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_187),
.A2(n_175),
.B(n_146),
.C(n_135),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_153),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_277),
.Y(n_313)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_153),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_157),
.A2(n_136),
.B1(n_173),
.B2(n_135),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_214),
.A2(n_135),
.B1(n_63),
.B2(n_157),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_132),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_150),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_285),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_214),
.B(n_135),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.C(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_206),
.B(n_214),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_253),
.Y(n_293)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_127),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_288),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_135),
.B(n_214),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_284),
.A2(n_253),
.B1(n_252),
.B2(n_227),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_311),
.B1(n_322),
.B2(n_323),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_293),
.B(n_291),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_295),
.B(n_272),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_300),
.Y(n_337)
);

AO21x2_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_224),
.B(n_242),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_298),
.A2(n_306),
.B1(n_232),
.B2(n_234),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_216),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_241),
.A2(n_251),
.B1(n_249),
.B2(n_229),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_217),
.A2(n_239),
.B1(n_227),
.B2(n_247),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_239),
.A2(n_276),
.B1(n_243),
.B2(n_254),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_225),
.A2(n_256),
.B1(n_286),
.B2(n_254),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_269),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_221),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_286),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_330),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_304),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_223),
.B(n_264),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_265),
.A2(n_246),
.B1(n_238),
.B2(n_237),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_333),
.B1(n_290),
.B2(n_323),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_219),
.A2(n_220),
.B1(n_235),
.B2(n_260),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_218),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_339),
.B(n_342),
.Y(n_377)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_288),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_315),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_343),
.B(n_353),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_R g344 ( 
.A(n_322),
.B(n_270),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_357),
.B(n_374),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_366),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_285),
.C(n_234),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_352),
.C(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_349),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_281),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_354),
.Y(n_384)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_240),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_314),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_355),
.A2(n_298),
.B1(n_331),
.B2(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

OR2x2_ASAP7_75t_SL g357 ( 
.A(n_307),
.B(n_278),
.Y(n_357)
);

AOI21xp33_ASAP7_75t_L g358 ( 
.A1(n_330),
.A2(n_236),
.B(n_282),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_335),
.A2(n_255),
.B1(n_262),
.B2(n_233),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_293),
.B(n_300),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_361),
.B(n_363),
.Y(n_397)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_309),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_365),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_295),
.B(n_317),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_367),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_329),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_326),
.Y(n_368)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_312),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g370 ( 
.A(n_312),
.B(n_304),
.CI(n_298),
.CON(n_370),
.SN(n_370)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_333),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_310),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_371),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_310),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_372),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_316),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_373),
.A2(n_319),
.B1(n_328),
.B2(n_324),
.Y(n_408)
);

AOI31xp33_ASAP7_75t_L g374 ( 
.A1(n_304),
.A2(n_298),
.A3(n_297),
.B(n_301),
.Y(n_374)
);

AO21x1_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_367),
.B(n_340),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_378),
.A2(n_390),
.B1(n_408),
.B2(n_336),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_388),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_371),
.Y(n_435)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_324),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_398),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_387),
.B(n_393),
.Y(n_429)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_400),
.Y(n_421)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_386),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_416),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_390),
.A2(n_378),
.B1(n_384),
.B2(n_354),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_389),
.B1(n_402),
.B2(n_400),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_384),
.A2(n_340),
.B1(n_365),
.B2(n_375),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_430),
.B1(n_387),
.B2(n_404),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_350),
.Y(n_415)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_407),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_407),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_417),
.A2(n_427),
.B1(n_429),
.B2(n_433),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_346),
.C(n_352),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_420),
.C(n_425),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_353),
.B1(n_370),
.B2(n_338),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_419),
.A2(n_422),
.B1(n_431),
.B2(n_393),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_338),
.C(n_405),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_397),
.A2(n_370),
.B1(n_337),
.B2(n_361),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_364),
.Y(n_424)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_342),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_343),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_401),
.A2(n_344),
.B1(n_369),
.B2(n_292),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_401),
.A2(n_373),
.B1(n_372),
.B2(n_339),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_357),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_398),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_377),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_382),
.B(n_368),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_434),
.B(n_406),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_399),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_379),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_379),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_321),
.C(n_308),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_412),
.C(n_418),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_440),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_441),
.B(n_443),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_433),
.B(n_399),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_442),
.B(n_447),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_455),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_446),
.A2(n_449),
.B1(n_421),
.B2(n_409),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_392),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_419),
.A2(n_404),
.B1(n_387),
.B2(n_395),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_392),
.Y(n_450)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_415),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_454),
.B(n_411),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_423),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_456),
.A2(n_458),
.B1(n_463),
.B2(n_421),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_430),
.A2(n_396),
.B1(n_389),
.B2(n_381),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_422),
.B(n_381),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_460),
.A2(n_436),
.B(n_299),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_416),
.B(n_376),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_462),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_417),
.B(n_376),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_380),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_443),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_420),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_472),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_451),
.A2(n_429),
.B1(n_435),
.B2(n_413),
.Y(n_469)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_438),
.C(n_435),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_473),
.C(n_461),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_414),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_426),
.C(n_432),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_431),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_484),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_475),
.A2(n_478),
.B1(n_462),
.B2(n_448),
.Y(n_496)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_446),
.A2(n_410),
.B1(n_437),
.B2(n_411),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_456),
.A2(n_436),
.B1(n_409),
.B2(n_380),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_448),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_483),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_494),
.C(n_499),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_466),
.B(n_440),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_486),
.B(n_489),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_468),
.B(n_439),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_441),
.C(n_463),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_470),
.C(n_481),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_467),
.B(n_461),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_482),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_480),
.B(n_449),
.Y(n_494)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_496),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_497),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_458),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_501),
.B(n_502),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_465),
.C(n_473),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_491),
.Y(n_504)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_504),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_487),
.A2(n_469),
.B1(n_491),
.B2(n_493),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_505),
.A2(n_493),
.B1(n_471),
.B2(n_478),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_509),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_485),
.C(n_465),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_498),
.C(n_499),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_487),
.A2(n_442),
.B(n_474),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_479),
.B1(n_460),
.B2(n_475),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_497),
.Y(n_512)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_512),
.Y(n_521)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_513),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_500),
.A2(n_453),
.B1(n_454),
.B2(n_459),
.Y(n_514)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_490),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_515),
.B(n_517),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_504),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_471),
.B(n_518),
.Y(n_524)
);

NOR2x1_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_459),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_522),
.A2(n_519),
.B(n_452),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_496),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_508),
.C(n_502),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_526),
.B(n_517),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_528),
.A2(n_530),
.B(n_531),
.Y(n_532)
);

AO21x1_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_523),
.B(n_521),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_527),
.A2(n_503),
.B1(n_516),
.B2(n_507),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_533),
.B(n_534),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_530),
.A2(n_522),
.B(n_525),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_532),
.Y(n_536)
);

AOI32xp33_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_524),
.A3(n_526),
.B1(n_457),
.B2(n_514),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_535),
.B(n_509),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_510),
.Y(n_539)
);


endmodule