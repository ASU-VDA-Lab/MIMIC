module fake_jpeg_18132_n_288 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2x1_ASAP7_75t_SL g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_32),
.B1(n_18),
.B2(n_23),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_57),
.B1(n_22),
.B2(n_20),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_32),
.B1(n_18),
.B2(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_27),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_61),
.B(n_70),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_33),
.B1(n_37),
.B2(n_36),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_62),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_14),
.B1(n_25),
.B2(n_31),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_25),
.B1(n_14),
.B2(n_31),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_65),
.Y(n_127)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_74),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_101),
.B1(n_92),
.B2(n_60),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_28),
.B(n_21),
.C(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_69),
.B(n_71),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_15),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_15),
.B1(n_20),
.B2(n_22),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_92),
.Y(n_114)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_79),
.B1(n_87),
.B2(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_19),
.B1(n_16),
.B2(n_26),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_28),
.B1(n_21),
.B2(n_13),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_38),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_44),
.C(n_43),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_96),
.C(n_99),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_21),
.B1(n_13),
.B2(n_12),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_98),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_44),
.C(n_43),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_47),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_41),
.B1(n_26),
.B2(n_40),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_66),
.B1(n_76),
.B2(n_65),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_111),
.B1(n_117),
.B2(n_126),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_44),
.A3(n_43),
.B1(n_42),
.B2(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_70),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_42),
.B1(n_38),
.B2(n_40),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_61),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_42),
.B1(n_19),
.B2(n_16),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_125),
.B1(n_3),
.B2(n_4),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_0),
.B(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_2),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_61),
.A2(n_19),
.B1(n_16),
.B2(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_99),
.C(n_68),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_144),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_79),
.B1(n_77),
.B2(n_88),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_104),
.B1(n_115),
.B2(n_124),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_154),
.B1(n_156),
.B2(n_133),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_60),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_138),
.B(n_145),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_70),
.B1(n_94),
.B2(n_68),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_82),
.B1(n_89),
.B2(n_98),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_147),
.B1(n_125),
.B2(n_110),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_150),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_67),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_26),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_148),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_83),
.B1(n_85),
.B2(n_12),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_3),
.B(n_4),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_27),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_159),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_27),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_19),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_73),
.C(n_16),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_114),
.B(n_3),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_103),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_3),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_182),
.B1(n_129),
.B2(n_140),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_141),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_180),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_121),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_183),
.B(n_181),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_179),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_102),
.B(n_118),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_158),
.B1(n_137),
.B2(n_126),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_180),
.B1(n_140),
.B2(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_192),
.B1(n_199),
.B2(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_112),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_200),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_135),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_193),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_178),
.B1(n_174),
.B2(n_186),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_210),
.B1(n_182),
.B2(n_130),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_143),
.B(n_116),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_170),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_209),
.B1(n_181),
.B2(n_164),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_204),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_177),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_144),
.C(n_152),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_208),
.C(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_167),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_120),
.C(n_156),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_154),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_154),
.B1(n_107),
.B2(n_131),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_194),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_212),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_196),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_179),
.B1(n_161),
.B2(n_163),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_226),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_201),
.B1(n_206),
.B2(n_190),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_161),
.B1(n_163),
.B2(n_176),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_221),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_184),
.B1(n_162),
.B2(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_184),
.C(n_169),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_225),
.C(n_229),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_131),
.C(n_123),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_171),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_228),
.B1(n_198),
.B2(n_187),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_115),
.B1(n_104),
.B2(n_109),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_112),
.C(n_109),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_210),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_203),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_212),
.B1(n_228),
.B2(n_214),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_203),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_236),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_240),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_196),
.CI(n_198),
.CON(n_241),
.SN(n_241)
);

NAND3xp33_ASAP7_75t_SL g248 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

OAI22x1_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_160),
.B1(n_5),
.B2(n_6),
.Y(n_255)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_229),
.C(n_217),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_224),
.C(n_227),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_224),
.B(n_197),
.C(n_202),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_237),
.B(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_197),
.C(n_104),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_243),
.B1(n_5),
.B2(n_6),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_261),
.A2(n_258),
.B1(n_251),
.B2(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_266),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_267),
.B(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_230),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_241),
.B(n_242),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_4),
.B(n_6),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_272),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_250),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_231),
.B1(n_248),
.B2(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_257),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_270),
.B(n_7),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_262),
.B1(n_260),
.B2(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_273),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_271),
.B(n_6),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_279),
.Y(n_284)
);

AOI31xp33_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_4),
.A3(n_7),
.B(n_9),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_283),
.B(n_9),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_286),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_7),
.Y(n_288)
);


endmodule