module fake_jpeg_14959_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_28),
.B1(n_21),
.B2(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_48),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_16),
.C(n_19),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_24),
.B(n_32),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_20),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_26),
.B(n_25),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_21),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_18),
.B1(n_28),
.B2(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_66),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_41),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_68),
.C(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_21),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_31),
.B(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_77),
.B1(n_41),
.B2(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_81),
.Y(n_88)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_34),
.B1(n_31),
.B2(n_23),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_25),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_47),
.B1(n_56),
.B2(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_102),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_96),
.B1(n_99),
.B2(n_0),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_67),
.B1(n_74),
.B2(n_84),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_78),
.B(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_70),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_56),
.C(n_26),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_104),
.C(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_53),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_47),
.B1(n_56),
.B2(n_23),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_111),
.B1(n_29),
.B2(n_33),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_66),
.B(n_26),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_29),
.B(n_26),
.C(n_17),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_86),
.B1(n_60),
.B2(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_138),
.B(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_130),
.B1(n_3),
.B2(n_4),
.Y(n_169)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_85),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_122),
.B(n_124),
.C(n_129),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_123),
.B(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_76),
.B1(n_33),
.B2(n_64),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_142),
.B1(n_96),
.B2(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_0),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_64),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_29),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_99),
.C(n_113),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_136),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_100),
.B(n_109),
.C(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_89),
.B(n_100),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_147),
.B(n_161),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_169),
.B1(n_171),
.B2(n_138),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_148),
.A2(n_154),
.B(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_151),
.Y(n_196)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_98),
.B(n_110),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_98),
.B(n_101),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_101),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.C(n_162),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_124),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_97),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_126),
.B1(n_116),
.B2(n_133),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_105),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_99),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_3),
.Y(n_165)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_11),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_132),
.C(n_141),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_5),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_120),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_161),
.B(n_158),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_191),
.B1(n_165),
.B2(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_148),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_127),
.B1(n_143),
.B2(n_137),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_144),
.B1(n_160),
.B2(n_147),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_10),
.C(n_6),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_203),
.C(n_170),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_5),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_5),
.Y(n_193)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_199),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_157),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_7),
.C(n_8),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_171),
.B1(n_177),
.B2(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_145),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_155),
.C(n_154),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_223),
.C(n_224),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_197),
.B1(n_195),
.B2(n_202),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_220),
.A2(n_225),
.B(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_145),
.C(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_231),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_233),
.B1(n_208),
.B2(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_182),
.C(n_186),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_177),
.B1(n_185),
.B2(n_178),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_188),
.C(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_238),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_198),
.B1(n_179),
.B2(n_178),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_213),
.B1(n_208),
.B2(n_218),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_198),
.C(n_192),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_179),
.C(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_240),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_168),
.C(n_149),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_168),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_243),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_214),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_212),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_255),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_252),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_217),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_150),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_209),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_232),
.B(n_221),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_255),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_227),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_147),
.Y(n_277)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_231),
.B(n_242),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_246),
.B(n_219),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_227),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_267),
.C(n_5),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.C(n_243),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_153),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_219),
.B1(n_222),
.B2(n_206),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_237),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_281),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_282),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_190),
.C(n_146),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_190),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_290),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_268),
.B(n_267),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_289),
.A2(n_279),
.B(n_280),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_274),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

OA21x2_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_8),
.B(n_12),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_284),
.C(n_285),
.Y(n_296)
);

AOI321xp33_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_298),
.A3(n_294),
.B1(n_14),
.B2(n_15),
.C(n_12),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_297),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_15),
.Y(n_302)
);


endmodule