module fake_jpeg_24953_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_21),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_8),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_18),
.A2(n_19),
.B(n_14),
.C(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx12_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_13),
.B(n_9),
.C(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_2),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_12),
.B1(n_14),
.B2(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_20),
.B(n_12),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_36),
.C(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_43),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_43),
.B(n_41),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_48),
.A3(n_42),
.B1(n_38),
.B2(n_34),
.C1(n_39),
.C2(n_32),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_34),
.B(n_6),
.Y(n_51)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_7),
.B(n_16),
.Y(n_52)
);


endmodule