module fake_netlist_1_5183_n_726 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_726);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_726;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx10_ASAP7_75t_L g92 ( .A(n_84), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_24), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_55), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_77), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_47), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_83), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_71), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_68), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_80), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_20), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_56), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_90), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_72), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_33), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_82), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_87), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_1), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_91), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_46), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_66), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_67), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_74), .Y(n_118) );
BUFx5_ASAP7_75t_L g119 ( .A(n_70), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_21), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_88), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_3), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_8), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_54), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_30), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_51), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_95), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_96), .A2(n_40), .B(n_85), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_119), .Y(n_131) );
BUFx8_ASAP7_75t_L g132 ( .A(n_125), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_111), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_96), .B(n_41), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_119), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_101), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_119), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_115), .A2(n_0), .B1(n_4), .B2(n_5), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_122), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_122), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_92), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_100), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_119), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_94), .B(n_97), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_143), .B(n_118), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_137), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
NOR2xp33_ASAP7_75t_SL g153 ( .A(n_135), .B(n_126), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_143), .B(n_102), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_133), .B(n_149), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g158 ( .A1(n_146), .A2(n_113), .B1(n_121), .B2(n_127), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_135), .B(n_119), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_143), .B(n_92), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_132), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_142), .B(n_92), .Y(n_163) );
AND3x2_ASAP7_75t_L g164 ( .A(n_132), .B(n_103), .C(n_104), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_128), .B(n_108), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_133), .A2(n_105), .B1(n_112), .B2(n_107), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_135), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_149), .B(n_108), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_144), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_145), .B(n_107), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_132), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_134), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_139), .A2(n_113), .B1(n_121), .B2(n_124), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_148), .B(n_109), .Y(n_183) );
CKINVDCx6p67_ASAP7_75t_R g184 ( .A(n_135), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_161), .B(n_116), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_168), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g187 ( .A(n_155), .B(n_141), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_176), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_176), .A2(n_135), .B1(n_141), .B2(n_147), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
INVxp67_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_177), .B(n_154), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_168), .B(n_130), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_153), .B(n_116), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_163), .A2(n_140), .B1(n_124), .B2(n_147), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_169), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_169), .B(n_99), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_153), .B(n_106), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_180), .A2(n_110), .B1(n_109), .B2(n_117), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_162), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_169), .B(n_183), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_169), .A2(n_130), .B1(n_110), .B2(n_120), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_150), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_182), .B(n_7), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_171), .B(n_130), .Y(n_212) );
AND2x6_ASAP7_75t_SL g213 ( .A(n_183), .B(n_9), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_168), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_179), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_180), .A2(n_101), .B1(n_11), .B2(n_12), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_156), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_173), .B(n_101), .Y(n_218) );
OAI22xp5_ASAP7_75t_SL g219 ( .A1(n_158), .A2(n_101), .B1(n_11), .B2(n_12), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_184), .A2(n_10), .B1(n_13), .B2(n_14), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_172), .B(n_45), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_184), .B(n_10), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_156), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_166), .B(n_13), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
AOI22x1_ASAP7_75t_L g226 ( .A1(n_194), .A2(n_181), .B1(n_178), .B2(n_167), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_188), .B(n_164), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_196), .B(n_174), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_191), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_209), .A2(n_160), .B(n_167), .Y(n_230) );
NOR3xp33_ASAP7_75t_L g231 ( .A(n_219), .B(n_166), .C(n_174), .Y(n_231) );
NOR2xp67_ASAP7_75t_L g232 ( .A(n_215), .B(n_14), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_192), .B(n_172), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_212), .A2(n_172), .B(n_181), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_SL g236 ( .A1(n_193), .A2(n_181), .B(n_178), .C(n_175), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_188), .B(n_178), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_205), .A2(n_175), .B(n_170), .C(n_165), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_205), .A2(n_175), .B1(n_170), .B2(n_165), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_189), .B(n_15), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_214), .A2(n_170), .B(n_165), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_211), .B(n_15), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_210), .B(n_16), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_211), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_214), .A2(n_157), .B(n_151), .Y(n_245) );
AOI21x1_ASAP7_75t_L g246 ( .A1(n_195), .A2(n_157), .B(n_151), .Y(n_246) );
BUFx12f_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_198), .A2(n_206), .B1(n_191), .B2(n_207), .Y(n_248) );
AO32x2_ASAP7_75t_L g249 ( .A1(n_220), .A2(n_16), .A3(n_17), .B1(n_151), .B2(n_19), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
OR2x6_ASAP7_75t_SL g251 ( .A(n_204), .B(n_17), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_198), .B(n_18), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_221), .A2(n_157), .B(n_23), .C(n_25), .Y(n_253) );
CKINVDCx10_ASAP7_75t_R g254 ( .A(n_213), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_185), .B(n_151), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_194), .B(n_218), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_238), .A2(n_200), .B(n_224), .C(n_206), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_238), .A2(n_187), .B(n_207), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_250), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_243), .A2(n_187), .B(n_208), .C(n_202), .Y(n_262) );
OAI21xp33_ASAP7_75t_L g263 ( .A1(n_243), .A2(n_202), .B(n_197), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_236), .A2(n_194), .B(n_208), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_244), .B(n_210), .Y(n_265) );
CKINVDCx11_ASAP7_75t_R g266 ( .A(n_247), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_235), .A2(n_203), .B(n_217), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_242), .B(n_199), .Y(n_268) );
BUFx8_ASAP7_75t_L g269 ( .A(n_225), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_227), .Y(n_270) );
OAI21xp33_ASAP7_75t_L g271 ( .A1(n_240), .A2(n_222), .B(n_190), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_231), .A2(n_216), .B(n_222), .C(n_217), .Y(n_273) );
AO32x2_ASAP7_75t_L g274 ( .A1(n_248), .A2(n_223), .A3(n_203), .B1(n_201), .B2(n_151), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_229), .A2(n_201), .B(n_223), .C(n_27), .Y(n_275) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_230), .A2(n_151), .B(n_26), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_229), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_226), .A2(n_22), .B(n_28), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_258), .A2(n_252), .B(n_245), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_263), .A2(n_232), .B1(n_233), .B2(n_256), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_272), .B(n_255), .Y(n_281) );
CKINVDCx11_ASAP7_75t_R g282 ( .A(n_266), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_277), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_261), .B(n_250), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_274), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_260), .B(n_233), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_261), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_269), .B(n_255), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_268), .B(n_239), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_264), .A2(n_246), .B(n_239), .Y(n_290) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_264), .A2(n_241), .B(n_253), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_257), .A2(n_253), .B(n_255), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_259), .B(n_249), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_270), .B(n_234), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_269), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_265), .B(n_251), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
BUFx8_ASAP7_75t_SL g300 ( .A(n_273), .Y(n_300) );
OA21x2_ASAP7_75t_L g301 ( .A1(n_257), .A2(n_249), .B(n_255), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_275), .A2(n_249), .B(n_234), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_283), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_289), .B(n_262), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_285), .Y(n_305) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_289), .A2(n_275), .B(n_267), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_283), .B(n_276), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_293), .B(n_249), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_293), .B(n_267), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_292), .A2(n_276), .B(n_271), .Y(n_315) );
OA21x2_ASAP7_75t_L g316 ( .A1(n_302), .A2(n_234), .B(n_31), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_292), .A2(n_234), .B(n_32), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_302), .A2(n_29), .B(n_34), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_302), .A2(n_35), .B(n_36), .Y(n_324) );
BUFx4f_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_301), .B(n_38), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_254), .B1(n_42), .B2(n_43), .Y(n_327) );
OAI211xp5_ASAP7_75t_L g328 ( .A1(n_288), .A2(n_39), .B(n_44), .C(n_48), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_291), .A2(n_49), .B(n_50), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_301), .B(n_52), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_301), .B(n_53), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_287), .B(n_57), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_286), .B(n_58), .Y(n_339) );
INVx4_ASAP7_75t_R g340 ( .A(n_297), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_322), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_318), .B(n_296), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_322), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_336), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_318), .B(n_296), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_310), .B(n_290), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_303), .B(n_294), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_312), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_310), .B(n_290), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_326), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_310), .B(n_286), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_304), .B(n_294), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_313), .B(n_290), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_313), .B(n_290), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_304), .B(n_294), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_317), .B(n_282), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_305), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_304), .B(n_294), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_305), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_290), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_305), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_313), .B(n_287), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_339), .B(n_287), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_320), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_327), .A2(n_284), .B1(n_280), .B2(n_287), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_313), .B(n_281), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_339), .B(n_311), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_313), .B(n_299), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_313), .B(n_299), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_334), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_323), .Y(n_383) );
NAND2x1_ASAP7_75t_L g384 ( .A(n_316), .B(n_280), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_307), .B(n_291), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_339), .B(n_279), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_307), .B(n_59), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
INVx5_ASAP7_75t_L g389 ( .A(n_326), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_323), .Y(n_390) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_328), .B(n_279), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_307), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_317), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_309), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_307), .B(n_86), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_308), .B(n_311), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_308), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_308), .B(n_61), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_308), .Y(n_400) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_308), .B(n_62), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_311), .B(n_63), .Y(n_402) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_328), .B(n_64), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_325), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_311), .B(n_65), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_311), .B(n_69), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_354), .B(n_338), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_394), .B(n_329), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_345), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_354), .B(n_338), .Y(n_410) );
OR2x6_ASAP7_75t_SL g411 ( .A(n_377), .B(n_340), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_348), .B(n_325), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_390), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_363), .B(n_338), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_350), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_348), .B(n_325), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_350), .Y(n_418) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_381), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_352), .B(n_325), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_394), .B(n_329), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_351), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_352), .B(n_335), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_351), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g426 ( .A(n_374), .B(n_327), .C(n_332), .D(n_326), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_343), .B(n_335), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_370), .B(n_337), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_357), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_370), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_357), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_343), .B(n_335), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_370), .B(n_337), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_347), .B(n_335), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_366), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_347), .B(n_329), .Y(n_438) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_353), .B(n_332), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_380), .B(n_329), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_370), .B(n_337), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_366), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_380), .B(n_337), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_341), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_381), .B(n_333), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_353), .B(n_333), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_341), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_344), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_344), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_349), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_356), .B(n_333), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_360), .Y(n_454) );
NAND2xp33_ASAP7_75t_L g455 ( .A(n_389), .B(n_332), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_346), .B(n_333), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_369), .B(n_365), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_367), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_382), .B(n_338), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_367), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_372), .Y(n_461) );
AND2x2_ASAP7_75t_SL g462 ( .A(n_401), .B(n_331), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_387), .Y(n_463) );
NOR2xp33_ASAP7_75t_SL g464 ( .A(n_393), .B(n_340), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_369), .B(n_331), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_371), .B(n_338), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_355), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_358), .B(n_331), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_358), .B(n_309), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_359), .B(n_309), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_372), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_359), .B(n_316), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_365), .B(n_316), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_378), .B(n_316), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_355), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_378), .B(n_316), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_376), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_355), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_397), .B(n_336), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_376), .B(n_306), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_379), .B(n_316), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_401), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_362), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_362), .B(n_306), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_379), .B(n_321), .Y(n_485) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_389), .B(n_73), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_397), .B(n_321), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_404), .B(n_319), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_404), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_404), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_364), .B(n_321), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_364), .B(n_321), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_364), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_451), .B(n_386), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_409), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_457), .B(n_342), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_457), .B(n_342), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_452), .B(n_373), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_443), .B(n_404), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_415), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_445), .B(n_373), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_412), .B(n_342), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_412), .B(n_392), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_417), .B(n_392), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_434), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_417), .B(n_392), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_420), .B(n_398), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_420), .B(n_398), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_469), .B(n_398), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_469), .B(n_400), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_470), .B(n_400), .Y(n_512) );
NOR2x1p5_ASAP7_75t_SL g513 ( .A(n_491), .B(n_375), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_470), .B(n_389), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_454), .B(n_368), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_482), .B(n_389), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_407), .B(n_368), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_448), .B(n_385), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_449), .B(n_385), .Y(n_519) );
AND2x4_ASAP7_75t_SL g520 ( .A(n_482), .B(n_431), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_424), .B(n_389), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_418), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_423), .B(n_383), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_424), .B(n_389), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_475), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_413), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_465), .B(n_375), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_425), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_426), .A2(n_361), .B1(n_401), .B2(n_406), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_430), .B(n_383), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_432), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_462), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_437), .B(n_388), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_462), .A2(n_321), .B1(n_403), .B2(n_406), .Y(n_535) );
NAND2x1_ASAP7_75t_L g536 ( .A(n_431), .B(n_403), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_410), .B(n_388), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_442), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_414), .B(n_405), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_458), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_460), .B(n_384), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_486), .B(n_405), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_465), .B(n_319), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_489), .B(n_319), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_464), .B(n_391), .C(n_384), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_468), .B(n_319), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_478), .Y(n_548) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_431), .B(n_324), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_461), .B(n_315), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_490), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_468), .B(n_319), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_453), .B(n_402), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_453), .B(n_399), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_428), .B(n_324), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_419), .B(n_466), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_471), .B(n_315), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_477), .B(n_315), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_479), .B(n_395), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_483), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_440), .B(n_315), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_440), .B(n_444), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_428), .B(n_315), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_444), .B(n_391), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_433), .B(n_324), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_480), .B(n_324), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_489), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_433), .B(n_324), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_436), .B(n_324), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_408), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_408), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_436), .B(n_330), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_438), .B(n_330), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_480), .B(n_330), .Y(n_575) );
AOI32xp33_ASAP7_75t_L g576 ( .A1(n_455), .A2(n_75), .A3(n_76), .B1(n_78), .B2(n_79), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_421), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_421), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_416), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_416), .Y(n_580) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_422), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_422), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_427), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_439), .B(n_81), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_496), .B(n_439), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_543), .B(n_472), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_500), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_571), .B(n_438), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_572), .B(n_485), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_523), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_563), .B(n_456), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_577), .B(n_485), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_529), .Y(n_594) );
AOI21xp33_ASAP7_75t_L g595 ( .A1(n_546), .A2(n_490), .B(n_488), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_532), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_538), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_497), .B(n_490), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_578), .B(n_487), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_530), .B(n_411), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_527), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_520), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_510), .B(n_447), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_540), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_533), .A2(n_411), .B1(n_463), .B2(n_459), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_584), .A2(n_472), .B1(n_473), .B2(n_476), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_557), .B(n_456), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_527), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_507), .B(n_447), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_580), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_537), .B(n_484), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_498), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_517), .B(n_484), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_473), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_547), .B(n_474), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_516), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_553), .B(n_474), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_494), .B(n_487), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_568), .B(n_429), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_499), .Y(n_623) );
NOR2x1_ASAP7_75t_SL g624 ( .A(n_584), .B(n_446), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_508), .B(n_481), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_502), .B(n_481), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_494), .B(n_446), .Y(n_627) );
OAI22xp33_ASAP7_75t_SL g628 ( .A1(n_536), .A2(n_488), .B1(n_492), .B2(n_435), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_518), .B(n_450), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_524), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_561), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_524), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_503), .B(n_476), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_531), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_531), .Y(n_635) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_542), .B(n_455), .Y(n_636) );
NAND2x1_ASAP7_75t_SL g637 ( .A(n_516), .B(n_488), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_499), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_534), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_580), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_504), .B(n_435), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_518), .B(n_450), .Y(n_643) );
NOR2x1p5_ASAP7_75t_L g644 ( .A(n_549), .B(n_493), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_501), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_561), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_600), .A2(n_511), .B1(n_512), .B2(n_506), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_602), .A2(n_535), .A3(n_551), .B1(n_570), .B2(n_569), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_630), .Y(n_649) );
AOI221xp5_ASAP7_75t_SL g650 ( .A1(n_606), .A2(n_535), .B1(n_514), .B2(n_519), .C(n_525), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_624), .A2(n_576), .B(n_581), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_632), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_608), .B(n_519), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_600), .A2(n_513), .B(n_551), .C(n_522), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_635), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_636), .A2(n_544), .B(n_581), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_605), .A2(n_544), .B1(n_556), .B2(n_566), .Y(n_658) );
OAI321xp33_ASAP7_75t_L g659 ( .A1(n_606), .A2(n_560), .A3(n_541), .B1(n_564), .B2(n_554), .C(n_555), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_607), .A2(n_573), .B1(n_574), .B2(n_539), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_623), .B(n_505), .Y(n_661) );
AOI211xp5_ASAP7_75t_SL g662 ( .A1(n_605), .A2(n_567), .B(n_541), .C(n_575), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_639), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_609), .B(n_641), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_615), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_628), .A2(n_575), .B(n_550), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_616), .B(n_515), .Y(n_667) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_621), .A2(n_562), .A3(n_567), .B1(n_501), .B2(n_559), .C1(n_558), .C2(n_550), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_631), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_607), .A2(n_562), .B(n_558), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_645), .B(n_582), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_585), .A2(n_579), .B1(n_559), .B2(n_583), .C1(n_552), .C2(n_548), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_605), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_588), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_619), .B(n_509), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_631), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_587), .B(n_583), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_638), .B(n_545), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_638), .B(n_526), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_591), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_594), .A2(n_521), .B1(n_435), .B2(n_441), .C(n_429), .Y(n_681) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_595), .A2(n_619), .B(n_586), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_665), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_659), .A2(n_604), .B1(n_597), .B2(n_596), .C(n_627), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_659), .A2(n_646), .B1(n_599), .B2(n_593), .C(n_590), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_666), .A2(n_644), .B1(n_622), .B2(n_646), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_651), .A2(n_622), .B(n_637), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_654), .A2(n_642), .B(n_625), .C(n_598), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_672), .B(n_587), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_650), .A2(n_643), .B1(n_629), .B2(n_589), .C(n_618), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g691 ( .A1(n_682), .A2(n_614), .B(n_610), .Y(n_691) );
NOR4xp25_ASAP7_75t_SL g692 ( .A(n_675), .B(n_592), .C(n_617), .D(n_633), .Y(n_692) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_660), .A2(n_620), .B(n_618), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g694 ( .A1(n_648), .A2(n_620), .B1(n_617), .B2(n_626), .C1(n_612), .C2(n_603), .Y(n_694) );
NOR2xp33_ASAP7_75t_SL g695 ( .A(n_676), .B(n_661), .Y(n_695) );
OAI22xp5_ASAP7_75t_SL g696 ( .A1(n_647), .A2(n_640), .B1(n_613), .B2(n_611), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_658), .A2(n_441), .B1(n_611), .B2(n_601), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_672), .B(n_670), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_662), .A2(n_657), .B(n_681), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_668), .A2(n_653), .B(n_671), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_669), .B(n_679), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_678), .A2(n_649), .B1(n_652), .B2(n_655), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_656), .B(n_663), .C(n_674), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_680), .B(n_664), .C(n_677), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_667), .B(n_672), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_647), .B(n_673), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_654), .A2(n_659), .B(n_651), .Y(n_707) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_687), .B(n_707), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_683), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_698), .B(n_706), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_705), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_700), .B(n_689), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_708), .B(n_694), .C(n_685), .D(n_684), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_712), .A2(n_699), .B1(n_686), .B2(n_693), .C(n_691), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_710), .B(n_690), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_714), .B(n_692), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_713), .B(n_711), .C(n_686), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_717), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_716), .Y(n_719) );
XNOR2xp5_ASAP7_75t_L g720 ( .A(n_719), .B(n_715), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_718), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_720), .A2(n_709), .B(n_695), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_722), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_721), .B(n_688), .Y(n_724) );
OA21x2_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_704), .B(n_703), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_697), .B1(n_696), .B2(n_702), .C(n_701), .Y(n_726) );
endmodule