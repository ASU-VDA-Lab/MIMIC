module real_jpeg_4963_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_487;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_0),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_0),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_0),
.Y(n_309)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_0),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_1),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_1),
.A2(n_151),
.B1(n_199),
.B2(n_268),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_1),
.A2(n_82),
.B1(n_268),
.B2(n_389),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g445 ( 
.A1(n_1),
.A2(n_268),
.B1(n_325),
.B2(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_2),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_2),
.Y(n_334)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_2),
.Y(n_349)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_2),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_2),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_55),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_3),
.A2(n_55),
.B1(n_127),
.B2(n_179),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_3),
.A2(n_55),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_4),
.Y(n_527)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_5),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_6),
.A2(n_68),
.B1(n_303),
.B2(n_306),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_6),
.A2(n_68),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_6),
.A2(n_68),
.B1(n_272),
.B2(n_391),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_7),
.A2(n_151),
.B1(n_153),
.B2(n_155),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_7),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_7),
.B(n_124),
.C(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_7),
.B(n_87),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_7),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_7),
.B(n_160),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_7),
.B(n_105),
.Y(n_256)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_8),
.Y(n_524)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_11),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_11),
.A2(n_49),
.B1(n_103),
.B2(n_107),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_49),
.B1(n_113),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_11),
.A2(n_49),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_12),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_200),
.B1(n_219),
.B2(n_222),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_12),
.A2(n_105),
.B1(n_200),
.B2(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_12),
.A2(n_65),
.B1(n_200),
.B2(n_353),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_13),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_13),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_113),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_14),
.A2(n_159),
.B1(n_189),
.B2(n_193),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_14),
.A2(n_159),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_14),
.A2(n_159),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_174),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_16),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_16),
.A2(n_178),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_16),
.A2(n_178),
.B1(n_294),
.B2(n_359),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_16),
.A2(n_67),
.B1(n_178),
.B2(n_397),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_17),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_17),
.A2(n_74),
.B1(n_166),
.B2(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_17),
.A2(n_74),
.B1(n_135),
.B2(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_17),
.A2(n_74),
.B1(n_273),
.B2(n_432),
.Y(n_431)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_522),
.B(n_525),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_58),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_50),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_24),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_24),
.B(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_25),
.B(n_155),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_25),
.A2(n_51),
.B1(n_396),
.B2(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_25)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_26),
.A2(n_319),
.A3(n_322),
.B1(n_326),
.B2(n_331),
.Y(n_318)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_38)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_30),
.Y(n_274)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_31),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_31),
.Y(n_262)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_34),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_37),
.A2(n_347),
.B(n_350),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_37),
.B(n_352),
.Y(n_448)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_43),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_50)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_50),
.B(n_60),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_69),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_69),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_51),
.A2(n_351),
.B(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_56),
.A2(n_420),
.B(n_448),
.Y(n_458)
);

AO21x1_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_140),
.B(n_521),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_136),
.C(n_137),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_61),
.A2(n_62),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_75),
.C(n_108),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_63),
.B(n_509),
.Y(n_508)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_75),
.A2(n_108),
.B1(n_109),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_75),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_95),
.B1(n_101),
.B2(n_102),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_76),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_76),
.A2(n_101),
.B1(n_293),
.B2(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_76),
.A2(n_101),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_76),
.A2(n_95),
.B1(n_101),
.B2(n_498),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_78),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_81),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_86),
.Y(n_254)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_86),
.Y(n_321)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_86),
.Y(n_330)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_86),
.Y(n_394)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_86),
.Y(n_433)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_87),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

AOI22x1_ASAP7_75t_L g421 ( 
.A1(n_87),
.A2(n_138),
.B1(n_298),
.B2(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_87),
.A2(n_138),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_94),
.Y(n_87)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_89),
.Y(n_276)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_90),
.Y(n_385)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_91),
.Y(n_381)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_101),
.B(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_101),
.A2(n_293),
.B(n_297),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_106),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_108),
.A2(n_109),
.B1(n_496),
.B2(n_497),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_108),
.B(n_493),
.C(n_496),
.Y(n_504)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_123),
.B(n_134),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_110),
.A2(n_150),
.B(n_156),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_110),
.A2(n_197),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_110),
.A2(n_156),
.B(n_247),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_110),
.A2(n_246),
.B1(n_363),
.B2(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_111),
.B(n_157),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_111),
.A2(n_160),
.B1(n_377),
.B2(n_382),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_111),
.A2(n_160),
.B1(n_382),
.B2(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_111),
.A2(n_160),
.B1(n_402),
.B2(n_436),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_123),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx5_ASAP7_75t_SL g250 ( 
.A(n_120),
.Y(n_250)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_123),
.A2(n_197),
.B(n_203),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_123),
.A2(n_203),
.B(n_363),
.Y(n_362)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_134),
.Y(n_436)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_135),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_136),
.B(n_137),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_138),
.A2(n_253),
.B(n_257),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_138),
.B(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_138),
.A2(n_257),
.B(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_515),
.B(n_520),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_487),
.B(n_512),
.Y(n_141)
);

OAI311xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_366),
.A3(n_463),
.B1(n_481),
.C1(n_486),
.Y(n_142)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_312),
.B(n_365),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_284),
.B(n_311),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_240),
.B(n_283),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_206),
.B(n_239),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_171),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_148),
.B(n_171),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_161),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_149),
.A2(n_161),
.B1(n_162),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_149),
.Y(n_237)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_153),
.B(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_153),
.Y(n_404)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g403 ( 
.A(n_154),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_155),
.A2(n_181),
.B(n_186),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g253 ( 
.A1(n_155),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_155),
.B(n_332),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_155),
.A2(n_331),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_194),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_195),
.C(n_205),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_181),
.B(n_186),
.Y(n_172)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_176),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_181),
.A2(n_212),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_181),
.A2(n_235),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_181),
.A2(n_373),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_188),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_182),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_182),
.A2(n_266),
.B1(n_302),
.B2(n_308),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_182),
.A2(n_339),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_184),
.Y(n_269)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_191),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_192),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_204),
.B2(n_205),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_230),
.B(n_238),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_216),
.B(n_229),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_225),
.B(n_227),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_219),
.Y(n_375)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_265),
.B(n_270),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_236),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_242),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_263),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_251),
.B2(n_252),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_251),
.C(n_263),
.Y(n_285)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI32xp33_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_272),
.A3(n_275),
.B1(n_277),
.B2(n_281),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_274),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_276),
.Y(n_378)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_285),
.B(n_286),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_310),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_290),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_292),
.B(n_300),
.C(n_301),
.Y(n_341)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_313),
.B(n_314),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_344),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_315)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_335),
.B2(n_336),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_318),
.B(n_335),
.Y(n_459)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_341),
.B(n_342),
.C(n_344),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_356),
.B2(n_364),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_345),
.B(n_357),
.C(n_362),
.Y(n_472)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_356),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_358),
.Y(n_461)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_449),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_367),
.A2(n_449),
.B(n_482),
.C(n_485),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_423),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_368),
.B(n_423),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_399),
.C(n_408),
.Y(n_368)
);

FAx1_ASAP7_75t_SL g462 ( 
.A(n_369),
.B(n_399),
.CI(n_408),
.CON(n_462),
.SN(n_462)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_386),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_370),
.B(n_387),
.C(n_395),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_371),
.B(n_376),
.Y(n_455)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_395),
.Y(n_386)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_405),
.B2(n_407),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_405),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_405),
.A2(n_407),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_405),
.A2(n_440),
.B(n_443),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_418),
.C(n_421),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_410),
.B(n_412),
.Y(n_471)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx8_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_418),
.A2(n_419),
.B1(n_421),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_421),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_424),
.B(n_427),
.C(n_438),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_438),
.B2(n_439),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_434),
.B(n_437),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_435),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_431),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_437),
.B(n_490),
.CI(n_491),
.CON(n_489),
.SN(n_489)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_490),
.C(n_491),
.Y(n_511)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_448),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_462),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_462),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_455),
.C(n_456),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_451),
.A2(n_452),
.B1(n_455),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_455),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.C(n_460),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_457),
.A2(n_458),
.B1(n_460),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_460),
.Y(n_469)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_462),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_476),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_465),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_473),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_473),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.C(n_472),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_479),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_471),
.B1(n_472),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_472),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_478),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_501),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_500),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_500),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_489),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_493),
.B1(n_495),
.B2(n_499),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_493),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_503),
.C(n_507),
.Y(n_519)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_495),
.Y(n_499)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_511),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_511),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_519),
.Y(n_520)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_523),
.Y(n_526)
);

INVx13_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.Y(n_525)
);


endmodule