module fake_jpeg_17445_n_174 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_53),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_50),
.B(n_62),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_81),
.Y(n_113)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_67),
.B1(n_62),
.B2(n_47),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_94),
.B1(n_51),
.B2(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_72),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_64),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_66),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_51),
.B1(n_65),
.B2(n_44),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_120),
.B1(n_59),
.B2(n_48),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_106),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_0),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_45),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_46),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_58),
.C(n_52),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_1),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_119),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_116),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_58),
.C(n_52),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_47),
.Y(n_125)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_131),
.B1(n_104),
.B2(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_97),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_138),
.Y(n_142)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_139),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_141),
.B1(n_96),
.B2(n_106),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_126),
.B1(n_132),
.B2(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_95),
.C(n_128),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_146),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_121),
.B1(n_108),
.B2(n_130),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_134),
.B(n_137),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_133),
.B(n_127),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_143),
.B(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_135),
.C(n_105),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_130),
.Y(n_158)
);

AOI211xp5_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_158),
.B(n_102),
.C(n_3),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_151),
.B1(n_127),
.B2(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_24),
.B1(n_43),
.B2(n_41),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_23),
.B(n_40),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_22),
.C(n_39),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_20),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_15),
.B(n_38),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_14),
.B(n_37),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_13),
.B(n_36),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_11),
.B(n_33),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_172),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_9),
.Y(n_174)
);


endmodule