module fake_jpeg_7732_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_12),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_58),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_12),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_19),
.B1(n_17),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_62),
.B1(n_29),
.B2(n_25),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_32),
.B1(n_35),
.B2(n_19),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_74),
.B1(n_21),
.B2(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_66),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_19),
.B1(n_34),
.B2(n_35),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_21),
.B1(n_35),
.B2(n_32),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_69),
.B1(n_23),
.B2(n_16),
.Y(n_114)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_71),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_47),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_21),
.B1(n_32),
.B2(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_16),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_34),
.B1(n_26),
.B2(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_80),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_46),
.C(n_39),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_4),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_15),
.B(n_14),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_53),
.A3(n_68),
.B1(n_13),
.B2(n_15),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_27),
.B(n_20),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_92),
.B(n_106),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_101),
.B1(n_112),
.B2(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_31),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_28),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NAND2x1p5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_109),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_61),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_24),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_39),
.B(n_33),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_65),
.B(n_56),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_14),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_33),
.B1(n_47),
.B2(n_45),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_5),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_66),
.B1(n_49),
.B2(n_47),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_124),
.A2(n_136),
.B1(n_140),
.B2(n_108),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_104),
.B1(n_107),
.B2(n_110),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_49),
.B1(n_45),
.B2(n_39),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_96),
.B1(n_80),
.B2(n_99),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_106),
.B(n_95),
.Y(n_150)
);

OAI211xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_45),
.B(n_33),
.C(n_65),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_115),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_87),
.B1(n_83),
.B2(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_144),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_56),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_82),
.B1(n_84),
.B2(n_93),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_5),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_151),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_148),
.A2(n_154),
.B1(n_157),
.B2(n_160),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_113),
.C(n_98),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_179),
.C(n_133),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_177),
.B(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_118),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_132),
.B1(n_134),
.B2(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_153),
.B(n_158),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_146),
.A2(n_95),
.B1(n_99),
.B2(n_85),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_156),
.Y(n_192)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_129),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_165),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_108),
.B1(n_105),
.B2(n_81),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_167),
.B1(n_178),
.B2(n_139),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_5),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_6),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_6),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_7),
.Y(n_174)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_123),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_141),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_90),
.C(n_78),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_182),
.A2(n_188),
.B1(n_205),
.B2(n_206),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_177),
.C(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_155),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_156),
.B1(n_168),
.B2(n_171),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_125),
.B1(n_135),
.B2(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_196),
.B(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_128),
.B(n_129),
.Y(n_196)
);

AO22x1_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_129),
.B1(n_123),
.B2(n_131),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_139),
.B1(n_131),
.B2(n_121),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_137),
.B1(n_142),
.B2(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_142),
.B1(n_127),
.B2(n_117),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_161),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_122),
.B1(n_77),
.B2(n_9),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_122),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_149),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_219),
.Y(n_241)
);

AOI22x1_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_150),
.B1(n_162),
.B2(n_153),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_240),
.B1(n_199),
.B2(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_218),
.B(n_220),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_222),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_172),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_234),
.B1(n_203),
.B2(n_205),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_238),
.B1(n_191),
.B2(n_181),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_158),
.C(n_8),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_7),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_7),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_7),
.C(n_8),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_216),
.B1(n_225),
.B2(n_223),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_199),
.B(n_196),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_246),
.B(n_216),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_188),
.B1(n_206),
.B2(n_182),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_249),
.B1(n_229),
.B2(n_230),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_260),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_203),
.B1(n_204),
.B2(n_197),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_258),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_180),
.B1(n_212),
.B2(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_212),
.B1(n_194),
.B2(n_193),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_208),
.B1(n_185),
.B2(n_186),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_186),
.B1(n_10),
.B2(n_11),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_239),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_213),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_272),
.Y(n_292)
);

AOI221xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_243),
.B1(n_254),
.B2(n_256),
.C(n_259),
.Y(n_288)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_241),
.C(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_277),
.C(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_221),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_273),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_219),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_242),
.B(n_261),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_217),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_278),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_222),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_229),
.B(n_234),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_235),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_251),
.B(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_217),
.C(n_240),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_11),
.C(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

AOI21x1_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_245),
.B(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_291),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_267),
.A2(n_246),
.B(n_242),
.C(n_261),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_273),
.B(n_10),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_265),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_257),
.B1(n_251),
.B2(n_11),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_9),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_270),
.C(n_264),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.C(n_304),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_277),
.C(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_281),
.C(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_266),
.C(n_282),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_284),
.B(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_296),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_11),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_290),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_293),
.B1(n_294),
.B2(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_312),
.B(n_314),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_306),
.B(n_303),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_295),
.B1(n_290),
.B2(n_289),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_316),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_303),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_317),
.C(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_307),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_313),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_312),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_329),
.B(n_325),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_314),
.B1(n_315),
.B2(n_304),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_327),
.Y(n_331)
);

AOI31xp33_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_325),
.A3(n_328),
.B(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_331),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_302),
.Y(n_336)
);


endmodule