module fake_jpeg_14941_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_3),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_3),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

AND2x2_ASAP7_75t_SL g11 ( 
.A(n_4),
.B(n_5),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

HAxp5_ASAP7_75t_SL g13 ( 
.A(n_4),
.B(n_3),
.CON(n_13),
.SN(n_13)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_18),
.B1(n_19),
.B2(n_7),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_11),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_1),
.B1(n_2),
.B2(n_8),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_12),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_7),
.C(n_12),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_26),
.B(n_24),
.Y(n_34)
);

BUFx24_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_10),
.B1(n_12),
.B2(n_21),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_12),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_24),
.C(n_28),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_22),
.C(n_26),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_37),
.C(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_32),
.Y(n_38)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_33),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_30),
.C(n_24),
.Y(n_41)
);


endmodule