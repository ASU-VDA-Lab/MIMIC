module fake_ibex_1515_n_4306 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4306);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4306;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_962;
wire n_1080;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3819;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4179;
wire n_3340;
wire n_4142;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3653;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_3904;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_2918;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3856;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3949;
wire n_3507;
wire n_3881;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3766;
wire n_2822;
wire n_3148;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3910;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3769;
wire n_2813;
wire n_2147;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_3217;
wire n_2511;
wire n_2782;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3887;
wire n_3800;
wire n_3963;
wire n_3317;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3983;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_4062;
wire n_2375;
wire n_2964;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_3331;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_4114;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_3558;
wire n_2751;
wire n_2785;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_4097;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_4215;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3797;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3584;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3646;
wire n_3477;
wire n_2635;
wire n_3070;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_3557;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_3495;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_3498;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_4278;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_4227;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_3902;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_4133;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1349;
wire n_1223;
wire n_1331;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_4138;
wire n_3499;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3828;
wire n_3240;
wire n_3336;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3673;
wire n_3476;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3746;
wire n_2758;
wire n_3480;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_4068;
wire n_1063;
wire n_3021;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_3512;
wire n_2963;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_4282;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3454;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3604;
wire n_1838;
wire n_3649;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_4032;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_3236;
wire n_2658;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_4265;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3013;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_1586;
wire n_1547;
wire n_1362;
wire n_946;
wire n_3497;
wire n_4178;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_3899;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_4281;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_4045;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3655;
wire n_3543;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_2371;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_1193;
wire n_3225;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3067;
wire n_1074;
wire n_3380;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3823;
wire n_3369;
wire n_3606;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_999;
wire n_2634;
wire n_2982;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_1762;
wire n_940;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3933;
wire n_2262;
wire n_3516;
wire n_3562;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_3193;
wire n_3635;
wire n_3501;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2349;
wire n_2100;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2673;
wire n_2430;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3494;
wire n_3040;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_300),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_480),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_914),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_757),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_710),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_357),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_79),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_400),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_106),
.Y(n_939)
);

BUFx10_ASAP7_75t_L g940 ( 
.A(n_771),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_164),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_847),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_305),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_488),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_263),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_618),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_688),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_659),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_135),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_477),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_908),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_267),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_113),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_724),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_64),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_385),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_544),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_108),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_884),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_278),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_454),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_503),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_906),
.Y(n_963)
);

CKINVDCx16_ASAP7_75t_R g964 ( 
.A(n_861),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_94),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_429),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_637),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_177),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_481),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_524),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_907),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_72),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_282),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_806),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_505),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_926),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_538),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_466),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_716),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_272),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_429),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_895),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_625),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_192),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_580),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_276),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_53),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_284),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_568),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_477),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_435),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_610),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_302),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_599),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_508),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_913),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_125),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_341),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_679),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_897),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_333),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_813),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_418),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_344),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_110),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_683),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_283),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_414),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_672),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_666),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_527),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_310),
.Y(n_1012)
);

BUFx10_ASAP7_75t_L g1013 ( 
.A(n_564),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_891),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_618),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_218),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_911),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_292),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_896),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_794),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_777),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_260),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_219),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_708),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_882),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_594),
.Y(n_1026)
);

BUFx5_ASAP7_75t_L g1027 ( 
.A(n_506),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_898),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_249),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_539),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_746),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_900),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_499),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_63),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_787),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_543),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_628),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_123),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_820),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_488),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_1),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_710),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_310),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_6),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_393),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_159),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_919),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_338),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_220),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_720),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_734),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_415),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_447),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_136),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_510),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_0),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_315),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_333),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_380),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_860),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_245),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_356),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_720),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_548),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_280),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_217),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_136),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_397),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_901),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_568),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_377),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_651),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_496),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_356),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_562),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_585),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_283),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_678),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_382),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_66),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_26),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_365),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_864),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_388),
.Y(n_1084)
);

CKINVDCx16_ASAP7_75t_R g1085 ( 
.A(n_905),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_161),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_466),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_656),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_890),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_337),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_889),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_404),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_416),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_732),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_727),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_829),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_650),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_783),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_711),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_903),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_473),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_405),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_211),
.Y(n_1103)
);

CKINVDCx16_ASAP7_75t_R g1104 ( 
.A(n_139),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_598),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_152),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_577),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_581),
.Y(n_1108)
);

CKINVDCx14_ASAP7_75t_R g1109 ( 
.A(n_495),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_639),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_926),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_28),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_662),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_888),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_886),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_714),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_763),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_483),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_764),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_541),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_285),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_621),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_684),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_860),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_513),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_697),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_645),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_902),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_604),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_704),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_754),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_481),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_139),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_435),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_885),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_7),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_19),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_783),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_326),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_77),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_394),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_641),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_899),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_81),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_894),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_450),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_53),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_830),
.Y(n_1149)
);

BUFx10_ASAP7_75t_L g1150 ( 
.A(n_358),
.Y(n_1150)
);

CKINVDCx16_ASAP7_75t_R g1151 ( 
.A(n_353),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_611),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_910),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_304),
.Y(n_1154)
);

BUFx5_ASAP7_75t_L g1155 ( 
.A(n_656),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_474),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_881),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_317),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_605),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_221),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_793),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_868),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_799),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_666),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_116),
.Y(n_1165)
);

BUFx5_ASAP7_75t_L g1166 ( 
.A(n_930),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_887),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_504),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_146),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_626),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_624),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_476),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_361),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_227),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_485),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_176),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_257),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_64),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_230),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_265),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_296),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_433),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_836),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_771),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_348),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_474),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_655),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_247),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_327),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_593),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_592),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_630),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_156),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_352),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_893),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_121),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_707),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_690),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_362),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_468),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_800),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_582),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_496),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_653),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_545),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_914),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_245),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_63),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_175),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_816),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_713),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_365),
.Y(n_1212)
);

BUFx5_ASAP7_75t_L g1213 ( 
.A(n_402),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_321),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_147),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_148),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_430),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_214),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_809),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_383),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_565),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_879),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_904),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_415),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_331),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_222),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_405),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_586),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_699),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_231),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_387),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_68),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_735),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_909),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_845),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_608),
.Y(n_1236)
);

BUFx5_ASAP7_75t_L g1237 ( 
.A(n_158),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_563),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_622),
.Y(n_1239)
);

BUFx5_ASAP7_75t_L g1240 ( 
.A(n_901),
.Y(n_1240)
);

INVxp33_ASAP7_75t_L g1241 ( 
.A(n_287),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_810),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_115),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_909),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_325),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_545),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_251),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_681),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_402),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_240),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_705),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_69),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_154),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_638),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_588),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_925),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_15),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_906),
.Y(n_1258)
);

CKINVDCx16_ASAP7_75t_R g1259 ( 
.A(n_885),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_847),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_522),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_198),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_142),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_510),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_551),
.Y(n_1265)
);

BUFx8_ASAP7_75t_SL g1266 ( 
.A(n_87),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_552),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_658),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_679),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_119),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_912),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_883),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_646),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_127),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_892),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_414),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_584),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_691),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_162),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_786),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_649),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_900),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_64),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_217),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_866),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_917),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_147),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_404),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_162),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_121),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_800),
.Y(n_1291)
);

CKINVDCx16_ASAP7_75t_R g1292 ( 
.A(n_864),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_54),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_653),
.Y(n_1294)
);

BUFx8_ASAP7_75t_SL g1295 ( 
.A(n_620),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_552),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_144),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_98),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_99),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_472),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_364),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_69),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_5),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_725),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_675),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_796),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_927),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_753),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_53),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_636),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_141),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_851),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_867),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_638),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_463),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_269),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_701),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_293),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_184),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_573),
.Y(n_1320)
);

CKINVDCx16_ASAP7_75t_R g1321 ( 
.A(n_804),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_463),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_184),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_482),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_779),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_309),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_752),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_267),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_527),
.Y(n_1329)
);

INVx4_ASAP7_75t_R g1330 ( 
.A(n_747),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_663),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_222),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_630),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_188),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_814),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_62),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_471),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_365),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_333),
.Y(n_1339)
);

CKINVDCx14_ASAP7_75t_R g1340 ( 
.A(n_464),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_6),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_645),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_205),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_849),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_657),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_105),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_620),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_483),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_308),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_105),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_233),
.Y(n_1351)
);

CKINVDCx16_ASAP7_75t_R g1352 ( 
.A(n_381),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_489),
.Y(n_1353)
);

BUFx10_ASAP7_75t_L g1354 ( 
.A(n_752),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_921),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_433),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_776),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_868),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_214),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_716),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1340),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1340),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1266),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1241),
.Y(n_1364)
);

CKINVDCx16_ASAP7_75t_R g1365 ( 
.A(n_1104),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1194),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1125),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_1008),
.B(n_0),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1346),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1052),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1103),
.B(n_0),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1245),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1109),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_941),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1295),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_949),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_941),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1241),
.B(n_1),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_952),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1178),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1295),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1178),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1151),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1352),
.B(n_2),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1029),
.B(n_2),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_984),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1169),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_955),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_947),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1169),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_984),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_931),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1213),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_958),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1120),
.B(n_2),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_960),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_R g1397 ( 
.A(n_1020),
.B(n_3),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_961),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_987),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1207),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_965),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1201),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1218),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_987),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_988),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_997),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1005),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_936),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_937),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1263),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_938),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_939),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1007),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1016),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_943),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_R g1416 ( 
.A(n_945),
.B(n_4),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_953),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1263),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_956),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1049),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1065),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_966),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1068),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1071),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1244),
.B(n_5),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_972),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1300),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_968),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1001),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1034),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_973),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1029),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1056),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1081),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1084),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1270),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1213),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_980),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_986),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1086),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1090),
.Y(n_1441)
);

INVxp67_ASAP7_75t_SL g1442 ( 
.A(n_1177),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1092),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1364),
.B(n_991),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1386),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1393),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1437),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1437),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1368),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1391),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1399),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1404),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1442),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1372),
.B(n_1029),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1366),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1392),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1369),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1389),
.B(n_1239),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1376),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1371),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1379),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1388),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1367),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1394),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1396),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1398),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1401),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1432),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1370),
.B(n_1335),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1361),
.B(n_1213),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1405),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1362),
.B(n_993),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1406),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1407),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1413),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1414),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1420),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1421),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1423),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1424),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1435),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1436),
.B(n_998),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1402),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1441),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1385),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1427),
.B(n_1150),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1371),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1408),
.Y(n_1488)
);

AND2x6_ASAP7_75t_L g1489 ( 
.A(n_1378),
.B(n_1177),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1395),
.Y(n_1490)
);

CKINVDCx8_ASAP7_75t_R g1491 ( 
.A(n_1363),
.Y(n_1491)
);

XOR2xp5_ASAP7_75t_L g1492 ( 
.A(n_1419),
.B(n_1121),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1374),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1365),
.B(n_1150),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1425),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1384),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1409),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1373),
.B(n_1004),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1411),
.Y(n_1499)
);

NAND2x1_ASAP7_75t_L g1500 ( 
.A(n_1397),
.B(n_1330),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1412),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1415),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1417),
.B(n_1012),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1416),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1422),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1416),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1428),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1431),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1438),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1439),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1377),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1383),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1375),
.B(n_1150),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1381),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1380),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1426),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1382),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1387),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1390),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1429),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1400),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1403),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1410),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1418),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1430),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1433),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1434),
.B(n_964),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1440),
.B(n_1213),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1443),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1364),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1367),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1386),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1386),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1366),
.B(n_1085),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1364),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1386),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1364),
.B(n_1018),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1364),
.B(n_1022),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1386),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1364),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1364),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1386),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1367),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1386),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1367),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1364),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1386),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1386),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1364),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1367),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1367),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1367),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1364),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1364),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1363),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1392),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1364),
.B(n_942),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1367),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1367),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1364),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1386),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1386),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1367),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1364),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1364),
.B(n_1023),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1364),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1392),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1364),
.B(n_1179),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1364),
.B(n_942),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1364),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1364),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1364),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1364),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1432),
.B(n_1237),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1393),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1386),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1393),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1393),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1386),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1393),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1386),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1367),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1386),
.Y(n_1583)
);

INVx6_ASAP7_75t_L g1584 ( 
.A(n_1371),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1367),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1364),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1455),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1487),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1468),
.B(n_1138),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1531),
.B(n_1259),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1457),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1545),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1460),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1495),
.B(n_1179),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1460),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1502),
.B(n_1140),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1485),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1450),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1568),
.B(n_1237),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1456),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1463),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1550),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1584),
.Y(n_1603)
);

INVx5_ASAP7_75t_L g1604 ( 
.A(n_1536),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1450),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1536),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1451),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1444),
.B(n_1537),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1543),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1556),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1451),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1567),
.B(n_1153),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1584),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1558),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1538),
.B(n_1237),
.Y(n_1615)
);

BUFx8_ASAP7_75t_SL g1616 ( 
.A(n_1493),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1548),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1516),
.B(n_1153),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1504),
.B(n_1196),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1551),
.B(n_1292),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1496),
.A2(n_1145),
.B1(n_1158),
.B2(n_1141),
.Y(n_1621)
);

AND2x6_ASAP7_75t_L g1622 ( 
.A(n_1506),
.B(n_1003),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1552),
.B(n_1321),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1582),
.Y(n_1625)
);

BUFx10_ASAP7_75t_L g1626 ( 
.A(n_1555),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1452),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1565),
.B(n_1237),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1454),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1559),
.B(n_1196),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1452),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1486),
.Y(n_1632)
);

OA22x2_ASAP7_75t_L g1633 ( 
.A1(n_1563),
.A2(n_1043),
.B1(n_1044),
.B2(n_1041),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1535),
.B(n_1045),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1542),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1469),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1542),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1453),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1453),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1532),
.Y(n_1640)
);

INVx6_ASAP7_75t_L g1641 ( 
.A(n_1514),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1464),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1511),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1492),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1464),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1585),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1483),
.B(n_940),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1464),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1482),
.B(n_940),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1488),
.B(n_1197),
.Y(n_1650)
);

INVx5_ASAP7_75t_L g1651 ( 
.A(n_1480),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1540),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1533),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1541),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1534),
.B(n_1048),
.C(n_1046),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1489),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1546),
.B(n_1053),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1549),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1553),
.B(n_1057),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1576),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1554),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1579),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1579),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1560),
.B(n_1058),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1503),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1564),
.A2(n_1359),
.B1(n_1059),
.B2(n_1062),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1566),
.A2(n_1066),
.B1(n_1067),
.B2(n_1061),
.Y(n_1667)
);

AND2x6_ASAP7_75t_L g1668 ( 
.A(n_1570),
.B(n_1038),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1571),
.B(n_1074),
.Y(n_1669)
);

NAND3x1_ASAP7_75t_L g1670 ( 
.A(n_1525),
.B(n_1222),
.C(n_1197),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1469),
.Y(n_1671)
);

BUFx10_ASAP7_75t_L g1672 ( 
.A(n_1458),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1586),
.B(n_1349),
.Y(n_1674)
);

NOR2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1500),
.B(n_1080),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1557),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1569),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1497),
.B(n_1028),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1462),
.B(n_1093),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_L g1680 ( 
.A(n_1489),
.B(n_1027),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1449),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1513),
.Y(n_1682)
);

INVx5_ASAP7_75t_L g1683 ( 
.A(n_1489),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1459),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1461),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1465),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1473),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1498),
.B(n_1038),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1499),
.B(n_1028),
.Y(n_1689)
);

CKINVDCx9p33_ASAP7_75t_R g1690 ( 
.A(n_1527),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1477),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1479),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1466),
.B(n_1102),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1484),
.Y(n_1694)
);

AND2x6_ASAP7_75t_L g1695 ( 
.A(n_1507),
.B(n_1082),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1491),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1467),
.B(n_1351),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1471),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1501),
.B(n_1106),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1474),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1475),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1476),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1478),
.B(n_1481),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1539),
.Y(n_1704)
);

INVx5_ASAP7_75t_L g1705 ( 
.A(n_1544),
.Y(n_1705)
);

INVx4_ASAP7_75t_SL g1706 ( 
.A(n_1508),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_1547),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1490),
.B(n_1112),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1505),
.B(n_1509),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1510),
.A2(n_1173),
.B1(n_1182),
.B2(n_1180),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1446),
.A2(n_1188),
.B1(n_1199),
.B2(n_1193),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1561),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1562),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1512),
.B(n_1170),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1528),
.B(n_1170),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1574),
.B(n_1135),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1520),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1470),
.B(n_1205),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1581),
.B(n_1137),
.Y(n_1719)
);

AND2x6_ASAP7_75t_L g1720 ( 
.A(n_1447),
.B(n_1082),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1529),
.B(n_940),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1448),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1575),
.B(n_1142),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1515),
.B(n_990),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1577),
.B(n_1147),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1578),
.B(n_1148),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1526),
.B(n_1205),
.Y(n_1727)
);

AND2x6_ASAP7_75t_L g1728 ( 
.A(n_1578),
.B(n_1257),
.Y(n_1728)
);

AND2x6_ASAP7_75t_L g1729 ( 
.A(n_1580),
.B(n_1257),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1519),
.B(n_1337),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1580),
.A2(n_1212),
.B1(n_1215),
.B2(n_1208),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1472),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1524),
.B(n_1154),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1517),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1517),
.A2(n_1231),
.B1(n_1232),
.B2(n_1217),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1518),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1521),
.B(n_1303),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1522),
.B(n_1337),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1523),
.Y(n_1739)
);

INVx4_ASAP7_75t_L g1740 ( 
.A(n_1468),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1468),
.B(n_1222),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1530),
.B(n_1160),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1530),
.B(n_1165),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1445),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1493),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1455),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1468),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1468),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1445),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1531),
.B(n_990),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1531),
.B(n_1079),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1468),
.Y(n_1752)
);

BUFx4_ASAP7_75t_L g1753 ( 
.A(n_1525),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1468),
.B(n_1234),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1468),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1455),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1531),
.B(n_1013),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1493),
.A2(n_1236),
.B1(n_1256),
.B2(n_1234),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1468),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1445),
.Y(n_1760)
);

AND2x4_ASAP7_75t_SL g1761 ( 
.A(n_1494),
.B(n_1013),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1468),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1495),
.B(n_1174),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1530),
.B(n_1176),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1495),
.B(n_1181),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1530),
.B(n_1185),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1487),
.B(n_1336),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1468),
.B(n_948),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1748),
.B(n_1236),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1598),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1755),
.B(n_1134),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1592),
.B(n_1256),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1614),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1608),
.B(n_1189),
.Y(n_1774)
);

AO22x2_ASAP7_75t_L g1775 ( 
.A1(n_1741),
.A2(n_1319),
.B1(n_1220),
.B2(n_1294),
.Y(n_1775)
);

BUFx8_ASAP7_75t_L g1776 ( 
.A(n_1696),
.Y(n_1776)
);

AO22x2_ASAP7_75t_L g1777 ( 
.A1(n_1754),
.A2(n_1294),
.B1(n_1360),
.B2(n_1268),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1605),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1607),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1611),
.Y(n_1780)
);

NAND2xp33_ASAP7_75t_L g1781 ( 
.A(n_1720),
.B(n_1230),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1616),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1627),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1592),
.Y(n_1784)
);

NAND2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1747),
.B(n_944),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1631),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1638),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1602),
.A2(n_1214),
.B1(n_1216),
.B2(n_1209),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1639),
.Y(n_1789)
);

AO22x2_ASAP7_75t_L g1790 ( 
.A1(n_1612),
.A2(n_1589),
.B1(n_1650),
.B2(n_1596),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1597),
.Y(n_1791)
);

AO22x2_ASAP7_75t_L g1792 ( 
.A1(n_1758),
.A2(n_1360),
.B1(n_1268),
.B2(n_1006),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1593),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1644),
.A2(n_933),
.B1(n_1305),
.B2(n_1091),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1625),
.B(n_1227),
.Y(n_1795)
);

AO22x2_ASAP7_75t_L g1796 ( 
.A1(n_1624),
.A2(n_975),
.B1(n_989),
.B2(n_962),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1595),
.Y(n_1797)
);

NAND2x1p5_ASAP7_75t_L g1798 ( 
.A(n_1759),
.B(n_1000),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1629),
.A2(n_1226),
.B1(n_1243),
.B2(n_1225),
.C(n_1224),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1602),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1752),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1759),
.B(n_1250),
.Y(n_1802)
);

NOR2xp67_ASAP7_75t_L g1803 ( 
.A(n_1601),
.B(n_7),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1752),
.B(n_1206),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1698),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1667),
.A2(n_1247),
.B1(n_1253),
.B2(n_1252),
.C(n_1249),
.Y(n_1806)
);

CKINVDCx14_ASAP7_75t_R g1807 ( 
.A(n_1618),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1643),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1700),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1646),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1609),
.B(n_1751),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1701),
.Y(n_1812)
);

NAND2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1762),
.B(n_1296),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1600),
.B(n_1310),
.Y(n_1814)
);

AO22x2_ASAP7_75t_L g1815 ( 
.A1(n_1610),
.A2(n_1333),
.B1(n_1325),
.B2(n_1356),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1763),
.B(n_1765),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1702),
.Y(n_1817)
);

NAND2x1p5_ASAP7_75t_L g1818 ( 
.A(n_1740),
.B(n_1283),
.Y(n_1818)
);

AO22x2_ASAP7_75t_L g1819 ( 
.A1(n_1590),
.A2(n_1341),
.B1(n_1343),
.B2(n_1339),
.Y(n_1819)
);

AO22x2_ASAP7_75t_L g1820 ( 
.A1(n_1620),
.A2(n_1350),
.B1(n_1288),
.B2(n_1290),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1591),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1665),
.B(n_1262),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1717),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1703),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1682),
.B(n_950),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1652),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1654),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1658),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1661),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1710),
.A2(n_1279),
.B1(n_1284),
.B2(n_1276),
.C(n_1274),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1630),
.A2(n_1293),
.B1(n_1297),
.B2(n_1289),
.Y(n_1831)
);

BUFx8_ASAP7_75t_L g1832 ( 
.A(n_1739),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1632),
.A2(n_1301),
.B1(n_1302),
.B2(n_1299),
.Y(n_1833)
);

NAND2xp33_ASAP7_75t_L g1834 ( 
.A(n_1720),
.B(n_1315),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1621),
.A2(n_1323),
.B1(n_1326),
.B2(n_1318),
.C(n_1316),
.Y(n_1835)
);

AO22x2_ASAP7_75t_L g1836 ( 
.A1(n_1670),
.A2(n_1298),
.B1(n_1309),
.B2(n_1287),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1649),
.A2(n_1338),
.B1(n_1334),
.B2(n_934),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1618),
.A2(n_1322),
.B1(n_1328),
.B2(n_1311),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1761),
.B(n_951),
.Y(n_1839)
);

AO22x2_ASAP7_75t_L g1840 ( 
.A1(n_1768),
.A2(n_1332),
.B1(n_959),
.B2(n_967),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1687),
.Y(n_1841)
);

AO22x2_ASAP7_75t_L g1842 ( 
.A1(n_1768),
.A2(n_969),
.B1(n_976),
.B2(n_957),
.Y(n_1842)
);

AO22x2_ASAP7_75t_L g1843 ( 
.A1(n_1666),
.A2(n_992),
.B1(n_995),
.B2(n_982),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1750),
.B(n_1354),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1668),
.A2(n_1054),
.B1(n_1077),
.B2(n_981),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1745),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1587),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1746),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1675),
.B(n_996),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1636),
.B(n_1009),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1683),
.B(n_932),
.Y(n_1851)
);

AO22x2_ASAP7_75t_L g1852 ( 
.A1(n_1736),
.A2(n_1011),
.B1(n_1021),
.B2(n_1010),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1757),
.B(n_935),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1673),
.A2(n_1025),
.B(n_1026),
.C(n_1024),
.Y(n_1854)
);

AO22x2_ASAP7_75t_L g1855 ( 
.A1(n_1753),
.A2(n_1035),
.B1(n_1036),
.B2(n_1032),
.Y(n_1855)
);

AO22x2_ASAP7_75t_L g1856 ( 
.A1(n_1753),
.A2(n_1040),
.B1(n_1042),
.B2(n_1037),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1756),
.Y(n_1857)
);

NAND2x1p5_ASAP7_75t_L g1858 ( 
.A(n_1617),
.B(n_981),
.Y(n_1858)
);

AO22x2_ASAP7_75t_L g1859 ( 
.A1(n_1706),
.A2(n_1055),
.B1(n_1060),
.B2(n_1047),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1647),
.Y(n_1860)
);

AO22x2_ASAP7_75t_L g1861 ( 
.A1(n_1706),
.A2(n_1064),
.B1(n_1075),
.B2(n_1063),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1676),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1683),
.B(n_946),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1677),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1685),
.Y(n_1865)
);

NOR2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1671),
.B(n_954),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1721),
.B(n_1076),
.Y(n_1867)
);

AO22x2_ASAP7_75t_L g1868 ( 
.A1(n_1734),
.A2(n_1083),
.B1(n_1088),
.B2(n_1078),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1686),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1691),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1692),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1694),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1668),
.B(n_1634),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1724),
.B(n_1089),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1641),
.Y(n_1875)
);

AO22x2_ASAP7_75t_L g1876 ( 
.A1(n_1730),
.A2(n_1097),
.B1(n_1100),
.B2(n_1096),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1714),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1714),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1683),
.B(n_963),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1684),
.Y(n_1880)
);

AO22x2_ASAP7_75t_L g1881 ( 
.A1(n_1730),
.A2(n_1105),
.B1(n_1107),
.B2(n_1101),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1678),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1689),
.Y(n_1883)
);

BUFx8_ASAP7_75t_L g1884 ( 
.A(n_1727),
.Y(n_1884)
);

AO22x2_ASAP7_75t_L g1885 ( 
.A1(n_1727),
.A2(n_1110),
.B1(n_1111),
.B2(n_1108),
.Y(n_1885)
);

AO22x2_ASAP7_75t_L g1886 ( 
.A1(n_1738),
.A2(n_1118),
.B1(n_1119),
.B2(n_1116),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1594),
.B(n_1122),
.Y(n_1887)
);

AO22x2_ASAP7_75t_L g1888 ( 
.A1(n_1738),
.A2(n_1126),
.B1(n_1127),
.B2(n_1123),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1709),
.B(n_1131),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1723),
.Y(n_1890)
);

NAND2x1p5_ASAP7_75t_L g1891 ( 
.A(n_1623),
.B(n_1054),
.Y(n_1891)
);

AO22x2_ASAP7_75t_L g1892 ( 
.A1(n_1681),
.A2(n_1136),
.B1(n_1139),
.B2(n_1133),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1725),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1726),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1695),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1709),
.B(n_1143),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1713),
.Y(n_1897)
);

AO22x2_ASAP7_75t_L g1898 ( 
.A1(n_1715),
.A2(n_1146),
.B1(n_1149),
.B2(n_1144),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1603),
.B(n_1152),
.Y(n_1899)
);

AO22x2_ASAP7_75t_L g1900 ( 
.A1(n_1715),
.A2(n_1159),
.B1(n_1162),
.B2(n_1157),
.Y(n_1900)
);

AO22x2_ASAP7_75t_L g1901 ( 
.A1(n_1732),
.A2(n_1164),
.B1(n_1171),
.B2(n_1163),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1672),
.B(n_970),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1711),
.A2(n_977),
.B1(n_978),
.B2(n_974),
.C(n_971),
.Y(n_1903)
);

AO22x2_ASAP7_75t_L g1904 ( 
.A1(n_1737),
.A2(n_1183),
.B1(n_1192),
.B2(n_1175),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1613),
.B(n_1054),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1704),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1599),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1619),
.B(n_1655),
.Y(n_1908)
);

OAI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1731),
.A2(n_985),
.B1(n_994),
.B2(n_983),
.C(n_979),
.Y(n_1909)
);

OAI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1659),
.A2(n_1015),
.B1(n_1019),
.B2(n_1002),
.C(n_999),
.Y(n_1910)
);

AO22x2_ASAP7_75t_L g1911 ( 
.A1(n_1733),
.A2(n_1238),
.B1(n_1242),
.B2(n_1235),
.Y(n_1911)
);

AO22x2_ASAP7_75t_L g1912 ( 
.A1(n_1633),
.A2(n_1695),
.B1(n_1688),
.B2(n_1728),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1679),
.Y(n_1913)
);

OAI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1669),
.A2(n_1764),
.B1(n_1766),
.B2(n_1743),
.C(n_1742),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1693),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1690),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1697),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1719),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1728),
.A2(n_1033),
.B1(n_1039),
.B2(n_1030),
.Y(n_1919)
);

NAND2x1p5_ASAP7_75t_L g1920 ( 
.A(n_1640),
.B(n_1054),
.Y(n_1920)
);

AO22x2_ASAP7_75t_L g1921 ( 
.A1(n_1708),
.A2(n_1269),
.B1(n_1271),
.B2(n_1264),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1657),
.B(n_1354),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1653),
.B(n_1275),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1588),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1660),
.B(n_1281),
.Y(n_1925)
);

AO22x2_ASAP7_75t_L g1926 ( 
.A1(n_1664),
.A2(n_1307),
.B1(n_1327),
.B2(n_1282),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1767),
.Y(n_1927)
);

OR2x6_ASAP7_75t_L g1928 ( 
.A(n_1674),
.B(n_1014),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1656),
.B(n_1722),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1656),
.A2(n_1336),
.B1(n_1347),
.B2(n_1077),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1728),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1699),
.A2(n_1073),
.B1(n_1087),
.B2(n_1069),
.C(n_1051),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1729),
.A2(n_1098),
.B1(n_1099),
.B2(n_1094),
.Y(n_1933)
);

AO22x2_ASAP7_75t_L g1934 ( 
.A1(n_1718),
.A2(n_1017),
.B1(n_1031),
.B2(n_1014),
.Y(n_1934)
);

NAND2x1p5_ASAP7_75t_L g1935 ( 
.A(n_1662),
.B(n_1077),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1729),
.B(n_1113),
.Y(n_1936)
);

AO22x2_ASAP7_75t_L g1937 ( 
.A1(n_1622),
.A2(n_1031),
.B1(n_1050),
.B2(n_1017),
.Y(n_1937)
);

BUFx8_ASAP7_75t_L g1938 ( 
.A(n_1663),
.Y(n_1938)
);

AO22x2_ASAP7_75t_L g1939 ( 
.A1(n_1707),
.A2(n_1072),
.B1(n_1115),
.B2(n_1070),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1615),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1705),
.B(n_1114),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1604),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1628),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1680),
.A2(n_1124),
.B1(n_1129),
.B2(n_1128),
.Y(n_1944)
);

AO22x2_ASAP7_75t_L g1945 ( 
.A1(n_1716),
.A2(n_1132),
.B1(n_1167),
.B2(n_1115),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1705),
.B(n_1156),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1604),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1604),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1712),
.B(n_1161),
.Y(n_1949)
);

AO22x2_ASAP7_75t_L g1950 ( 
.A1(n_1606),
.A2(n_1229),
.B1(n_1280),
.B2(n_1184),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1651),
.B(n_1168),
.Y(n_1951)
);

OR2x2_ASAP7_75t_SL g1952 ( 
.A(n_1635),
.B(n_1280),
.Y(n_1952)
);

AO22x2_ASAP7_75t_L g1953 ( 
.A1(n_1637),
.A2(n_1342),
.B1(n_10),
.B2(n_8),
.Y(n_1953)
);

AO22x2_ASAP7_75t_L g1954 ( 
.A1(n_1744),
.A2(n_1342),
.B1(n_10),
.B2(n_8),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1642),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1645),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1648),
.Y(n_1957)
);

AO22x2_ASAP7_75t_L g1958 ( 
.A1(n_1749),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1651),
.B(n_1172),
.Y(n_1959)
);

AO22x2_ASAP7_75t_L g1960 ( 
.A1(n_1760),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1625),
.B(n_1186),
.Y(n_1961)
);

CKINVDCx11_ASAP7_75t_R g1962 ( 
.A(n_1626),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1598),
.Y(n_1963)
);

BUFx8_ASAP7_75t_L g1964 ( 
.A(n_1696),
.Y(n_1964)
);

AO22x2_ASAP7_75t_L g1965 ( 
.A1(n_1612),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1598),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1592),
.A2(n_1190),
.B1(n_1191),
.B2(n_1187),
.Y(n_1967)
);

OAI221xp5_ASAP7_75t_L g1968 ( 
.A1(n_1735),
.A2(n_1198),
.B1(n_1202),
.B2(n_1200),
.C(n_1195),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1592),
.A2(n_1204),
.B1(n_1210),
.B2(n_1203),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1747),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1625),
.B(n_1211),
.Y(n_1971)
);

AO22x2_ASAP7_75t_L g1972 ( 
.A1(n_1612),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1592),
.Y(n_1973)
);

AO22x2_ASAP7_75t_L g1974 ( 
.A1(n_1741),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1592),
.B(n_1219),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1616),
.Y(n_1976)
);

AO22x2_ASAP7_75t_L g1977 ( 
.A1(n_1741),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1977)
);

AO22x2_ASAP7_75t_L g1978 ( 
.A1(n_1741),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1978)
);

AO22x2_ASAP7_75t_L g1979 ( 
.A1(n_1741),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1979)
);

OAI22xp33_ASAP7_75t_SL g1980 ( 
.A1(n_1618),
.A2(n_1223),
.B1(n_1228),
.B2(n_1221),
.Y(n_1980)
);

AO22x2_ASAP7_75t_L g1981 ( 
.A1(n_1741),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1981)
);

NAND2x1p5_ASAP7_75t_L g1982 ( 
.A(n_1748),
.B(n_1117),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1811),
.B(n_1233),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_SL g1984 ( 
.A(n_1931),
.B(n_1117),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_SL g1985 ( 
.A(n_1824),
.B(n_1117),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1800),
.B(n_1345),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1973),
.B(n_1348),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1890),
.B(n_20),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1773),
.B(n_1355),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1810),
.B(n_1357),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1784),
.B(n_1358),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1771),
.B(n_1246),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1804),
.B(n_1324),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1788),
.B(n_1329),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1936),
.B(n_1248),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1970),
.B(n_1306),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1970),
.B(n_1308),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1893),
.B(n_1894),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1774),
.B(n_1251),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1772),
.B(n_1975),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1818),
.B(n_1313),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1832),
.B(n_1314),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1813),
.B(n_1317),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1822),
.B(n_1320),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1814),
.B(n_1254),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1873),
.B(n_1130),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1913),
.B(n_21),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1816),
.B(n_1915),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1801),
.B(n_1344),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1833),
.B(n_1353),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1919),
.B(n_1255),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1933),
.B(n_1267),
.Y(n_2012)
);

NAND2xp33_ASAP7_75t_SL g2013 ( 
.A(n_1940),
.B(n_1095),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1967),
.B(n_1272),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1969),
.B(n_1273),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1831),
.B(n_1277),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1785),
.B(n_1278),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1798),
.B(n_1285),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1803),
.B(n_1286),
.Y(n_2019)
);

NAND2xp33_ASAP7_75t_SL g2020 ( 
.A(n_1943),
.B(n_1095),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1769),
.B(n_1291),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1917),
.B(n_1826),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1841),
.B(n_1304),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1872),
.B(n_1837),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1941),
.B(n_1258),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1860),
.B(n_1312),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1827),
.B(n_1260),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1819),
.B(n_1261),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1828),
.B(n_1829),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1820),
.B(n_1265),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_SL g2031 ( 
.A(n_1805),
.B(n_1095),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1840),
.B(n_1775),
.Y(n_2032)
);

NAND2xp33_ASAP7_75t_SL g2033 ( 
.A(n_1809),
.B(n_1117),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_SL g2034 ( 
.A(n_1942),
.B(n_1130),
.Y(n_2034)
);

NAND2xp33_ASAP7_75t_SL g2035 ( 
.A(n_1916),
.B(n_1130),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1914),
.B(n_1844),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1884),
.B(n_1155),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_SL g2038 ( 
.A(n_1866),
.B(n_1331),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1918),
.B(n_22),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1815),
.B(n_1842),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1812),
.B(n_23),
.Y(n_2041)
);

NAND2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1823),
.B(n_1331),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1795),
.B(n_23),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1980),
.B(n_1166),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1902),
.B(n_1853),
.Y(n_2045)
);

NAND2xp33_ASAP7_75t_SL g2046 ( 
.A(n_1817),
.B(n_23),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1938),
.B(n_1240),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1895),
.B(n_1949),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_SL g2049 ( 
.A(n_1907),
.B(n_24),
.Y(n_2049)
);

NAND2xp33_ASAP7_75t_SL g2050 ( 
.A(n_1821),
.B(n_24),
.Y(n_2050)
);

NAND2xp33_ASAP7_75t_SL g2051 ( 
.A(n_1770),
.B(n_25),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1778),
.B(n_25),
.Y(n_2052)
);

NAND2xp33_ASAP7_75t_SL g2053 ( 
.A(n_1779),
.B(n_25),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_SL g2054 ( 
.A(n_1780),
.B(n_26),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1922),
.B(n_27),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1961),
.B(n_27),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1971),
.B(n_27),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1783),
.B(n_1786),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1944),
.B(n_28),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1867),
.B(n_28),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_SL g2061 ( 
.A(n_1787),
.B(n_26),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1874),
.B(n_30),
.Y(n_2062)
);

NAND2xp33_ASAP7_75t_SL g2063 ( 
.A(n_1789),
.B(n_29),
.Y(n_2063)
);

NAND2xp33_ASAP7_75t_SL g2064 ( 
.A(n_1963),
.B(n_29),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1908),
.B(n_31),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1825),
.B(n_31),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1966),
.B(n_29),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1839),
.B(n_32),
.Y(n_2068)
);

XNOR2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1794),
.B(n_32),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1791),
.B(n_33),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1886),
.B(n_33),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1858),
.B(n_34),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1891),
.B(n_36),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1793),
.B(n_35),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1889),
.B(n_36),
.Y(n_2075)
);

NAND2xp33_ASAP7_75t_SL g2076 ( 
.A(n_1947),
.B(n_35),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1896),
.B(n_36),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1886),
.B(n_1888),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1868),
.B(n_35),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1923),
.B(n_38),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1925),
.B(n_38),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_1928),
.B(n_37),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1797),
.B(n_37),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1951),
.B(n_40),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1959),
.B(n_40),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1875),
.B(n_41),
.Y(n_2086)
);

NAND2xp33_ASAP7_75t_SL g2087 ( 
.A(n_1948),
.B(n_39),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1911),
.B(n_41),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_1847),
.B(n_42),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1899),
.B(n_43),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1849),
.B(n_43),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1946),
.B(n_44),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1808),
.B(n_44),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1888),
.B(n_42),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1846),
.B(n_44),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1926),
.B(n_42),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1887),
.B(n_1920),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1935),
.B(n_46),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1850),
.B(n_46),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1848),
.B(n_47),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1857),
.B(n_47),
.Y(n_2101)
);

NAND2xp33_ASAP7_75t_SL g2102 ( 
.A(n_1865),
.B(n_45),
.Y(n_2102)
);

NAND2xp33_ASAP7_75t_SL g2103 ( 
.A(n_1869),
.B(n_45),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_SL g2104 ( 
.A(n_1870),
.B(n_45),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1871),
.B(n_49),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1928),
.B(n_48),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1982),
.B(n_50),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1930),
.B(n_51),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1905),
.B(n_51),
.Y(n_2109)
);

NAND2xp33_ASAP7_75t_SL g2110 ( 
.A(n_1782),
.B(n_49),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1885),
.B(n_52),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1862),
.B(n_52),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1877),
.B(n_55),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1878),
.B(n_55),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1882),
.B(n_56),
.Y(n_2115)
);

NAND2xp33_ASAP7_75t_SL g2116 ( 
.A(n_1781),
.B(n_52),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1864),
.B(n_56),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1883),
.B(n_57),
.Y(n_2118)
);

NAND2xp33_ASAP7_75t_SL g2119 ( 
.A(n_1834),
.B(n_56),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1897),
.B(n_58),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_SL g2121 ( 
.A(n_1906),
.B(n_58),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_1880),
.B(n_59),
.Y(n_2122)
);

NAND2xp33_ASAP7_75t_SL g2123 ( 
.A(n_1929),
.B(n_59),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1845),
.B(n_61),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1802),
.B(n_61),
.Y(n_2125)
);

NAND2xp33_ASAP7_75t_SL g2126 ( 
.A(n_1851),
.B(n_60),
.Y(n_2126)
);

NAND2xp33_ASAP7_75t_SL g2127 ( 
.A(n_1863),
.B(n_65),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1854),
.B(n_66),
.Y(n_2128)
);

NAND2xp33_ASAP7_75t_SL g2129 ( 
.A(n_1879),
.B(n_65),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1776),
.B(n_67),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1964),
.B(n_67),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1885),
.B(n_65),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1806),
.B(n_68),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1796),
.B(n_70),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1924),
.B(n_71),
.Y(n_2135)
);

NAND2xp33_ASAP7_75t_SL g2136 ( 
.A(n_1976),
.B(n_70),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1921),
.B(n_73),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1876),
.B(n_1881),
.Y(n_2138)
);

NAND2xp33_ASAP7_75t_SL g2139 ( 
.A(n_1955),
.B(n_73),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1927),
.B(n_74),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1956),
.B(n_74),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1876),
.B(n_73),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_SL g2143 ( 
.A(n_1957),
.B(n_75),
.Y(n_2143)
);

XNOR2xp5_ASAP7_75t_L g2144 ( 
.A(n_1777),
.B(n_75),
.Y(n_2144)
);

NAND2xp33_ASAP7_75t_SL g2145 ( 
.A(n_1912),
.B(n_76),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1945),
.B(n_76),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1799),
.B(n_79),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1838),
.B(n_80),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1881),
.B(n_78),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1807),
.B(n_80),
.Y(n_2150)
);

NAND2xp33_ASAP7_75t_SL g2151 ( 
.A(n_1912),
.B(n_78),
.Y(n_2151)
);

NAND2xp33_ASAP7_75t_SL g2152 ( 
.A(n_1859),
.B(n_80),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1861),
.B(n_82),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1855),
.B(n_1856),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1950),
.B(n_82),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1898),
.B(n_81),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1898),
.B(n_1900),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1900),
.B(n_81),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1950),
.B(n_83),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1830),
.B(n_83),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1835),
.B(n_83),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_1904),
.B(n_84),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1937),
.B(n_84),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1843),
.B(n_82),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1852),
.B(n_85),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1892),
.B(n_85),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1952),
.B(n_86),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_SL g2168 ( 
.A(n_1953),
.B(n_85),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1939),
.B(n_88),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1790),
.B(n_88),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1962),
.B(n_89),
.Y(n_2171)
);

AND2x4_ASAP7_75t_SL g2172 ( 
.A(n_1974),
.B(n_1977),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1932),
.B(n_89),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_1777),
.B(n_87),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1934),
.B(n_87),
.Y(n_2175)
);

NAND2xp33_ASAP7_75t_SL g2176 ( 
.A(n_1974),
.B(n_90),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1965),
.B(n_90),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1901),
.B(n_91),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1972),
.B(n_91),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1910),
.B(n_93),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1903),
.B(n_93),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1909),
.B(n_93),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1836),
.B(n_92),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1977),
.B(n_92),
.Y(n_2184)
);

NAND2xp33_ASAP7_75t_SL g2185 ( 
.A(n_1978),
.B(n_92),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1968),
.B(n_95),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_1978),
.B(n_94),
.Y(n_2187)
);

NAND2xp33_ASAP7_75t_SL g2188 ( 
.A(n_1979),
.B(n_95),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1981),
.B(n_97),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1981),
.B(n_1954),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1958),
.B(n_1960),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1792),
.B(n_99),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1800),
.B(n_100),
.Y(n_2193)
);

NAND2xp33_ASAP7_75t_SL g2194 ( 
.A(n_1931),
.B(n_96),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1800),
.B(n_100),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1800),
.B(n_101),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_1800),
.B(n_101),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1811),
.B(n_96),
.Y(n_2198)
);

NAND2xp33_ASAP7_75t_SL g2199 ( 
.A(n_1931),
.B(n_102),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1811),
.B(n_102),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1824),
.B(n_102),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1811),
.B(n_103),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1800),
.B(n_104),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_1800),
.B(n_104),
.Y(n_2204)
);

NAND2xp33_ASAP7_75t_SL g2205 ( 
.A(n_1931),
.B(n_103),
.Y(n_2205)
);

NAND2xp33_ASAP7_75t_SL g2206 ( 
.A(n_1931),
.B(n_104),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_SL g2207 ( 
.A(n_1800),
.B(n_106),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1800),
.B(n_106),
.Y(n_2208)
);

NAND2xp33_ASAP7_75t_SL g2209 ( 
.A(n_1931),
.B(n_105),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1824),
.B(n_107),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1800),
.B(n_108),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1824),
.B(n_107),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1800),
.B(n_108),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1800),
.B(n_109),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_SL g2215 ( 
.A(n_1931),
.B(n_107),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1824),
.B(n_109),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1824),
.B(n_109),
.Y(n_2217)
);

NAND2xp33_ASAP7_75t_SL g2218 ( 
.A(n_1931),
.B(n_110),
.Y(n_2218)
);

NAND2xp33_ASAP7_75t_SL g2219 ( 
.A(n_1931),
.B(n_111),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_1800),
.B(n_112),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1824),
.B(n_111),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1800),
.B(n_112),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1800),
.B(n_112),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_1800),
.B(n_113),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1824),
.B(n_111),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1800),
.B(n_114),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1800),
.B(n_114),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1800),
.B(n_114),
.Y(n_2228)
);

OR2x2_ASAP7_75t_L g2229 ( 
.A(n_1773),
.B(n_113),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_1800),
.B(n_116),
.Y(n_2230)
);

NAND2xp33_ASAP7_75t_SL g2231 ( 
.A(n_1931),
.B(n_115),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1800),
.B(n_117),
.Y(n_2232)
);

NAND2xp33_ASAP7_75t_SL g2233 ( 
.A(n_1931),
.B(n_116),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1824),
.B(n_117),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1824),
.B(n_117),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1824),
.B(n_118),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1824),
.B(n_119),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1824),
.B(n_119),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1800),
.B(n_121),
.Y(n_2239)
);

NAND2xp33_ASAP7_75t_SL g2240 ( 
.A(n_1931),
.B(n_120),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1800),
.B(n_122),
.Y(n_2241)
);

NAND2xp33_ASAP7_75t_SL g2242 ( 
.A(n_1931),
.B(n_120),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1811),
.B(n_120),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1824),
.B(n_122),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_1800),
.B(n_124),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_1800),
.B(n_124),
.Y(n_2246)
);

XNOR2x2_ASAP7_75t_L g2247 ( 
.A(n_1775),
.B(n_123),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1800),
.B(n_124),
.Y(n_2248)
);

NAND2xp33_ASAP7_75t_SL g2249 ( 
.A(n_1931),
.B(n_123),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_1800),
.B(n_126),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1800),
.B(n_126),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1800),
.B(n_126),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1800),
.B(n_127),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_1800),
.B(n_127),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_1800),
.B(n_128),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1811),
.B(n_125),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1824),
.B(n_128),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_1800),
.B(n_129),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1811),
.B(n_128),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_1800),
.B(n_130),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1824),
.B(n_129),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_SL g2262 ( 
.A(n_1931),
.B(n_129),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1824),
.B(n_130),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_1800),
.B(n_132),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1800),
.B(n_132),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1800),
.B(n_133),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_1800),
.B(n_133),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_1800),
.B(n_133),
.Y(n_2268)
);

AND2x2_ASAP7_75t_SL g2269 ( 
.A(n_1781),
.B(n_131),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_1800),
.B(n_135),
.Y(n_2270)
);

NAND2xp33_ASAP7_75t_SL g2271 ( 
.A(n_1931),
.B(n_134),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1824),
.B(n_134),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_1800),
.B(n_137),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1824),
.B(n_136),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1811),
.B(n_137),
.Y(n_2275)
);

NAND2xp33_ASAP7_75t_SL g2276 ( 
.A(n_1931),
.B(n_138),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_1811),
.B(n_138),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_1800),
.B(n_140),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1824),
.B(n_139),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1824),
.B(n_140),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1800),
.B(n_141),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1800),
.B(n_142),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1811),
.B(n_140),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_SL g2284 ( 
.A(n_1931),
.B(n_142),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_1800),
.B(n_144),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1824),
.B(n_143),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_1800),
.B(n_146),
.Y(n_2287)
);

NAND2xp33_ASAP7_75t_SL g2288 ( 
.A(n_1931),
.B(n_145),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1800),
.B(n_146),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_1800),
.B(n_148),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_1800),
.B(n_149),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1824),
.B(n_145),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1824),
.B(n_145),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_1824),
.B(n_149),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1811),
.B(n_150),
.Y(n_2295)
);

NAND2xp33_ASAP7_75t_SL g2296 ( 
.A(n_1931),
.B(n_150),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_1800),
.B(n_151),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_1800),
.B(n_152),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_SL g2299 ( 
.A(n_1931),
.B(n_150),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_1824),
.B(n_153),
.Y(n_2300)
);

AND2x2_ASAP7_75t_SL g2301 ( 
.A(n_1781),
.B(n_153),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_1800),
.B(n_154),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_1800),
.B(n_156),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_1800),
.B(n_156),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_1800),
.B(n_157),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_1800),
.B(n_157),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_SL g2307 ( 
.A(n_1931),
.B(n_155),
.Y(n_2307)
);

NAND2xp33_ASAP7_75t_SL g2308 ( 
.A(n_1931),
.B(n_155),
.Y(n_2308)
);

XNOR2xp5_ASAP7_75t_L g2309 ( 
.A(n_1823),
.B(n_157),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1800),
.B(n_159),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1824),
.B(n_158),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_1800),
.B(n_160),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_1800),
.B(n_160),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1824),
.B(n_158),
.Y(n_2314)
);

NAND2xp33_ASAP7_75t_SL g2315 ( 
.A(n_1931),
.B(n_161),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_1800),
.B(n_162),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_1800),
.B(n_163),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_1824),
.B(n_161),
.Y(n_2318)
);

NAND2xp33_ASAP7_75t_SL g2319 ( 
.A(n_1931),
.B(n_163),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_1800),
.B(n_165),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1824),
.B(n_164),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_1800),
.B(n_165),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_1800),
.B(n_165),
.Y(n_2323)
);

NAND2xp33_ASAP7_75t_SL g2324 ( 
.A(n_1931),
.B(n_164),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1824),
.B(n_166),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1800),
.B(n_167),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_1800),
.B(n_168),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_SL g2328 ( 
.A(n_1931),
.B(n_166),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_1773),
.B(n_166),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1824),
.B(n_168),
.Y(n_2330)
);

NAND2xp33_ASAP7_75t_SL g2331 ( 
.A(n_1931),
.B(n_168),
.Y(n_2331)
);

NAND2xp33_ASAP7_75t_SL g2332 ( 
.A(n_1931),
.B(n_169),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_1800),
.B(n_170),
.Y(n_2333)
);

NAND2xp33_ASAP7_75t_R g2334 ( 
.A(n_1976),
.B(n_169),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_1800),
.B(n_170),
.Y(n_2335)
);

NAND2xp33_ASAP7_75t_SL g2336 ( 
.A(n_1931),
.B(n_169),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_1811),
.B(n_170),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1811),
.B(n_171),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_1800),
.B(n_172),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1800),
.B(n_173),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_1800),
.B(n_173),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_1800),
.B(n_173),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1800),
.B(n_174),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_1824),
.B(n_171),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_1800),
.B(n_175),
.Y(n_2345)
);

NAND2xp33_ASAP7_75t_SL g2346 ( 
.A(n_1931),
.B(n_171),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_1800),
.B(n_177),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_1800),
.B(n_177),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1824),
.B(n_176),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_1811),
.B(n_178),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_SL g2351 ( 
.A(n_1931),
.B(n_178),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_1811),
.B(n_178),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_1811),
.B(n_179),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_1800),
.B(n_181),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_1800),
.B(n_182),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_1800),
.B(n_182),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1800),
.B(n_182),
.Y(n_2357)
);

NAND2xp33_ASAP7_75t_SL g2358 ( 
.A(n_1931),
.B(n_180),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_SL g2359 ( 
.A(n_1931),
.B(n_180),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_1800),
.B(n_183),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_1824),
.B(n_180),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1800),
.B(n_184),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_1800),
.B(n_185),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1824),
.B(n_183),
.Y(n_2364)
);

NAND2xp33_ASAP7_75t_SL g2365 ( 
.A(n_1931),
.B(n_183),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_1800),
.B(n_186),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_1800),
.B(n_186),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_1800),
.B(n_186),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_1800),
.B(n_187),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_1800),
.B(n_188),
.Y(n_2370)
);

NAND2xp33_ASAP7_75t_SL g2371 ( 
.A(n_1931),
.B(n_185),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1811),
.B(n_185),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1824),
.B(n_189),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_1811),
.B(n_189),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1824),
.B(n_190),
.Y(n_2375)
);

NAND2xp33_ASAP7_75t_SL g2376 ( 
.A(n_1931),
.B(n_191),
.Y(n_2376)
);

NAND2xp33_ASAP7_75t_SL g2377 ( 
.A(n_1931),
.B(n_191),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_1800),
.B(n_192),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1824),
.B(n_191),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_1800),
.B(n_193),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1824),
.B(n_192),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1824),
.B(n_193),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_1800),
.B(n_194),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_1824),
.B(n_193),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_1800),
.B(n_196),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1824),
.B(n_195),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_1800),
.B(n_196),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_1800),
.B(n_197),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_1800),
.B(n_197),
.Y(n_2389)
);

NAND2xp33_ASAP7_75t_SL g2390 ( 
.A(n_1931),
.B(n_195),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_1800),
.B(n_198),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_SL g2392 ( 
.A(n_1931),
.B(n_195),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_1800),
.B(n_200),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_1800),
.B(n_200),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_1800),
.B(n_200),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_1800),
.B(n_201),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_1800),
.B(n_201),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_1811),
.B(n_199),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1824),
.B(n_199),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_1800),
.B(n_203),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_1800),
.B(n_203),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_1800),
.B(n_203),
.Y(n_2402)
);

A2O1A1Ixp33_ASAP7_75t_L g2403 ( 
.A1(n_1985),
.A2(n_205),
.B(n_202),
.C(n_204),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1998),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2058),
.Y(n_2405)
);

OR2x6_ASAP7_75t_L g2406 ( 
.A(n_2138),
.B(n_202),
.Y(n_2406)
);

BUFx8_ASAP7_75t_L g2407 ( 
.A(n_2177),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_2210),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2210),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2013),
.A2(n_206),
.B(n_207),
.Y(n_2410)
);

NOR2xp67_ASAP7_75t_L g2411 ( 
.A(n_1993),
.B(n_208),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1998),
.Y(n_2412)
);

O2A1O1Ixp5_ASAP7_75t_L g2413 ( 
.A1(n_2020),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1998),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2008),
.B(n_208),
.Y(n_2415)
);

INVxp67_ASAP7_75t_L g2416 ( 
.A(n_2078),
.Y(n_2416)
);

CKINVDCx5p33_ASAP7_75t_R g2417 ( 
.A(n_2334),
.Y(n_2417)
);

INVx3_ASAP7_75t_L g2418 ( 
.A(n_2210),
.Y(n_2418)
);

OA21x2_ASAP7_75t_L g2419 ( 
.A1(n_2155),
.A2(n_2159),
.B(n_2191),
.Y(n_2419)
);

HB1xp67_ASAP7_75t_L g2420 ( 
.A(n_2216),
.Y(n_2420)
);

AO31x2_ASAP7_75t_L g2421 ( 
.A1(n_2146),
.A2(n_214),
.A3(n_212),
.B(n_213),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2216),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2000),
.B(n_215),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_2216),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2002),
.Y(n_2425)
);

AOI22xp5_ASAP7_75t_L g2426 ( 
.A1(n_2036),
.A2(n_218),
.B1(n_215),
.B2(n_216),
.Y(n_2426)
);

BUFx2_ASAP7_75t_L g2427 ( 
.A(n_2042),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2022),
.B(n_219),
.Y(n_2428)
);

AOI221xp5_ASAP7_75t_SL g2429 ( 
.A1(n_2190),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.C(n_223),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2294),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2052),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2198),
.B(n_226),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2052),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2200),
.B(n_227),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2398),
.B(n_227),
.Y(n_2435)
);

CKINVDCx16_ASAP7_75t_R g2436 ( 
.A(n_2069),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2082),
.Y(n_2437)
);

BUFx2_ASAP7_75t_L g2438 ( 
.A(n_2294),
.Y(n_2438)
);

NOR2xp67_ASAP7_75t_SL g2439 ( 
.A(n_2154),
.B(n_228),
.Y(n_2439)
);

A2O1A1Ixp33_ASAP7_75t_L g2440 ( 
.A1(n_2031),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_L g2441 ( 
.A(n_2045),
.B(n_231),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_2110),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_SL g2443 ( 
.A(n_2269),
.B(n_467),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2202),
.B(n_232),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2165),
.B(n_232),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2033),
.A2(n_233),
.B(n_234),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2029),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2067),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2243),
.B(n_235),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2269),
.B(n_467),
.Y(n_2450)
);

INVx5_ASAP7_75t_L g2451 ( 
.A(n_2294),
.Y(n_2451)
);

OAI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2201),
.A2(n_2217),
.B(n_2212),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2301),
.B(n_468),
.Y(n_2453)
);

INVxp67_ASAP7_75t_SL g2454 ( 
.A(n_2300),
.Y(n_2454)
);

NOR2xp67_ASAP7_75t_SL g2455 ( 
.A(n_2040),
.B(n_236),
.Y(n_2455)
);

NAND3xp33_ASAP7_75t_SL g2456 ( 
.A(n_2176),
.B(n_2188),
.C(n_2185),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2021),
.B(n_237),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2300),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2300),
.Y(n_2459)
);

INVxp67_ASAP7_75t_L g2460 ( 
.A(n_2229),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2256),
.B(n_237),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2259),
.B(n_237),
.Y(n_2462)
);

OAI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2221),
.A2(n_2234),
.B(n_2225),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_SL g2464 ( 
.A1(n_2173),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.C(n_241),
.Y(n_2464)
);

OA21x2_ASAP7_75t_L g2465 ( 
.A1(n_2162),
.A2(n_238),
.B(n_239),
.Y(n_2465)
);

OR2x6_ASAP7_75t_L g2466 ( 
.A(n_2361),
.B(n_238),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2361),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2275),
.B(n_239),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2111),
.B(n_240),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2041),
.Y(n_2470)
);

OAI21x1_ASAP7_75t_SL g2471 ( 
.A1(n_2157),
.A2(n_2247),
.B(n_2088),
.Y(n_2471)
);

OAI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2235),
.A2(n_242),
.B(n_243),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_2007),
.B(n_242),
.Y(n_2473)
);

BUFx3_ASAP7_75t_L g2474 ( 
.A(n_2361),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_2136),
.B(n_243),
.C(n_244),
.Y(n_2475)
);

O2A1O1Ixp5_ASAP7_75t_L g2476 ( 
.A1(n_2006),
.A2(n_247),
.B(n_244),
.C(n_246),
.Y(n_2476)
);

A2O1A1Ixp33_ASAP7_75t_L g2477 ( 
.A1(n_2049),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2007),
.B(n_248),
.Y(n_2478)
);

AO32x2_ASAP7_75t_L g2479 ( 
.A1(n_2168),
.A2(n_252),
.A3(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2277),
.B(n_2283),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2301),
.B(n_469),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2384),
.Y(n_2482)
);

BUFx10_ASAP7_75t_L g2483 ( 
.A(n_2384),
.Y(n_2483)
);

OAI21x1_ASAP7_75t_SL g2484 ( 
.A1(n_2166),
.A2(n_254),
.B(n_255),
.Y(n_2484)
);

OAI21x1_ASAP7_75t_SL g2485 ( 
.A1(n_2178),
.A2(n_2079),
.B(n_2156),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2295),
.B(n_254),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2236),
.A2(n_255),
.B(n_256),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_2384),
.Y(n_2488)
);

AND2x2_ASAP7_75t_SL g2489 ( 
.A(n_2172),
.B(n_257),
.Y(n_2489)
);

NOR2xp67_ASAP7_75t_L g2490 ( 
.A(n_1992),
.B(n_258),
.Y(n_2490)
);

INVx4_ASAP7_75t_L g2491 ( 
.A(n_2172),
.Y(n_2491)
);

INVx1_ASAP7_75t_SL g2492 ( 
.A(n_2329),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2132),
.B(n_259),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_1988),
.Y(n_2494)
);

INVx3_ASAP7_75t_L g2495 ( 
.A(n_1988),
.Y(n_2495)
);

AOI221xp5_ASAP7_75t_SL g2496 ( 
.A1(n_2180),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.C(n_264),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2089),
.Y(n_2497)
);

OAI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2237),
.A2(n_265),
.B(n_266),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_1984),
.B(n_470),
.Y(n_2499)
);

INVx2_ASAP7_75t_SL g2500 ( 
.A(n_2007),
.Y(n_2500)
);

NOR2x1_ASAP7_75t_L g2501 ( 
.A(n_2003),
.B(n_266),
.Y(n_2501)
);

OAI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_2238),
.A2(n_267),
.B(n_268),
.Y(n_2502)
);

A2O1A1Ixp33_ASAP7_75t_L g2503 ( 
.A1(n_2046),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_2503)
);

AO31x2_ASAP7_75t_L g2504 ( 
.A1(n_2070),
.A2(n_2096),
.A3(n_2137),
.B(n_2117),
.Y(n_2504)
);

OAI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_1988),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_2505)
);

OAI21xp5_ASAP7_75t_SL g2506 ( 
.A1(n_2144),
.A2(n_271),
.B(n_272),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2005),
.B(n_271),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2337),
.B(n_273),
.Y(n_2508)
);

BUFx2_ASAP7_75t_L g2509 ( 
.A(n_2034),
.Y(n_2509)
);

AOI221xp5_ASAP7_75t_SL g2510 ( 
.A1(n_2163),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2338),
.B(n_275),
.Y(n_2511)
);

AOI221xp5_ASAP7_75t_L g2512 ( 
.A1(n_2032),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.C(n_279),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2024),
.B(n_277),
.Y(n_2513)
);

CKINVDCx11_ASAP7_75t_R g2514 ( 
.A(n_2039),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2350),
.B(n_279),
.Y(n_2515)
);

OAI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2244),
.A2(n_280),
.B(n_281),
.Y(n_2516)
);

OAI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2039),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2352),
.B(n_2353),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2120),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2142),
.B(n_282),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2149),
.B(n_284),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_1984),
.A2(n_285),
.B(n_286),
.Y(n_2522)
);

AOI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2039),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2074),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2071),
.B(n_286),
.Y(n_2525)
);

OA21x2_ASAP7_75t_L g2526 ( 
.A1(n_2189),
.A2(n_288),
.B(n_289),
.Y(n_2526)
);

OR2x6_ASAP7_75t_L g2527 ( 
.A(n_2074),
.B(n_289),
.Y(n_2527)
);

INVx5_ASAP7_75t_L g2528 ( 
.A(n_2074),
.Y(n_2528)
);

OAI21xp5_ASAP7_75t_SL g2529 ( 
.A1(n_2134),
.A2(n_290),
.B(n_291),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2372),
.B(n_292),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2374),
.B(n_292),
.Y(n_2531)
);

OAI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2257),
.A2(n_293),
.B(n_294),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2083),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2133),
.B(n_295),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_1983),
.B(n_296),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2094),
.B(n_297),
.Y(n_2536)
);

NAND3xp33_ASAP7_75t_L g2537 ( 
.A(n_2145),
.B(n_2151),
.C(n_2143),
.Y(n_2537)
);

BUFx4_ASAP7_75t_SL g2538 ( 
.A(n_2130),
.Y(n_2538)
);

O2A1O1Ixp33_ASAP7_75t_SL g2539 ( 
.A1(n_2072),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2083),
.Y(n_2540)
);

OAI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2122),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2055),
.B(n_299),
.Y(n_2542)
);

INVx5_ASAP7_75t_L g2543 ( 
.A(n_2122),
.Y(n_2543)
);

OAI21xp5_ASAP7_75t_L g2544 ( 
.A1(n_2261),
.A2(n_301),
.B(n_302),
.Y(n_2544)
);

AOI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2152),
.A2(n_304),
.B1(n_301),
.B2(n_303),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2263),
.B(n_301),
.Y(n_2546)
);

O2A1O1Ixp5_ASAP7_75t_L g2547 ( 
.A1(n_2044),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_2122),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_2097),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2272),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2274),
.B(n_306),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2279),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2019),
.A2(n_2161),
.B(n_2160),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_2001),
.B(n_307),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2280),
.B(n_308),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2028),
.Y(n_2556)
);

OAI22x1_ASAP7_75t_L g2557 ( 
.A1(n_2184),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2557)
);

AO31x2_ASAP7_75t_L g2558 ( 
.A1(n_2112),
.A2(n_2175),
.A3(n_2292),
.B(n_2286),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_1994),
.B(n_312),
.Y(n_2559)
);

OAI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2293),
.A2(n_312),
.B(n_313),
.Y(n_2560)
);

A2O1A1Ixp33_ASAP7_75t_L g2561 ( 
.A1(n_2139),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_2311),
.B(n_315),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2314),
.B(n_316),
.Y(n_2563)
);

INVx2_ASAP7_75t_SL g2564 ( 
.A(n_2047),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2106),
.Y(n_2565)
);

AO32x2_ASAP7_75t_L g2566 ( 
.A1(n_2176),
.A2(n_2185),
.A3(n_2188),
.B1(n_2151),
.B2(n_2145),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2318),
.Y(n_2567)
);

NOR3xp33_ASAP7_75t_L g2568 ( 
.A(n_2148),
.B(n_318),
.C(n_319),
.Y(n_2568)
);

AOI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_2321),
.A2(n_319),
.B(n_320),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2325),
.A2(n_319),
.B(n_320),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2330),
.B(n_320),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_2073),
.Y(n_2572)
);

OAI21xp33_ASAP7_75t_L g2573 ( 
.A1(n_1999),
.A2(n_321),
.B(n_322),
.Y(n_2573)
);

AOI221x1_ASAP7_75t_L g2574 ( 
.A1(n_2152),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.C(n_324),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2344),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2349),
.B(n_322),
.Y(n_2576)
);

AOI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2364),
.A2(n_323),
.B(n_324),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2373),
.Y(n_2578)
);

INVx1_ASAP7_75t_SL g2579 ( 
.A(n_2076),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_1995),
.B(n_323),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_SL g2581 ( 
.A(n_2174),
.B(n_324),
.Y(n_2581)
);

CKINVDCx20_ASAP7_75t_R g2582 ( 
.A(n_2309),
.Y(n_2582)
);

NAND2x1p5_ASAP7_75t_L g2583 ( 
.A(n_2153),
.B(n_325),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2375),
.B(n_328),
.Y(n_2584)
);

OAI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2379),
.A2(n_328),
.B(n_329),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2381),
.Y(n_2586)
);

OAI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2382),
.A2(n_329),
.B(n_330),
.Y(n_2587)
);

CKINVDCx14_ASAP7_75t_R g2588 ( 
.A(n_2179),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2386),
.Y(n_2589)
);

NOR2x1_ASAP7_75t_L g2590 ( 
.A(n_2150),
.B(n_330),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2399),
.B(n_331),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2038),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2164),
.B(n_332),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2183),
.B(n_332),
.Y(n_2594)
);

NOR4xp25_ASAP7_75t_L g2595 ( 
.A(n_2192),
.B(n_336),
.C(n_334),
.D(n_335),
.Y(n_2595)
);

OR2x2_ASAP7_75t_L g2596 ( 
.A(n_2030),
.B(n_334),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2135),
.Y(n_2597)
);

A2O1A1Ixp33_ASAP7_75t_L g2598 ( 
.A1(n_2139),
.A2(n_337),
.B(n_335),
.C(n_336),
.Y(n_2598)
);

A2O1A1Ixp33_ASAP7_75t_L g2599 ( 
.A1(n_2143),
.A2(n_2119),
.B(n_2116),
.C(n_2053),
.Y(n_2599)
);

AOI221xp5_ASAP7_75t_SL g2600 ( 
.A1(n_2169),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.C(n_340),
.Y(n_2600)
);

BUFx12f_ASAP7_75t_L g2601 ( 
.A(n_2187),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2066),
.B(n_338),
.Y(n_2602)
);

BUFx6f_ASAP7_75t_L g2603 ( 
.A(n_2098),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2107),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2090),
.B(n_339),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2027),
.B(n_340),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2141),
.Y(n_2607)
);

NAND3x1_ASAP7_75t_L g2608 ( 
.A(n_2158),
.B(n_341),
.C(n_342),
.Y(n_2608)
);

OR2x2_ASAP7_75t_L g2609 ( 
.A(n_2068),
.B(n_342),
.Y(n_2609)
);

OAI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2181),
.A2(n_343),
.B(n_344),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2182),
.A2(n_343),
.B(n_344),
.Y(n_2611)
);

BUFx6f_ASAP7_75t_L g2612 ( 
.A(n_2109),
.Y(n_2612)
);

O2A1O1Ixp5_ASAP7_75t_L g2613 ( 
.A1(n_2092),
.A2(n_2085),
.B(n_2084),
.C(n_2167),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2194),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2199),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2035),
.B(n_475),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2037),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2043),
.B(n_345),
.Y(n_2618)
);

AOI21xp5_ASAP7_75t_SL g2619 ( 
.A1(n_2100),
.A2(n_346),
.B(n_347),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2060),
.B(n_347),
.Y(n_2620)
);

AOI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2186),
.A2(n_347),
.B(n_348),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_R g2622 ( 
.A(n_2205),
.B(n_349),
.Y(n_2622)
);

A2O1A1Ixp33_ASAP7_75t_L g2623 ( 
.A1(n_2051),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_2062),
.B(n_350),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2050),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2048),
.B(n_351),
.Y(n_2626)
);

NAND3xp33_ASAP7_75t_L g2627 ( 
.A(n_2054),
.B(n_354),
.C(n_355),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2075),
.B(n_354),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2205),
.B(n_475),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2077),
.B(n_2091),
.Y(n_2630)
);

AO21x1_ASAP7_75t_L g2631 ( 
.A1(n_2206),
.A2(n_478),
.B(n_476),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2056),
.B(n_355),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2065),
.A2(n_2059),
.B1(n_2128),
.B2(n_2101),
.Y(n_2633)
);

OAI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2147),
.A2(n_355),
.B(n_357),
.Y(n_2634)
);

BUFx12f_ASAP7_75t_L g2635 ( 
.A(n_2171),
.Y(n_2635)
);

AO32x2_ASAP7_75t_L g2636 ( 
.A1(n_2061),
.A2(n_360),
.A3(n_358),
.B1(n_359),
.B2(n_361),
.Y(n_2636)
);

AOI211x1_ASAP7_75t_L g2637 ( 
.A1(n_2193),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2113),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2099),
.B(n_363),
.Y(n_2639)
);

NAND2x1_ASAP7_75t_L g2640 ( 
.A(n_2206),
.B(n_364),
.Y(n_2640)
);

NAND2x1_ASAP7_75t_L g2641 ( 
.A(n_2209),
.B(n_364),
.Y(n_2641)
);

A2O1A1Ixp33_ASAP7_75t_L g2642 ( 
.A1(n_2063),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_2642)
);

OR2x2_ASAP7_75t_L g2643 ( 
.A(n_2080),
.B(n_366),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2195),
.B(n_368),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2196),
.B(n_368),
.Y(n_2645)
);

AOI22xp5_ASAP7_75t_L g2646 ( 
.A1(n_2102),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_SL g2647 ( 
.A(n_2209),
.B(n_369),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2081),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2014),
.B(n_369),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_SL g2650 ( 
.A(n_2215),
.B(n_370),
.Y(n_2650)
);

OAI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2114),
.A2(n_370),
.B(n_371),
.Y(n_2651)
);

INVxp67_ASAP7_75t_L g2652 ( 
.A(n_2087),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_SL g2653 ( 
.A(n_2215),
.B(n_2218),
.Y(n_2653)
);

BUFx6f_ASAP7_75t_L g2654 ( 
.A(n_2124),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2115),
.Y(n_2655)
);

AO31x2_ASAP7_75t_L g2656 ( 
.A1(n_2064),
.A2(n_374),
.A3(n_372),
.B(n_373),
.Y(n_2656)
);

CKINVDCx11_ASAP7_75t_R g2657 ( 
.A(n_2131),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2197),
.B(n_372),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2170),
.B(n_373),
.Y(n_2659)
);

AND2x4_ASAP7_75t_L g2660 ( 
.A(n_2057),
.B(n_374),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2093),
.B(n_374),
.Y(n_2661)
);

AOI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2140),
.A2(n_375),
.B(n_376),
.Y(n_2662)
);

OAI21x1_ASAP7_75t_SL g2663 ( 
.A1(n_2218),
.A2(n_375),
.B(n_376),
.Y(n_2663)
);

OAI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2118),
.A2(n_377),
.B(n_378),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2121),
.A2(n_378),
.B(n_379),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2105),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2219),
.B(n_479),
.Y(n_2667)
);

BUFx12f_ASAP7_75t_L g2668 ( 
.A(n_2025),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2103),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_2669)
);

A2O1A1Ixp33_ASAP7_75t_L g2670 ( 
.A1(n_2104),
.A2(n_386),
.B(n_384),
.C(n_385),
.Y(n_2670)
);

NAND3xp33_ASAP7_75t_L g2671 ( 
.A(n_2126),
.B(n_388),
.C(n_389),
.Y(n_2671)
);

INVx5_ASAP7_75t_L g2672 ( 
.A(n_2231),
.Y(n_2672)
);

NAND2x1p5_ASAP7_75t_L g2673 ( 
.A(n_2017),
.B(n_389),
.Y(n_2673)
);

AOI21xp33_ASAP7_75t_L g2674 ( 
.A1(n_2004),
.A2(n_390),
.B(n_391),
.Y(n_2674)
);

A2O1A1Ixp33_ASAP7_75t_L g2675 ( 
.A1(n_2231),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_2675)
);

NAND3xp33_ASAP7_75t_L g2676 ( 
.A(n_2127),
.B(n_392),
.C(n_393),
.Y(n_2676)
);

AOI22x1_ASAP7_75t_L g2677 ( 
.A1(n_2123),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_2677)
);

AND2x4_ASAP7_75t_L g2678 ( 
.A(n_2125),
.B(n_395),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2203),
.B(n_398),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2204),
.B(n_398),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_R g2681 ( 
.A(n_2233),
.B(n_2240),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2240),
.Y(n_2682)
);

NOR4xp25_ASAP7_75t_L g2683 ( 
.A(n_2207),
.B(n_401),
.C(n_399),
.D(n_400),
.Y(n_2683)
);

BUFx6f_ASAP7_75t_L g2684 ( 
.A(n_2108),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2208),
.Y(n_2685)
);

HB1xp67_ASAP7_75t_L g2686 ( 
.A(n_2211),
.Y(n_2686)
);

BUFx2_ASAP7_75t_L g2687 ( 
.A(n_2242),
.Y(n_2687)
);

OR2x2_ASAP7_75t_L g2688 ( 
.A(n_1991),
.B(n_1989),
.Y(n_2688)
);

AOI21xp5_ASAP7_75t_SL g2689 ( 
.A1(n_2213),
.A2(n_399),
.B(n_401),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2214),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2015),
.B(n_401),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2095),
.B(n_403),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2220),
.Y(n_2693)
);

OAI21xp5_ASAP7_75t_L g2694 ( 
.A1(n_2222),
.A2(n_405),
.B(n_406),
.Y(n_2694)
);

A2O1A1Ixp33_ASAP7_75t_L g2695 ( 
.A1(n_2242),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_2695)
);

BUFx2_ASAP7_75t_R g2696 ( 
.A(n_2016),
.Y(n_2696)
);

AO31x2_ASAP7_75t_L g2697 ( 
.A1(n_2249),
.A2(n_408),
.A3(n_406),
.B(n_407),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2018),
.Y(n_2698)
);

NAND2x1p5_ASAP7_75t_L g2699 ( 
.A(n_2086),
.B(n_2223),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2249),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_2224),
.Y(n_2701)
);

AND2x4_ASAP7_75t_L g2702 ( 
.A(n_1996),
.B(n_411),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2226),
.B(n_2227),
.Y(n_2703)
);

A2O1A1Ixp33_ASAP7_75t_L g2704 ( 
.A1(n_2262),
.A2(n_415),
.B(n_412),
.C(n_413),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2228),
.B(n_412),
.Y(n_2705)
);

INVx5_ASAP7_75t_L g2706 ( 
.A(n_2262),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2230),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2129),
.A2(n_413),
.B(n_416),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2232),
.B(n_416),
.Y(n_2709)
);

BUFx12f_ASAP7_75t_L g2710 ( 
.A(n_1997),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2239),
.B(n_417),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_L g2712 ( 
.A(n_2271),
.B(n_418),
.C(n_419),
.Y(n_2712)
);

BUFx4_ASAP7_75t_SL g2713 ( 
.A(n_2271),
.Y(n_2713)
);

BUFx2_ASAP7_75t_L g2714 ( 
.A(n_2276),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2241),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_2715)
);

BUFx4_ASAP7_75t_R g2716 ( 
.A(n_2276),
.Y(n_2716)
);

BUFx3_ASAP7_75t_L g2717 ( 
.A(n_2009),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_SL g2718 ( 
.A1(n_2245),
.A2(n_420),
.B(n_421),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2246),
.B(n_422),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2248),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2250),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2402),
.A2(n_422),
.B(n_423),
.Y(n_2722)
);

OAI21x1_ASAP7_75t_SL g2723 ( 
.A1(n_2284),
.A2(n_2296),
.B(n_2288),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2251),
.B(n_423),
.Y(n_2724)
);

OA21x2_ASAP7_75t_L g2725 ( 
.A1(n_2252),
.A2(n_2254),
.B(n_2253),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2255),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2401),
.A2(n_423),
.B(n_424),
.Y(n_2727)
);

OR2x2_ASAP7_75t_L g2728 ( 
.A(n_1990),
.B(n_424),
.Y(n_2728)
);

OAI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2258),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2260),
.B(n_2264),
.Y(n_2730)
);

AOI22x1_ASAP7_75t_L g2731 ( 
.A1(n_2284),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2400),
.B(n_425),
.Y(n_2732)
);

BUFx3_ASAP7_75t_L g2733 ( 
.A(n_2288),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2265),
.Y(n_2734)
);

BUFx2_ASAP7_75t_L g2735 ( 
.A(n_2299),
.Y(n_2735)
);

BUFx2_ASAP7_75t_L g2736 ( 
.A(n_2307),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2266),
.A2(n_427),
.B(n_428),
.Y(n_2737)
);

NAND3xp33_ASAP7_75t_L g2738 ( 
.A(n_2308),
.B(n_2319),
.C(n_2315),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2267),
.Y(n_2739)
);

OAI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2268),
.A2(n_427),
.B(n_428),
.Y(n_2740)
);

INVxp67_ASAP7_75t_SL g2741 ( 
.A(n_2270),
.Y(n_2741)
);

OAI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2273),
.A2(n_429),
.B(n_430),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2010),
.B(n_430),
.Y(n_2743)
);

BUFx8_ASAP7_75t_L g2744 ( 
.A(n_2315),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2278),
.Y(n_2745)
);

OAI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2281),
.A2(n_431),
.B(n_432),
.Y(n_2746)
);

OAI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2282),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2285),
.A2(n_436),
.B(n_437),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2287),
.B(n_437),
.Y(n_2749)
);

NOR4xp25_ASAP7_75t_L g2750 ( 
.A(n_2289),
.B(n_439),
.C(n_437),
.D(n_438),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2290),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2291),
.A2(n_438),
.B(n_439),
.Y(n_2752)
);

AOI211x1_ASAP7_75t_L g2753 ( 
.A1(n_2297),
.A2(n_442),
.B(n_440),
.C(n_441),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_2319),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_1986),
.B(n_442),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_1987),
.B(n_443),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2298),
.B(n_443),
.Y(n_2757)
);

INVx1_ASAP7_75t_SL g2758 ( 
.A(n_2023),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2324),
.B(n_484),
.Y(n_2759)
);

INVx1_ASAP7_75t_SL g2760 ( 
.A(n_2328),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2302),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2303),
.B(n_444),
.Y(n_2762)
);

OAI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2304),
.A2(n_2306),
.B(n_2305),
.Y(n_2763)
);

INVx2_ASAP7_75t_SL g2764 ( 
.A(n_2310),
.Y(n_2764)
);

NOR4xp25_ASAP7_75t_L g2765 ( 
.A(n_2312),
.B(n_447),
.C(n_445),
.D(n_446),
.Y(n_2765)
);

AO31x2_ASAP7_75t_L g2766 ( 
.A1(n_2328),
.A2(n_448),
.A3(n_445),
.B(n_447),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2313),
.B(n_448),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_SL g2768 ( 
.A(n_2331),
.B(n_448),
.Y(n_2768)
);

NOR4xp25_ASAP7_75t_L g2769 ( 
.A(n_2316),
.B(n_451),
.C(n_449),
.D(n_450),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2331),
.B(n_2332),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2332),
.B(n_485),
.Y(n_2771)
);

OAI21xp5_ASAP7_75t_L g2772 ( 
.A1(n_2317),
.A2(n_451),
.B(n_452),
.Y(n_2772)
);

AO32x2_ASAP7_75t_L g2773 ( 
.A1(n_2336),
.A2(n_454),
.A3(n_452),
.B1(n_453),
.B2(n_455),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2320),
.B(n_453),
.Y(n_2774)
);

OA21x2_ASAP7_75t_L g2775 ( 
.A1(n_2322),
.A2(n_454),
.B(n_455),
.Y(n_2775)
);

OAI21xp5_ASAP7_75t_L g2776 ( 
.A1(n_2613),
.A2(n_2326),
.B(n_2323),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2451),
.B(n_2327),
.Y(n_2777)
);

BUFx2_ASAP7_75t_SL g2778 ( 
.A(n_2491),
.Y(n_2778)
);

OAI21x1_ASAP7_75t_SL g2779 ( 
.A1(n_2723),
.A2(n_2346),
.B(n_2336),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2482),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2454),
.A2(n_2351),
.B(n_2346),
.Y(n_2781)
);

OA21x2_ASAP7_75t_L g2782 ( 
.A1(n_2537),
.A2(n_2335),
.B(n_2333),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2447),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2405),
.B(n_2339),
.Y(n_2784)
);

AOI221xp5_ASAP7_75t_L g2785 ( 
.A1(n_2595),
.A2(n_2342),
.B1(n_2343),
.B2(n_2341),
.C(n_2340),
.Y(n_2785)
);

AOI221xp5_ASAP7_75t_L g2786 ( 
.A1(n_2534),
.A2(n_2529),
.B1(n_2750),
.B2(n_2765),
.C(n_2683),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2405),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2466),
.A2(n_2358),
.B1(n_2359),
.B2(n_2351),
.Y(n_2788)
);

OAI21x1_ASAP7_75t_L g2789 ( 
.A1(n_2485),
.A2(n_2347),
.B(n_2345),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2469),
.B(n_2348),
.Y(n_2790)
);

AOI21xp33_ASAP7_75t_SL g2791 ( 
.A1(n_2489),
.A2(n_2385),
.B(n_2383),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2482),
.Y(n_2792)
);

INVx1_ASAP7_75t_SL g2793 ( 
.A(n_2514),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2493),
.B(n_2389),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2566),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2566),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2451),
.B(n_2354),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2566),
.Y(n_2798)
);

NAND3xp33_ASAP7_75t_L g2799 ( 
.A(n_2647),
.B(n_2768),
.C(n_2650),
.Y(n_2799)
);

HB1xp67_ASAP7_75t_L g2800 ( 
.A(n_2527),
.Y(n_2800)
);

OAI21x1_ASAP7_75t_L g2801 ( 
.A1(n_2614),
.A2(n_2356),
.B(n_2355),
.Y(n_2801)
);

CKINVDCx6p67_ASAP7_75t_R g2802 ( 
.A(n_2436),
.Y(n_2802)
);

OAI21x1_ASAP7_75t_L g2803 ( 
.A1(n_2614),
.A2(n_2360),
.B(n_2357),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2615),
.A2(n_2363),
.B(n_2362),
.Y(n_2804)
);

INVx8_ASAP7_75t_L g2805 ( 
.A(n_2466),
.Y(n_2805)
);

OAI21x1_ASAP7_75t_L g2806 ( 
.A1(n_2682),
.A2(n_2367),
.B(n_2366),
.Y(n_2806)
);

AO21x2_ASAP7_75t_L g2807 ( 
.A1(n_2471),
.A2(n_2369),
.B(n_2368),
.Y(n_2807)
);

AOI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2527),
.A2(n_2359),
.B1(n_2365),
.B2(n_2358),
.Y(n_2808)
);

NOR2xp67_ASAP7_75t_L g2809 ( 
.A(n_2672),
.B(n_2706),
.Y(n_2809)
);

NOR2xp67_ASAP7_75t_L g2810 ( 
.A(n_2672),
.B(n_2370),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2480),
.B(n_2378),
.Y(n_2811)
);

NOR2xp67_ASAP7_75t_L g2812 ( 
.A(n_2672),
.B(n_2380),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_2538),
.Y(n_2813)
);

AO21x2_ASAP7_75t_L g2814 ( 
.A1(n_2599),
.A2(n_2388),
.B(n_2387),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2518),
.B(n_2391),
.Y(n_2815)
);

OR2x2_ASAP7_75t_L g2816 ( 
.A(n_2492),
.B(n_2393),
.Y(n_2816)
);

AOI221xp5_ASAP7_75t_L g2817 ( 
.A1(n_2769),
.A2(n_2396),
.B1(n_2397),
.B2(n_2395),
.C(n_2394),
.Y(n_2817)
);

AND2x4_ASAP7_75t_L g2818 ( 
.A(n_2451),
.B(n_2011),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2575),
.Y(n_2819)
);

BUFx8_ASAP7_75t_SL g2820 ( 
.A(n_2635),
.Y(n_2820)
);

AO21x2_ASAP7_75t_L g2821 ( 
.A1(n_2663),
.A2(n_2012),
.B(n_2026),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2408),
.Y(n_2822)
);

AOI22xp33_ASAP7_75t_L g2823 ( 
.A1(n_2406),
.A2(n_2371),
.B1(n_2376),
.B2(n_2365),
.Y(n_2823)
);

AND2x4_ASAP7_75t_L g2824 ( 
.A(n_2528),
.B(n_2371),
.Y(n_2824)
);

O2A1O1Ixp33_ASAP7_75t_L g2825 ( 
.A1(n_2443),
.A2(n_2377),
.B(n_2390),
.C(n_2376),
.Y(n_2825)
);

INVx1_ASAP7_75t_SL g2826 ( 
.A(n_2528),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2406),
.A2(n_2390),
.B1(n_2392),
.B2(n_2377),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2578),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2499),
.A2(n_2653),
.B(n_2463),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2473),
.Y(n_2830)
);

NAND2x1p5_ASAP7_75t_L g2831 ( 
.A(n_2528),
.B(n_2392),
.Y(n_2831)
);

AOI21xp33_ASAP7_75t_SL g2832 ( 
.A1(n_2450),
.A2(n_455),
.B(n_456),
.Y(n_2832)
);

AOI22xp33_ASAP7_75t_L g2833 ( 
.A1(n_2456),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_2833)
);

AOI21x1_ASAP7_75t_L g2834 ( 
.A1(n_2592),
.A2(n_487),
.B(n_486),
.Y(n_2834)
);

AOI22xp33_ASAP7_75t_L g2835 ( 
.A1(n_2453),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_2835)
);

O2A1O1Ixp33_ASAP7_75t_L g2836 ( 
.A1(n_2481),
.A2(n_461),
.B(n_459),
.C(n_460),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2483),
.Y(n_2837)
);

BUFx3_ASAP7_75t_L g2838 ( 
.A(n_2710),
.Y(n_2838)
);

AOI22xp33_ASAP7_75t_L g2839 ( 
.A1(n_2491),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2483),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2520),
.B(n_459),
.Y(n_2841)
);

INVx2_ASAP7_75t_SL g2842 ( 
.A(n_2713),
.Y(n_2842)
);

OAI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2543),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2465),
.Y(n_2844)
);

OAI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2543),
.A2(n_465),
.B1(n_462),
.B2(n_464),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2581),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2465),
.Y(n_2847)
);

NAND5xp2_ASAP7_75t_SL g2848 ( 
.A(n_2417),
.B(n_493),
.C(n_491),
.D(n_492),
.E(n_494),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2697),
.Y(n_2849)
);

INVx3_ASAP7_75t_L g2850 ( 
.A(n_2408),
.Y(n_2850)
);

AOI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2452),
.A2(n_494),
.B(n_495),
.Y(n_2851)
);

OAI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2553),
.A2(n_497),
.B(n_498),
.Y(n_2852)
);

OAI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2413),
.A2(n_497),
.B(n_498),
.Y(n_2853)
);

AOI22xp33_ASAP7_75t_L g2854 ( 
.A1(n_2744),
.A2(n_501),
.B1(n_499),
.B2(n_500),
.Y(n_2854)
);

HB1xp67_ASAP7_75t_L g2855 ( 
.A(n_2473),
.Y(n_2855)
);

INVxp67_ASAP7_75t_SL g2856 ( 
.A(n_2420),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2697),
.Y(n_2857)
);

INVx8_ASAP7_75t_L g2858 ( 
.A(n_2543),
.Y(n_2858)
);

INVx4_ASAP7_75t_SL g2859 ( 
.A(n_2478),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2474),
.B(n_502),
.Y(n_2860)
);

AO21x2_ASAP7_75t_L g2861 ( 
.A1(n_2770),
.A2(n_502),
.B(n_503),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2697),
.Y(n_2862)
);

AO32x2_ASAP7_75t_L g2863 ( 
.A1(n_2409),
.A2(n_509),
.A3(n_507),
.B1(n_508),
.B2(n_511),
.Y(n_2863)
);

CKINVDCx20_ASAP7_75t_R g2864 ( 
.A(n_2657),
.Y(n_2864)
);

OAI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2611),
.A2(n_507),
.B(n_509),
.Y(n_2865)
);

BUFx8_ASAP7_75t_L g2866 ( 
.A(n_2668),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_L g2867 ( 
.A(n_2408),
.Y(n_2867)
);

INVxp67_ASAP7_75t_L g2868 ( 
.A(n_2423),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2521),
.B(n_512),
.Y(n_2869)
);

OA21x2_ASAP7_75t_L g2870 ( 
.A1(n_2738),
.A2(n_514),
.B(n_515),
.Y(n_2870)
);

OAI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2621),
.A2(n_516),
.B(n_517),
.Y(n_2871)
);

CKINVDCx6p67_ASAP7_75t_R g2872 ( 
.A(n_2601),
.Y(n_2872)
);

BUFx3_ASAP7_75t_L g2873 ( 
.A(n_2407),
.Y(n_2873)
);

AOI22x1_ASAP7_75t_L g2874 ( 
.A1(n_2410),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2766),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2525),
.B(n_521),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2766),
.Y(n_2877)
);

O2A1O1Ixp33_ASAP7_75t_L g2878 ( 
.A1(n_2475),
.A2(n_525),
.B(n_523),
.C(n_524),
.Y(n_2878)
);

OAI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2438),
.A2(n_528),
.B1(n_525),
.B2(n_526),
.Y(n_2879)
);

INVx3_ASAP7_75t_L g2880 ( 
.A(n_2424),
.Y(n_2880)
);

BUFx6f_ASAP7_75t_L g2881 ( 
.A(n_2424),
.Y(n_2881)
);

AOI21xp33_ASAP7_75t_L g2882 ( 
.A1(n_2633),
.A2(n_526),
.B(n_528),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2437),
.B(n_930),
.Y(n_2883)
);

BUFx6f_ASAP7_75t_L g2884 ( 
.A(n_2424),
.Y(n_2884)
);

INVx3_ASAP7_75t_L g2885 ( 
.A(n_2706),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2407),
.Y(n_2886)
);

AOI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2500),
.A2(n_529),
.B(n_530),
.Y(n_2887)
);

AO21x2_ASAP7_75t_L g2888 ( 
.A1(n_2484),
.A2(n_531),
.B(n_532),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2467),
.A2(n_532),
.B(n_533),
.Y(n_2889)
);

CKINVDCx20_ASAP7_75t_R g2890 ( 
.A(n_2582),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2766),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2412),
.B(n_2706),
.Y(n_2892)
);

OR2x6_ASAP7_75t_L g2893 ( 
.A(n_2478),
.B(n_533),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2656),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_L g2895 ( 
.A1(n_2744),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2552),
.B(n_929),
.Y(n_2896)
);

AO31x2_ASAP7_75t_L g2897 ( 
.A1(n_2631),
.A2(n_539),
.A3(n_536),
.B(n_537),
.Y(n_2897)
);

AOI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_2488),
.A2(n_537),
.B(n_540),
.Y(n_2898)
);

OAI21x1_ASAP7_75t_L g2899 ( 
.A1(n_2418),
.A2(n_2459),
.B(n_2458),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2656),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2536),
.B(n_542),
.Y(n_2901)
);

INVx3_ASAP7_75t_L g2902 ( 
.A(n_2548),
.Y(n_2902)
);

AOI21x1_ASAP7_75t_L g2903 ( 
.A1(n_2687),
.A2(n_546),
.B(n_547),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2556),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_2904)
);

OAI21xp5_ASAP7_75t_SL g2905 ( 
.A1(n_2506),
.A2(n_549),
.B(n_553),
.Y(n_2905)
);

CKINVDCx20_ASAP7_75t_R g2906 ( 
.A(n_2588),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2445),
.B(n_553),
.Y(n_2907)
);

NAND2x1p5_ASAP7_75t_L g2908 ( 
.A(n_2640),
.B(n_554),
.Y(n_2908)
);

INVxp33_ASAP7_75t_SL g2909 ( 
.A(n_2622),
.Y(n_2909)
);

OAI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2610),
.A2(n_554),
.B(n_555),
.Y(n_2910)
);

BUFx3_ASAP7_75t_L g2911 ( 
.A(n_2717),
.Y(n_2911)
);

INVx2_ASAP7_75t_SL g2912 ( 
.A(n_2548),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2568),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2714),
.A2(n_559),
.B1(n_556),
.B2(n_558),
.Y(n_2914)
);

AOI22xp33_ASAP7_75t_L g2915 ( 
.A1(n_2681),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_2915)
);

HB1xp67_ASAP7_75t_L g2916 ( 
.A(n_2548),
.Y(n_2916)
);

OAI21x1_ASAP7_75t_L g2917 ( 
.A1(n_2459),
.A2(n_2495),
.B(n_2494),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2442),
.Y(n_2918)
);

OR2x6_ASAP7_75t_L g2919 ( 
.A(n_2641),
.B(n_561),
.Y(n_2919)
);

BUFx3_ASAP7_75t_L g2920 ( 
.A(n_2698),
.Y(n_2920)
);

OA21x2_ASAP7_75t_L g2921 ( 
.A1(n_2574),
.A2(n_562),
.B(n_563),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2565),
.B(n_564),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2567),
.B(n_566),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2586),
.B(n_928),
.Y(n_2924)
);

INVx4_ASAP7_75t_L g2925 ( 
.A(n_2716),
.Y(n_2925)
);

AOI221xp5_ASAP7_75t_L g2926 ( 
.A1(n_2535),
.A2(n_570),
.B1(n_567),
.B2(n_569),
.C(n_571),
.Y(n_2926)
);

O2A1O1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_2648),
.A2(n_571),
.B(n_569),
.C(n_570),
.Y(n_2927)
);

AOI21xp33_ASAP7_75t_SL g2928 ( 
.A1(n_2557),
.A2(n_572),
.B(n_574),
.Y(n_2928)
);

INVx4_ASAP7_75t_L g2929 ( 
.A(n_2540),
.Y(n_2929)
);

OR2x6_ASAP7_75t_L g2930 ( 
.A(n_2689),
.B(n_572),
.Y(n_2930)
);

INVxp67_ASAP7_75t_SL g2931 ( 
.A(n_2540),
.Y(n_2931)
);

A2O1A1Ixp33_ASAP7_75t_L g2932 ( 
.A1(n_2522),
.A2(n_576),
.B(n_574),
.C(n_575),
.Y(n_2932)
);

AOI221xp5_ASAP7_75t_L g2933 ( 
.A1(n_2460),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.C(n_582),
.Y(n_2933)
);

AO31x2_ASAP7_75t_L g2934 ( 
.A1(n_2403),
.A2(n_585),
.A3(n_583),
.B(n_584),
.Y(n_2934)
);

AO32x2_ASAP7_75t_L g2935 ( 
.A1(n_2422),
.A2(n_589),
.A3(n_587),
.B1(n_588),
.B2(n_590),
.Y(n_2935)
);

BUFx3_ASAP7_75t_L g2936 ( 
.A(n_2425),
.Y(n_2936)
);

NAND3xp33_ASAP7_75t_L g2937 ( 
.A(n_2731),
.B(n_589),
.C(n_590),
.Y(n_2937)
);

BUFx2_ASAP7_75t_L g2938 ( 
.A(n_2733),
.Y(n_2938)
);

OAI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2547),
.A2(n_591),
.B(n_592),
.Y(n_2939)
);

BUFx3_ASAP7_75t_L g2940 ( 
.A(n_2702),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2735),
.A2(n_595),
.B1(n_591),
.B2(n_593),
.Y(n_2941)
);

AOI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2448),
.A2(n_595),
.B(n_596),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2754),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2416),
.B(n_596),
.Y(n_2944)
);

OR2x6_ASAP7_75t_SL g2945 ( 
.A(n_2596),
.B(n_597),
.Y(n_2945)
);

OAI22xp5_ASAP7_75t_L g2946 ( 
.A1(n_2736),
.A2(n_2760),
.B1(n_2523),
.B2(n_2700),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2526),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2589),
.B(n_597),
.Y(n_2948)
);

OR2x2_ASAP7_75t_L g2949 ( 
.A(n_2593),
.B(n_598),
.Y(n_2949)
);

INVx4_ASAP7_75t_L g2950 ( 
.A(n_2626),
.Y(n_2950)
);

OR2x2_ASAP7_75t_L g2951 ( 
.A(n_2594),
.B(n_600),
.Y(n_2951)
);

AO31x2_ASAP7_75t_L g2952 ( 
.A1(n_2440),
.A2(n_603),
.A3(n_601),
.B(n_602),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2696),
.B(n_601),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2526),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_L g2955 ( 
.A(n_2549),
.Y(n_2955)
);

OAI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2476),
.A2(n_605),
.B(n_606),
.Y(n_2956)
);

INVx1_ASAP7_75t_SL g2957 ( 
.A(n_2758),
.Y(n_2957)
);

INVx1_ASAP7_75t_SL g2958 ( 
.A(n_2688),
.Y(n_2958)
);

AO21x1_ASAP7_75t_L g2959 ( 
.A1(n_2629),
.A2(n_606),
.B(n_607),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2415),
.B(n_925),
.Y(n_2960)
);

CKINVDCx6p67_ASAP7_75t_R g2961 ( 
.A(n_2702),
.Y(n_2961)
);

AND2x4_ASAP7_75t_L g2962 ( 
.A(n_2404),
.B(n_2414),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2470),
.A2(n_609),
.B(n_610),
.Y(n_2963)
);

AOI21xp33_ASAP7_75t_L g2964 ( 
.A1(n_2741),
.A2(n_609),
.B(n_611),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2550),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_SL g2966 ( 
.A1(n_2731),
.A2(n_612),
.B(n_615),
.Y(n_2966)
);

AND2x6_ASAP7_75t_L g2967 ( 
.A(n_2497),
.B(n_615),
.Y(n_2967)
);

OR2x6_ASAP7_75t_L g2968 ( 
.A(n_2718),
.B(n_616),
.Y(n_2968)
);

AO21x2_ASAP7_75t_L g2969 ( 
.A1(n_2472),
.A2(n_924),
.B(n_616),
.Y(n_2969)
);

AND2x4_ASAP7_75t_L g2970 ( 
.A(n_2519),
.B(n_2524),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2579),
.A2(n_621),
.B1(n_617),
.B2(n_619),
.Y(n_2971)
);

INVx2_ASAP7_75t_SL g2972 ( 
.A(n_2626),
.Y(n_2972)
);

OR2x2_ASAP7_75t_L g2973 ( 
.A(n_2432),
.B(n_2434),
.Y(n_2973)
);

AO22x1_ASAP7_75t_L g2974 ( 
.A1(n_2590),
.A2(n_626),
.B1(n_623),
.B2(n_625),
.Y(n_2974)
);

HB1xp67_ASAP7_75t_L g2975 ( 
.A(n_2411),
.Y(n_2975)
);

NOR4xp25_ASAP7_75t_L g2976 ( 
.A(n_2608),
.B(n_629),
.C(n_627),
.D(n_628),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2479),
.Y(n_2977)
);

HB1xp67_ASAP7_75t_L g2978 ( 
.A(n_2490),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2435),
.B(n_631),
.Y(n_2979)
);

AOI221xp5_ASAP7_75t_SL g2980 ( 
.A1(n_2675),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.C(n_635),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2630),
.B(n_634),
.Y(n_2981)
);

NOR2x1_ASAP7_75t_R g2982 ( 
.A(n_2427),
.B(n_635),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2428),
.B(n_924),
.Y(n_2983)
);

BUFx3_ASAP7_75t_L g2984 ( 
.A(n_2549),
.Y(n_2984)
);

INVxp67_ASAP7_75t_SL g2985 ( 
.A(n_2431),
.Y(n_2985)
);

O2A1O1Ixp33_ASAP7_75t_SL g2986 ( 
.A1(n_2695),
.A2(n_2704),
.B(n_2503),
.C(n_2561),
.Y(n_2986)
);

CKINVDCx20_ASAP7_75t_R g2987 ( 
.A(n_2728),
.Y(n_2987)
);

INVx1_ASAP7_75t_SL g2988 ( 
.A(n_2509),
.Y(n_2988)
);

BUFx4_ASAP7_75t_R g2989 ( 
.A(n_2690),
.Y(n_2989)
);

CKINVDCx20_ASAP7_75t_R g2990 ( 
.A(n_2533),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2550),
.A2(n_643),
.B1(n_640),
.B2(n_642),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2479),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2441),
.B(n_640),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2661),
.B(n_2692),
.Y(n_2994)
);

AND2x4_ASAP7_75t_L g2995 ( 
.A(n_2433),
.B(n_642),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2562),
.B(n_2606),
.Y(n_2996)
);

OR2x2_ASAP7_75t_L g2997 ( 
.A(n_2444),
.B(n_644),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2562),
.B(n_923),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2479),
.Y(n_2999)
);

NAND3xp33_ASAP7_75t_L g3000 ( 
.A(n_2429),
.B(n_646),
.C(n_647),
.Y(n_3000)
);

OR2x6_ASAP7_75t_L g3001 ( 
.A(n_2637),
.B(n_648),
.Y(n_3001)
);

INVx1_ASAP7_75t_SL g3002 ( 
.A(n_2549),
.Y(n_3002)
);

OA21x2_ASAP7_75t_L g3003 ( 
.A1(n_2464),
.A2(n_652),
.B(n_654),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2513),
.A2(n_662),
.B1(n_660),
.B2(n_661),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2487),
.A2(n_664),
.B(n_665),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2419),
.Y(n_3006)
);

OAI222xp33_ASAP7_75t_L g3007 ( 
.A1(n_2455),
.A2(n_667),
.B1(n_669),
.B2(n_664),
.C1(n_665),
.C2(n_668),
.Y(n_3007)
);

A2O1A1Ixp33_ASAP7_75t_L g3008 ( 
.A1(n_2446),
.A2(n_670),
.B(n_667),
.C(n_669),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2609),
.B(n_670),
.Y(n_3009)
);

AO21x2_ASAP7_75t_L g3010 ( 
.A1(n_2498),
.A2(n_2516),
.B(n_2502),
.Y(n_3010)
);

OR2x2_ASAP7_75t_L g3011 ( 
.A(n_2449),
.B(n_671),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2659),
.B(n_673),
.Y(n_3012)
);

O2A1O1Ixp33_ASAP7_75t_SL g3013 ( 
.A1(n_2598),
.A2(n_2759),
.B(n_2771),
.C(n_2667),
.Y(n_3013)
);

NOR2xp67_ASAP7_75t_L g3014 ( 
.A(n_2712),
.B(n_673),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2673),
.Y(n_3015)
);

OR2x6_ASAP7_75t_L g3016 ( 
.A(n_2753),
.B(n_674),
.Y(n_3016)
);

BUFx2_ASAP7_75t_L g3017 ( 
.A(n_2652),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_2654),
.Y(n_3018)
);

AO31x2_ASAP7_75t_L g3019 ( 
.A1(n_2477),
.A2(n_678),
.A3(n_676),
.B(n_677),
.Y(n_3019)
);

CKINVDCx5p33_ASAP7_75t_R g3020 ( 
.A(n_2507),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2439),
.A2(n_682),
.B1(n_680),
.B2(n_681),
.Y(n_3021)
);

BUFx12f_ASAP7_75t_L g3022 ( 
.A(n_2617),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2686),
.B(n_923),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2421),
.Y(n_3024)
);

BUFx3_ASAP7_75t_L g3025 ( 
.A(n_2632),
.Y(n_3025)
);

INVx3_ASAP7_75t_L g3026 ( 
.A(n_2572),
.Y(n_3026)
);

AND2x4_ASAP7_75t_L g3027 ( 
.A(n_2597),
.B(n_683),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_2701),
.A2(n_687),
.B1(n_685),
.B2(n_686),
.Y(n_3028)
);

NAND2x1p5_ASAP7_75t_L g3029 ( 
.A(n_2501),
.B(n_688),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_2725),
.A2(n_691),
.B1(n_689),
.B2(n_690),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2607),
.B(n_692),
.Y(n_3031)
);

BUFx5_ASAP7_75t_L g3032 ( 
.A(n_2638),
.Y(n_3032)
);

OAI21x1_ASAP7_75t_SL g3033 ( 
.A1(n_2677),
.A2(n_693),
.B(n_694),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2504),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2461),
.B(n_922),
.Y(n_3035)
);

INVx3_ASAP7_75t_L g3036 ( 
.A(n_2572),
.Y(n_3036)
);

BUFx3_ASAP7_75t_L g3037 ( 
.A(n_2632),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_SL g3038 ( 
.A1(n_2583),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_3038)
);

OA21x2_ASAP7_75t_L g3039 ( 
.A1(n_2496),
.A2(n_2510),
.B(n_2600),
.Y(n_3039)
);

AOI221xp5_ASAP7_75t_L g3040 ( 
.A1(n_2457),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.C(n_702),
.Y(n_3040)
);

INVx3_ASAP7_75t_L g3041 ( 
.A(n_2572),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2775),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2504),
.Y(n_3043)
);

AO21x2_ASAP7_75t_L g3044 ( 
.A1(n_2532),
.A2(n_703),
.B(n_705),
.Y(n_3044)
);

NAND2xp33_ASAP7_75t_R g3045 ( 
.A(n_2660),
.B(n_706),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2725),
.A2(n_709),
.B1(n_707),
.B2(n_708),
.Y(n_3046)
);

HB1xp67_ASAP7_75t_L g3047 ( 
.A(n_2660),
.Y(n_3047)
);

BUFx2_ASAP7_75t_L g3048 ( 
.A(n_2678),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2504),
.Y(n_3049)
);

AND2x4_ASAP7_75t_L g3050 ( 
.A(n_2666),
.B(n_712),
.Y(n_3050)
);

CKINVDCx5p33_ASAP7_75t_R g3051 ( 
.A(n_2580),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2612),
.Y(n_3052)
);

INVx1_ASAP7_75t_SL g3053 ( 
.A(n_2684),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_2430),
.A2(n_718),
.B1(n_715),
.B2(n_717),
.Y(n_3054)
);

BUFx4f_ASAP7_75t_SL g3055 ( 
.A(n_2624),
.Y(n_3055)
);

AO21x2_ASAP7_75t_L g3056 ( 
.A1(n_2544),
.A2(n_2585),
.B(n_2560),
.Y(n_3056)
);

NAND3xp33_ASAP7_75t_L g3057 ( 
.A(n_2677),
.B(n_2627),
.C(n_2623),
.Y(n_3057)
);

OAI22xp33_ASAP7_75t_L g3058 ( 
.A1(n_2545),
.A2(n_718),
.B1(n_715),
.B2(n_717),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2636),
.Y(n_3059)
);

OAI211xp5_ASAP7_75t_SL g3060 ( 
.A1(n_2618),
.A2(n_722),
.B(n_719),
.C(n_721),
.Y(n_3060)
);

OAI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_2625),
.A2(n_724),
.B1(n_722),
.B2(n_723),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2462),
.B(n_725),
.Y(n_3062)
);

AOI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2505),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_3063)
);

CKINVDCx20_ASAP7_75t_R g3064 ( 
.A(n_2541),
.Y(n_3064)
);

INVx2_ASAP7_75t_SL g3065 ( 
.A(n_2628),
.Y(n_3065)
);

INVxp67_ASAP7_75t_L g3066 ( 
.A(n_2554),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2654),
.Y(n_3067)
);

A2O1A1Ixp33_ASAP7_75t_L g3068 ( 
.A1(n_2665),
.A2(n_729),
.B(n_726),
.C(n_728),
.Y(n_3068)
);

AO21x1_ASAP7_75t_L g3069 ( 
.A1(n_2517),
.A2(n_729),
.B(n_730),
.Y(n_3069)
);

A2O1A1Ixp33_ASAP7_75t_L g3070 ( 
.A1(n_2708),
.A2(n_2670),
.B(n_2642),
.C(n_2587),
.Y(n_3070)
);

OR2x2_ASAP7_75t_L g3071 ( 
.A(n_2468),
.B(n_730),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2546),
.A2(n_731),
.B(n_732),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2678),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2654),
.Y(n_3074)
);

O2A1O1Ixp33_ASAP7_75t_SL g3075 ( 
.A1(n_2616),
.A2(n_735),
.B(n_733),
.C(n_734),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2636),
.Y(n_3076)
);

OAI21x1_ASAP7_75t_SL g3077 ( 
.A1(n_2694),
.A2(n_736),
.B(n_737),
.Y(n_3077)
);

HB1xp67_ASAP7_75t_L g3078 ( 
.A(n_2643),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2486),
.B(n_922),
.Y(n_3079)
);

HB1xp67_ASAP7_75t_L g3080 ( 
.A(n_2508),
.Y(n_3080)
);

AND2x4_ASAP7_75t_L g3081 ( 
.A(n_2655),
.B(n_736),
.Y(n_3081)
);

OR2x2_ASAP7_75t_L g3082 ( 
.A(n_2511),
.B(n_738),
.Y(n_3082)
);

OR2x2_ASAP7_75t_L g3083 ( 
.A(n_2515),
.B(n_739),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2636),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_SL g3085 ( 
.A1(n_2573),
.A2(n_739),
.B(n_740),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_2755),
.Y(n_3086)
);

NOR2xp67_ASAP7_75t_L g3087 ( 
.A(n_2685),
.B(n_740),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2530),
.B(n_741),
.Y(n_3088)
);

OA21x2_ASAP7_75t_L g3089 ( 
.A1(n_2634),
.A2(n_741),
.B(n_742),
.Y(n_3089)
);

OAI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_2646),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2551),
.A2(n_744),
.B(n_745),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2558),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_2569),
.A2(n_746),
.B(n_747),
.Y(n_3093)
);

OAI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2763),
.A2(n_748),
.B(n_749),
.Y(n_3094)
);

INVxp33_ASAP7_75t_L g3095 ( 
.A(n_2531),
.Y(n_3095)
);

BUFx12f_ASAP7_75t_L g3096 ( 
.A(n_2603),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2555),
.A2(n_748),
.B(n_749),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2773),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2764),
.B(n_750),
.Y(n_3099)
);

BUFx2_ASAP7_75t_L g3100 ( 
.A(n_2612),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2756),
.B(n_750),
.Y(n_3101)
);

NAND3x1_ASAP7_75t_L g3102 ( 
.A(n_2426),
.B(n_751),
.C(n_753),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_2732),
.Y(n_3103)
);

BUFx2_ASAP7_75t_R g3104 ( 
.A(n_2620),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_2570),
.A2(n_751),
.B(n_754),
.Y(n_3105)
);

OAI21x1_ASAP7_75t_L g3106 ( 
.A1(n_2577),
.A2(n_755),
.B(n_756),
.Y(n_3106)
);

BUFx3_ASAP7_75t_L g3107 ( 
.A(n_2612),
.Y(n_3107)
);

OAI221xp5_ASAP7_75t_L g3108 ( 
.A1(n_2703),
.A2(n_755),
.B1(n_756),
.B2(n_757),
.C(n_758),
.Y(n_3108)
);

NAND2xp33_ASAP7_75t_L g3109 ( 
.A(n_2603),
.B(n_920),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2707),
.B(n_759),
.Y(n_3110)
);

O2A1O1Ixp33_ASAP7_75t_L g3111 ( 
.A1(n_2730),
.A2(n_762),
.B(n_760),
.C(n_761),
.Y(n_3111)
);

INVx3_ASAP7_75t_L g3112 ( 
.A(n_2603),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2684),
.Y(n_3113)
);

OAI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_2662),
.A2(n_2727),
.B(n_2722),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2684),
.Y(n_3115)
);

OR2x2_ASAP7_75t_L g3116 ( 
.A(n_2563),
.B(n_763),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2571),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_2602),
.Y(n_3118)
);

OAI221xp5_ASAP7_75t_L g3119 ( 
.A1(n_2740),
.A2(n_764),
.B1(n_765),
.B2(n_766),
.C(n_767),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_2576),
.A2(n_2591),
.B(n_2584),
.Y(n_3120)
);

BUFx3_ASAP7_75t_L g3121 ( 
.A(n_2604),
.Y(n_3121)
);

AND2x4_ASAP7_75t_L g3122 ( 
.A(n_2693),
.B(n_765),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_2559),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.Y(n_3123)
);

BUFx3_ASAP7_75t_L g3124 ( 
.A(n_2604),
.Y(n_3124)
);

OA21x2_ASAP7_75t_L g3125 ( 
.A1(n_2651),
.A2(n_768),
.B(n_769),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2539),
.Y(n_3126)
);

INVx3_ASAP7_75t_L g3127 ( 
.A(n_2604),
.Y(n_3127)
);

BUFx3_ASAP7_75t_L g3128 ( 
.A(n_2564),
.Y(n_3128)
);

BUFx12f_ASAP7_75t_L g3129 ( 
.A(n_2699),
.Y(n_3129)
);

INVx1_ASAP7_75t_SL g3130 ( 
.A(n_2639),
.Y(n_3130)
);

OAI221xp5_ASAP7_75t_L g3131 ( 
.A1(n_2742),
.A2(n_770),
.B1(n_772),
.B2(n_773),
.C(n_774),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2605),
.Y(n_3132)
);

AOI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_2720),
.A2(n_774),
.B(n_775),
.Y(n_3133)
);

AOI22x1_ASAP7_75t_L g3134 ( 
.A1(n_2737),
.A2(n_778),
.B1(n_775),
.B2(n_776),
.Y(n_3134)
);

NOR2x1_ASAP7_75t_L g3135 ( 
.A(n_2671),
.B(n_779),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2669),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2734),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2721),
.Y(n_3138)
);

AOI21x1_ASAP7_75t_L g3139 ( 
.A1(n_2726),
.A2(n_780),
.B(n_781),
.Y(n_3139)
);

OAI22xp33_ASAP7_75t_L g3140 ( 
.A1(n_2676),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_3140)
);

OA21x2_ASAP7_75t_L g3141 ( 
.A1(n_2664),
.A2(n_784),
.B(n_785),
.Y(n_3141)
);

NAND2xp33_ASAP7_75t_L g3142 ( 
.A(n_2805),
.B(n_2746),
.Y(n_3142)
);

INVx2_ASAP7_75t_SL g3143 ( 
.A(n_2866),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2894),
.Y(n_3144)
);

BUFx6f_ASAP7_75t_L g3145 ( 
.A(n_2858),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2841),
.B(n_784),
.Y(n_3146)
);

CKINVDCx5p33_ASAP7_75t_R g3147 ( 
.A(n_2866),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2894),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2900),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2783),
.B(n_2542),
.Y(n_3150)
);

CKINVDCx8_ASAP7_75t_R g3151 ( 
.A(n_2813),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2819),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2900),
.Y(n_3153)
);

INVx2_ASAP7_75t_SL g3154 ( 
.A(n_2873),
.Y(n_3154)
);

BUFx12f_ASAP7_75t_L g3155 ( 
.A(n_2842),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2868),
.B(n_2644),
.Y(n_3156)
);

BUFx6f_ASAP7_75t_L g3157 ( 
.A(n_2858),
.Y(n_3157)
);

INVx2_ASAP7_75t_SL g3158 ( 
.A(n_2886),
.Y(n_3158)
);

OR2x6_ASAP7_75t_L g3159 ( 
.A(n_2805),
.B(n_2619),
.Y(n_3159)
);

HB1xp67_ASAP7_75t_L g3160 ( 
.A(n_2830),
.Y(n_3160)
);

AO21x2_ASAP7_75t_L g3161 ( 
.A1(n_2966),
.A2(n_2752),
.B(n_2748),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2828),
.Y(n_3162)
);

OR2x6_ASAP7_75t_L g3163 ( 
.A(n_2805),
.B(n_2772),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2849),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2849),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2907),
.B(n_785),
.Y(n_3166)
);

INVx2_ASAP7_75t_SL g3167 ( 
.A(n_2838),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2994),
.B(n_2869),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2787),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2857),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2857),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2862),
.Y(n_3172)
);

AND2x2_ASAP7_75t_L g3173 ( 
.A(n_2876),
.B(n_786),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2862),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_3137),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3138),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3138),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2875),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2909),
.B(n_2649),
.Y(n_3179)
);

INVx3_ASAP7_75t_L g3180 ( 
.A(n_2858),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2875),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2877),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2877),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2911),
.Y(n_3184)
);

AND2x2_ASAP7_75t_L g3185 ( 
.A(n_2901),
.B(n_787),
.Y(n_3185)
);

INVx4_ASAP7_75t_L g3186 ( 
.A(n_2859),
.Y(n_3186)
);

BUFx2_ASAP7_75t_L g3187 ( 
.A(n_2925),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2891),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_2820),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2891),
.Y(n_3190)
);

NAND2x1p5_ASAP7_75t_L g3191 ( 
.A(n_2793),
.B(n_2739),
.Y(n_3191)
);

BUFx10_ASAP7_75t_L g3192 ( 
.A(n_2893),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2949),
.B(n_788),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2951),
.B(n_788),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3078),
.B(n_2512),
.Y(n_3195)
);

BUFx3_ASAP7_75t_L g3196 ( 
.A(n_2906),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_3117),
.Y(n_3197)
);

HB1xp67_ASAP7_75t_L g3198 ( 
.A(n_2855),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_2859),
.B(n_2745),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3103),
.Y(n_3200)
);

OR2x2_ASAP7_75t_L g3201 ( 
.A(n_2958),
.B(n_2645),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3118),
.Y(n_3202)
);

INVx2_ASAP7_75t_SL g3203 ( 
.A(n_2872),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2995),
.Y(n_3204)
);

OR2x6_ASAP7_75t_L g3205 ( 
.A(n_2778),
.B(n_2925),
.Y(n_3205)
);

HB1xp67_ASAP7_75t_L g3206 ( 
.A(n_3048),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2995),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_SL g3208 ( 
.A(n_3104),
.B(n_2674),
.Y(n_3208)
);

AND2x4_ASAP7_75t_L g3209 ( 
.A(n_2809),
.B(n_2751),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3027),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_3080),
.B(n_789),
.Y(n_3211)
);

BUFx2_ASAP7_75t_L g3212 ( 
.A(n_3096),
.Y(n_3212)
);

INVxp67_ASAP7_75t_SL g3213 ( 
.A(n_2985),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3027),
.Y(n_3214)
);

HB1xp67_ASAP7_75t_L g3215 ( 
.A(n_3073),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3095),
.B(n_2893),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_2802),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_3129),
.Y(n_3218)
);

OR2x6_ASAP7_75t_L g3219 ( 
.A(n_2919),
.B(n_2715),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3031),
.Y(n_3220)
);

BUFx3_ASAP7_75t_L g3221 ( 
.A(n_2864),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3031),
.Y(n_3222)
);

NAND3xp33_ASAP7_75t_L g3223 ( 
.A(n_2786),
.B(n_2691),
.C(n_2743),
.Y(n_3223)
);

CKINVDCx5p33_ASAP7_75t_R g3224 ( 
.A(n_2890),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_3047),
.Y(n_3225)
);

BUFx3_ASAP7_75t_L g3226 ( 
.A(n_2920),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3050),
.Y(n_3227)
);

AND2x2_ASAP7_75t_L g3228 ( 
.A(n_2961),
.B(n_789),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3050),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3081),
.Y(n_3230)
);

BUFx6f_ASAP7_75t_L g3231 ( 
.A(n_2822),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3081),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3122),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2844),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3122),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3065),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_3055),
.B(n_2658),
.Y(n_3237)
);

INVx2_ASAP7_75t_SL g3238 ( 
.A(n_2936),
.Y(n_3238)
);

HB1xp67_ASAP7_75t_L g3239 ( 
.A(n_2800),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2844),
.Y(n_3240)
);

HB1xp67_ASAP7_75t_L g3241 ( 
.A(n_2940),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3136),
.B(n_2996),
.Y(n_3242)
);

NAND2x1p5_ASAP7_75t_L g3243 ( 
.A(n_2860),
.B(n_2761),
.Y(n_3243)
);

BUFx3_ASAP7_75t_L g3244 ( 
.A(n_3022),
.Y(n_3244)
);

OAI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_2799),
.A2(n_2747),
.B(n_2729),
.Y(n_3245)
);

NAND4xp25_ASAP7_75t_L g3246 ( 
.A(n_3045),
.B(n_2679),
.C(n_2705),
.D(n_2680),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2847),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_2847),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2947),
.Y(n_3249)
);

INVx3_ASAP7_75t_L g3250 ( 
.A(n_2885),
.Y(n_3250)
);

AND2x4_ASAP7_75t_L g3251 ( 
.A(n_2809),
.B(n_2709),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3066),
.B(n_790),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2947),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_2990),
.A2(n_2719),
.B1(n_2724),
.B2(n_2711),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_2954),
.Y(n_3255)
);

CKINVDCx5p33_ASAP7_75t_R g3256 ( 
.A(n_2918),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3017),
.Y(n_3257)
);

BUFx2_ASAP7_75t_L g3258 ( 
.A(n_2938),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3001),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_3006),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3006),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3001),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3012),
.B(n_790),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3016),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3016),
.Y(n_3265)
);

INVxp67_ASAP7_75t_R g3266 ( 
.A(n_3038),
.Y(n_3266)
);

OR2x2_ASAP7_75t_L g3267 ( 
.A(n_2957),
.B(n_2749),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2780),
.Y(n_3268)
);

BUFx3_ASAP7_75t_L g3269 ( 
.A(n_3128),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_3015),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2896),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_L g3272 ( 
.A1(n_3064),
.A2(n_2774),
.B1(n_2762),
.B2(n_2767),
.Y(n_3272)
);

NAND2x1p5_ASAP7_75t_L g3273 ( 
.A(n_2860),
.B(n_2757),
.Y(n_3273)
);

INVx1_ASAP7_75t_SL g3274 ( 
.A(n_2989),
.Y(n_3274)
);

INVx3_ASAP7_75t_L g3275 ( 
.A(n_2780),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2790),
.B(n_919),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_2987),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_L g3278 ( 
.A1(n_3136),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.Y(n_3278)
);

AND2x4_ASAP7_75t_L g3279 ( 
.A(n_2824),
.B(n_791),
.Y(n_3279)
);

INVx1_ASAP7_75t_SL g3280 ( 
.A(n_2826),
.Y(n_3280)
);

BUFx2_ASAP7_75t_L g3281 ( 
.A(n_2950),
.Y(n_3281)
);

CKINVDCx5p33_ASAP7_75t_R g3282 ( 
.A(n_2945),
.Y(n_3282)
);

OR2x2_ASAP7_75t_L g3283 ( 
.A(n_2950),
.B(n_795),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_2794),
.B(n_795),
.Y(n_3284)
);

BUFx4f_ASAP7_75t_SL g3285 ( 
.A(n_3025),
.Y(n_3285)
);

INVxp67_ASAP7_75t_SL g3286 ( 
.A(n_2799),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_2824),
.B(n_797),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2923),
.Y(n_3288)
);

OR2x2_ASAP7_75t_L g3289 ( 
.A(n_2856),
.B(n_798),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_2944),
.B(n_801),
.Y(n_3290)
);

OA21x2_ASAP7_75t_L g3291 ( 
.A1(n_3024),
.A2(n_801),
.B(n_802),
.Y(n_3291)
);

BUFx2_ASAP7_75t_L g3292 ( 
.A(n_3037),
.Y(n_3292)
);

BUFx3_ASAP7_75t_L g3293 ( 
.A(n_3107),
.Y(n_3293)
);

BUFx3_ASAP7_75t_L g3294 ( 
.A(n_3121),
.Y(n_3294)
);

BUFx3_ASAP7_75t_L g3295 ( 
.A(n_3124),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2972),
.B(n_802),
.Y(n_3296)
);

INVx1_ASAP7_75t_SL g3297 ( 
.A(n_2826),
.Y(n_3297)
);

BUFx2_ASAP7_75t_L g3298 ( 
.A(n_2792),
.Y(n_3298)
);

INVxp67_ASAP7_75t_L g3299 ( 
.A(n_2982),
.Y(n_3299)
);

BUFx3_ASAP7_75t_L g3300 ( 
.A(n_2792),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3092),
.Y(n_3301)
);

BUFx6f_ASAP7_75t_L g3302 ( 
.A(n_2822),
.Y(n_3302)
);

BUFx2_ASAP7_75t_SL g3303 ( 
.A(n_2943),
.Y(n_3303)
);

OR2x2_ASAP7_75t_L g3304 ( 
.A(n_2973),
.B(n_803),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_2943),
.B(n_803),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3130),
.B(n_918),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3092),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3034),
.Y(n_3308)
);

INVx3_ASAP7_75t_L g3309 ( 
.A(n_2831),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3034),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3043),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3043),
.Y(n_3312)
);

INVx3_ASAP7_75t_L g3313 ( 
.A(n_2929),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3049),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3049),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2795),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2784),
.B(n_804),
.Y(n_3317)
);

INVx4_ASAP7_75t_L g3318 ( 
.A(n_2837),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_2823),
.A2(n_807),
.B1(n_805),
.B2(n_806),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2924),
.Y(n_3320)
);

AO21x1_ASAP7_75t_SL g3321 ( 
.A1(n_2788),
.A2(n_805),
.B(n_807),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2948),
.Y(n_3322)
);

INVx2_ASAP7_75t_SL g3323 ( 
.A(n_2840),
.Y(n_3323)
);

BUFx3_ASAP7_75t_L g3324 ( 
.A(n_2840),
.Y(n_3324)
);

BUFx3_ASAP7_75t_L g3325 ( 
.A(n_2984),
.Y(n_3325)
);

AND2x4_ASAP7_75t_L g3326 ( 
.A(n_2929),
.B(n_808),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2934),
.Y(n_3327)
);

AOI22xp33_ASAP7_75t_L g3328 ( 
.A1(n_2827),
.A2(n_2808),
.B1(n_2968),
.B2(n_2930),
.Y(n_3328)
);

BUFx12f_ASAP7_75t_L g3329 ( 
.A(n_3020),
.Y(n_3329)
);

INVx3_ASAP7_75t_L g3330 ( 
.A(n_2892),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3132),
.B(n_808),
.Y(n_3331)
);

OAI21x1_ASAP7_75t_SL g3332 ( 
.A1(n_2779),
.A2(n_809),
.B(n_810),
.Y(n_3332)
);

AOI21x1_ASAP7_75t_L g3333 ( 
.A1(n_2829),
.A2(n_811),
.B(n_812),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2934),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2934),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2952),
.Y(n_3336)
);

HB1xp67_ASAP7_75t_L g3337 ( 
.A(n_2988),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_2905),
.A2(n_811),
.B1(n_812),
.B2(n_813),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_2811),
.B(n_814),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2952),
.Y(n_3340)
);

OA21x2_ASAP7_75t_L g3341 ( 
.A1(n_3042),
.A2(n_815),
.B(n_817),
.Y(n_3341)
);

AOI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_2781),
.A2(n_818),
.B(n_819),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2952),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_2988),
.B(n_818),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_2892),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3009),
.B(n_918),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3019),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3019),
.Y(n_3348)
);

OR2x2_ASAP7_75t_L g3349 ( 
.A(n_2816),
.B(n_821),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_2922),
.B(n_821),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2815),
.B(n_822),
.Y(n_3351)
);

NAND2x1p5_ASAP7_75t_L g3352 ( 
.A(n_2846),
.B(n_2818),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_2998),
.B(n_822),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3019),
.Y(n_3354)
);

AO21x2_ASAP7_75t_L g3355 ( 
.A1(n_3033),
.A2(n_823),
.B(n_824),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_2982),
.Y(n_3356)
);

BUFx3_ASAP7_75t_L g3357 ( 
.A(n_3100),
.Y(n_3357)
);

BUFx2_ASAP7_75t_L g3358 ( 
.A(n_2822),
.Y(n_3358)
);

OA21x2_ASAP7_75t_L g3359 ( 
.A1(n_3059),
.A2(n_823),
.B(n_825),
.Y(n_3359)
);

BUFx12f_ASAP7_75t_L g3360 ( 
.A(n_3051),
.Y(n_3360)
);

BUFx3_ASAP7_75t_L g3361 ( 
.A(n_2867),
.Y(n_3361)
);

INVx2_ASAP7_75t_SL g3362 ( 
.A(n_2919),
.Y(n_3362)
);

HB1xp67_ASAP7_75t_L g3363 ( 
.A(n_2916),
.Y(n_3363)
);

AND2x4_ASAP7_75t_L g3364 ( 
.A(n_2850),
.B(n_825),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2967),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_2846),
.B(n_917),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2967),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_2867),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_2967),
.Y(n_3369)
);

OA21x2_ASAP7_75t_L g3370 ( 
.A1(n_3059),
.A2(n_3084),
.B(n_3076),
.Y(n_3370)
);

OAI21x1_ASAP7_75t_SL g3371 ( 
.A1(n_2905),
.A2(n_826),
.B(n_827),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_2930),
.A2(n_826),
.B1(n_827),
.B2(n_828),
.Y(n_3372)
);

BUFx6f_ASAP7_75t_L g3373 ( 
.A(n_2867),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_2883),
.B(n_828),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_2881),
.Y(n_3375)
);

OR2x6_ASAP7_75t_L g3376 ( 
.A(n_2968),
.B(n_2908),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_2981),
.B(n_2979),
.Y(n_3377)
);

INVx3_ASAP7_75t_L g3378 ( 
.A(n_2881),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_2997),
.B(n_916),
.Y(n_3379)
);

INVx2_ASAP7_75t_SL g3380 ( 
.A(n_2975),
.Y(n_3380)
);

BUFx2_ASAP7_75t_L g3381 ( 
.A(n_2881),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_2977),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2897),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2977),
.Y(n_3384)
);

HB1xp67_ASAP7_75t_L g3385 ( 
.A(n_2884),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3011),
.B(n_831),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_3071),
.B(n_831),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_2897),
.Y(n_3388)
);

INVx3_ASAP7_75t_L g3389 ( 
.A(n_2884),
.Y(n_3389)
);

BUFx2_ASAP7_75t_L g3390 ( 
.A(n_2884),
.Y(n_3390)
);

HB1xp67_ASAP7_75t_SL g3391 ( 
.A(n_2978),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2992),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2992),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_2999),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_2999),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3115),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_2897),
.Y(n_3397)
);

AO21x2_ASAP7_75t_L g3398 ( 
.A1(n_2937),
.A2(n_3014),
.B(n_2852),
.Y(n_3398)
);

OR2x6_ASAP7_75t_L g3399 ( 
.A(n_2974),
.B(n_3029),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_2962),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3076),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2962),
.Y(n_3402)
);

HB1xp67_ASAP7_75t_L g3403 ( 
.A(n_2912),
.Y(n_3403)
);

BUFx2_ASAP7_75t_L g3404 ( 
.A(n_2850),
.Y(n_3404)
);

INVx2_ASAP7_75t_SL g3405 ( 
.A(n_2880),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3082),
.B(n_832),
.Y(n_3406)
);

INVx1_ASAP7_75t_SL g3407 ( 
.A(n_3086),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2795),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2796),
.Y(n_3409)
);

HB1xp67_ASAP7_75t_L g3410 ( 
.A(n_3113),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_2825),
.A2(n_833),
.B(n_834),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2796),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2798),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2798),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3098),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3098),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3084),
.Y(n_3417)
);

INVx3_ASAP7_75t_L g3418 ( 
.A(n_2777),
.Y(n_3418)
);

BUFx4f_ASAP7_75t_SL g3419 ( 
.A(n_3002),
.Y(n_3419)
);

BUFx3_ASAP7_75t_L g3420 ( 
.A(n_2880),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3083),
.B(n_916),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3032),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3099),
.B(n_833),
.Y(n_3423)
);

INVx2_ASAP7_75t_SL g3424 ( 
.A(n_2902),
.Y(n_3424)
);

O2A1O1Ixp33_ASAP7_75t_SL g3425 ( 
.A1(n_3007),
.A2(n_834),
.B(n_835),
.C(n_836),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3032),
.Y(n_3426)
);

INVx4_ASAP7_75t_SL g3427 ( 
.A(n_3038),
.Y(n_3427)
);

HB1xp67_ASAP7_75t_L g3428 ( 
.A(n_3113),
.Y(n_3428)
);

BUFx2_ASAP7_75t_L g3429 ( 
.A(n_2902),
.Y(n_3429)
);

INVx3_ASAP7_75t_L g3430 ( 
.A(n_2777),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3116),
.B(n_915),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_2993),
.B(n_837),
.Y(n_3432)
);

INVx2_ASAP7_75t_SL g3433 ( 
.A(n_3026),
.Y(n_3433)
);

AND2x4_ASAP7_75t_L g3434 ( 
.A(n_2931),
.B(n_838),
.Y(n_3434)
);

INVx3_ASAP7_75t_L g3435 ( 
.A(n_2797),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3101),
.B(n_839),
.Y(n_3436)
);

HB1xp67_ASAP7_75t_L g3437 ( 
.A(n_3053),
.Y(n_3437)
);

OR2x2_ASAP7_75t_L g3438 ( 
.A(n_3023),
.B(n_840),
.Y(n_3438)
);

NOR2xp67_ASAP7_75t_SL g3439 ( 
.A(n_3085),
.B(n_841),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3053),
.Y(n_3440)
);

BUFx10_ASAP7_75t_L g3441 ( 
.A(n_2953),
.Y(n_3441)
);

HB1xp67_ASAP7_75t_L g3442 ( 
.A(n_3002),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3120),
.B(n_841),
.Y(n_3443)
);

HB1xp67_ASAP7_75t_L g3444 ( 
.A(n_3026),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3035),
.B(n_915),
.Y(n_3445)
);

BUFx4f_ASAP7_75t_SL g3446 ( 
.A(n_2955),
.Y(n_3446)
);

AO21x2_ASAP7_75t_L g3447 ( 
.A1(n_3014),
.A2(n_842),
.B(n_843),
.Y(n_3447)
);

AND2x4_ASAP7_75t_L g3448 ( 
.A(n_2970),
.B(n_842),
.Y(n_3448)
);

HB1xp67_ASAP7_75t_L g3449 ( 
.A(n_3036),
.Y(n_3449)
);

BUFx4f_ASAP7_75t_SL g3450 ( 
.A(n_2955),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2946),
.A2(n_843),
.B1(n_844),
.B2(n_845),
.Y(n_3451)
);

OAI21x1_ASAP7_75t_L g3452 ( 
.A1(n_2899),
.A2(n_844),
.B(n_846),
.Y(n_3452)
);

CKINVDCx20_ASAP7_75t_R g3453 ( 
.A(n_3189),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_3147),
.Y(n_3454)
);

INVxp67_ASAP7_75t_L g3455 ( 
.A(n_3258),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3202),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_R g3457 ( 
.A(n_3143),
.B(n_2848),
.Y(n_3457)
);

NAND2xp33_ASAP7_75t_R g3458 ( 
.A(n_3282),
.B(n_2791),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3197),
.B(n_2976),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_SL g3460 ( 
.A(n_3274),
.B(n_2976),
.Y(n_3460)
);

XNOR2xp5_ASAP7_75t_L g3461 ( 
.A(n_3224),
.B(n_3102),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3200),
.Y(n_3462)
);

NAND2xp33_ASAP7_75t_R g3463 ( 
.A(n_3356),
.B(n_2791),
.Y(n_3463)
);

OR2x6_ASAP7_75t_L g3464 ( 
.A(n_3205),
.B(n_3376),
.Y(n_3464)
);

AND2x4_ASAP7_75t_L g3465 ( 
.A(n_3205),
.B(n_3036),
.Y(n_3465)
);

AND2x4_ASAP7_75t_L g3466 ( 
.A(n_3186),
.B(n_3041),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_R g3467 ( 
.A(n_3151),
.B(n_2903),
.Y(n_3467)
);

AND2x4_ASAP7_75t_L g3468 ( 
.A(n_3186),
.B(n_3041),
.Y(n_3468)
);

INVxp67_ASAP7_75t_L g3469 ( 
.A(n_3391),
.Y(n_3469)
);

OR2x6_ASAP7_75t_L g3470 ( 
.A(n_3376),
.B(n_3303),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_R g3471 ( 
.A(n_3218),
.B(n_2834),
.Y(n_3471)
);

NAND2xp33_ASAP7_75t_R g3472 ( 
.A(n_3187),
.B(n_2870),
.Y(n_3472)
);

NAND2xp33_ASAP7_75t_R g3473 ( 
.A(n_3212),
.B(n_2870),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3176),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3177),
.Y(n_3475)
);

AND2x4_ASAP7_75t_L g3476 ( 
.A(n_3281),
.B(n_3052),
.Y(n_3476)
);

AND2x4_ASAP7_75t_SL g3477 ( 
.A(n_3145),
.B(n_2818),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_SL g3478 ( 
.A(n_3318),
.B(n_2810),
.Y(n_3478)
);

XNOR2xp5_ASAP7_75t_L g3479 ( 
.A(n_3217),
.B(n_2854),
.Y(n_3479)
);

NAND2x1p5_ASAP7_75t_L g3480 ( 
.A(n_3145),
.B(n_3054),
.Y(n_3480)
);

OR2x2_ASAP7_75t_L g3481 ( 
.A(n_3337),
.B(n_3052),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3168),
.B(n_2970),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_R g3483 ( 
.A(n_3203),
.B(n_3109),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3242),
.B(n_3010),
.Y(n_3484)
);

INVxp67_ASAP7_75t_L g3485 ( 
.A(n_3239),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_3145),
.B(n_3112),
.Y(n_3486)
);

AND2x4_ASAP7_75t_L g3487 ( 
.A(n_3157),
.B(n_3112),
.Y(n_3487)
);

NOR2xp33_ASAP7_75t_R g3488 ( 
.A(n_3256),
.B(n_2895),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3257),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3152),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_3269),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3236),
.B(n_3127),
.Y(n_3492)
);

NAND2xp33_ASAP7_75t_R g3493 ( 
.A(n_3180),
.B(n_3125),
.Y(n_3493)
);

NAND2xp33_ASAP7_75t_R g3494 ( 
.A(n_3180),
.B(n_3125),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3169),
.Y(n_3495)
);

INVxp67_ASAP7_75t_L g3496 ( 
.A(n_3216),
.Y(n_3496)
);

NAND2xp33_ASAP7_75t_R g3497 ( 
.A(n_3228),
.B(n_3141),
.Y(n_3497)
);

BUFx24_ASAP7_75t_SL g3498 ( 
.A(n_3254),
.Y(n_3498)
);

AND2x4_ASAP7_75t_L g3499 ( 
.A(n_3157),
.B(n_3127),
.Y(n_3499)
);

INVxp67_ASAP7_75t_L g3500 ( 
.A(n_3241),
.Y(n_3500)
);

XNOR2xp5_ASAP7_75t_L g3501 ( 
.A(n_3221),
.B(n_3196),
.Y(n_3501)
);

BUFx10_ASAP7_75t_L g3502 ( 
.A(n_3157),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3162),
.B(n_3010),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3213),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3280),
.Y(n_3505)
);

NAND2xp33_ASAP7_75t_R g3506 ( 
.A(n_3399),
.B(n_3141),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3297),
.B(n_2888),
.Y(n_3507)
);

BUFx3_ASAP7_75t_L g3508 ( 
.A(n_3226),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3160),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3175),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3198),
.Y(n_3511)
);

BUFx10_ASAP7_75t_L g3512 ( 
.A(n_3167),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3396),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3225),
.Y(n_3514)
);

BUFx12f_ASAP7_75t_L g3515 ( 
.A(n_3155),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_R g3516 ( 
.A(n_3192),
.B(n_846),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3206),
.B(n_3215),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_R g3518 ( 
.A(n_3192),
.B(n_848),
.Y(n_3518)
);

CKINVDCx20_ASAP7_75t_R g3519 ( 
.A(n_3244),
.Y(n_3519)
);

BUFx3_ASAP7_75t_L g3520 ( 
.A(n_3184),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3146),
.B(n_2888),
.Y(n_3521)
);

NAND2xp33_ASAP7_75t_R g3522 ( 
.A(n_3399),
.B(n_2921),
.Y(n_3522)
);

CKINVDCx16_ASAP7_75t_R g3523 ( 
.A(n_3329),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3417),
.Y(n_3524)
);

OR2x6_ASAP7_75t_L g3525 ( 
.A(n_3159),
.B(n_2810),
.Y(n_3525)
);

INVxp67_ASAP7_75t_L g3526 ( 
.A(n_3298),
.Y(n_3526)
);

BUFx3_ASAP7_75t_L g3527 ( 
.A(n_3154),
.Y(n_3527)
);

NAND2xp33_ASAP7_75t_R g3528 ( 
.A(n_3279),
.B(n_2921),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3417),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3271),
.B(n_3056),
.Y(n_3530)
);

CKINVDCx6p67_ASAP7_75t_R g3531 ( 
.A(n_3360),
.Y(n_3531)
);

AND2x4_ASAP7_75t_L g3532 ( 
.A(n_3313),
.B(n_2812),
.Y(n_3532)
);

INVx2_ASAP7_75t_SL g3533 ( 
.A(n_3158),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_R g3534 ( 
.A(n_3142),
.B(n_848),
.Y(n_3534)
);

INVxp67_ASAP7_75t_L g3535 ( 
.A(n_3363),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3288),
.B(n_3056),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3407),
.B(n_3299),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3260),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3415),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_R g3540 ( 
.A(n_3285),
.B(n_3208),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3415),
.Y(n_3541)
);

CKINVDCx12_ASAP7_75t_R g3542 ( 
.A(n_3163),
.Y(n_3542)
);

CKINVDCx16_ASAP7_75t_R g3543 ( 
.A(n_3277),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3261),
.Y(n_3544)
);

NAND2xp33_ASAP7_75t_R g3545 ( 
.A(n_3279),
.B(n_3089),
.Y(n_3545)
);

NAND2x1p5_ASAP7_75t_L g3546 ( 
.A(n_3326),
.B(n_3054),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3320),
.B(n_2928),
.Y(n_3547)
);

AND2x4_ASAP7_75t_L g3548 ( 
.A(n_3313),
.B(n_2812),
.Y(n_3548)
);

NAND2xp33_ASAP7_75t_R g3549 ( 
.A(n_3287),
.B(n_3089),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3401),
.Y(n_3550)
);

INVxp67_ASAP7_75t_L g3551 ( 
.A(n_3304),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3322),
.B(n_2928),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3276),
.B(n_2861),
.Y(n_3553)
);

NAND2xp33_ASAP7_75t_R g3554 ( 
.A(n_3287),
.B(n_3039),
.Y(n_3554)
);

NAND2xp33_ASAP7_75t_R g3555 ( 
.A(n_3163),
.B(n_3039),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3301),
.Y(n_3556)
);

AND2x4_ASAP7_75t_L g3557 ( 
.A(n_3300),
.B(n_2797),
.Y(n_3557)
);

NAND2xp33_ASAP7_75t_R g3558 ( 
.A(n_3326),
.B(n_3309),
.Y(n_3558)
);

NAND2xp33_ASAP7_75t_R g3559 ( 
.A(n_3309),
.B(n_2832),
.Y(n_3559)
);

NOR2xp33_ASAP7_75t_R g3560 ( 
.A(n_3362),
.B(n_849),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3230),
.B(n_2980),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_R g3562 ( 
.A(n_3419),
.B(n_850),
.Y(n_3562)
);

NOR2x1_ASAP7_75t_L g3563 ( 
.A(n_3318),
.B(n_3000),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3284),
.B(n_3400),
.Y(n_3564)
);

BUFx3_ASAP7_75t_L g3565 ( 
.A(n_3238),
.Y(n_3565)
);

BUFx3_ASAP7_75t_L g3566 ( 
.A(n_3270),
.Y(n_3566)
);

NAND2xp33_ASAP7_75t_R g3567 ( 
.A(n_3159),
.B(n_2832),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_R g3568 ( 
.A(n_3259),
.B(n_850),
.Y(n_3568)
);

INVxp67_ASAP7_75t_L g3569 ( 
.A(n_3211),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3232),
.B(n_2980),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3301),
.Y(n_3571)
);

NAND2xp33_ASAP7_75t_R g3572 ( 
.A(n_3305),
.B(n_3003),
.Y(n_3572)
);

NAND2xp33_ASAP7_75t_SL g3573 ( 
.A(n_3262),
.B(n_2969),
.Y(n_3573)
);

AND2x4_ASAP7_75t_L g3574 ( 
.A(n_3357),
.B(n_2955),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_R g3575 ( 
.A(n_3264),
.B(n_851),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3427),
.B(n_3018),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3292),
.B(n_3018),
.Y(n_3577)
);

AND2x4_ASAP7_75t_L g3578 ( 
.A(n_3293),
.B(n_3018),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_R g3579 ( 
.A(n_3265),
.B(n_852),
.Y(n_3579)
);

BUFx6f_ASAP7_75t_L g3580 ( 
.A(n_3294),
.Y(n_3580)
);

XNOR2xp5_ASAP7_75t_L g3581 ( 
.A(n_3191),
.B(n_2843),
.Y(n_3581)
);

XNOR2xp5_ASAP7_75t_L g3582 ( 
.A(n_3328),
.B(n_2845),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3234),
.Y(n_3583)
);

NAND2xp33_ASAP7_75t_R g3584 ( 
.A(n_3305),
.B(n_3003),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_R g3585 ( 
.A(n_3446),
.B(n_853),
.Y(n_3585)
);

CKINVDCx11_ASAP7_75t_R g3586 ( 
.A(n_3441),
.Y(n_3586)
);

AND2x4_ASAP7_75t_L g3587 ( 
.A(n_3295),
.B(n_3067),
.Y(n_3587)
);

INVxp67_ASAP7_75t_L g3588 ( 
.A(n_3403),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3402),
.B(n_2863),
.Y(n_3589)
);

OR2x6_ASAP7_75t_L g3590 ( 
.A(n_3219),
.B(n_3094),
.Y(n_3590)
);

XNOR2xp5_ASAP7_75t_L g3591 ( 
.A(n_3377),
.B(n_3252),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_R g3592 ( 
.A(n_3450),
.B(n_853),
.Y(n_3592)
);

NAND2xp33_ASAP7_75t_R g3593 ( 
.A(n_3219),
.B(n_854),
.Y(n_3593)
);

INVxp67_ASAP7_75t_L g3594 ( 
.A(n_3166),
.Y(n_3594)
);

NAND2xp33_ASAP7_75t_R g3595 ( 
.A(n_3283),
.B(n_854),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3325),
.Y(n_3596)
);

AND2x4_ASAP7_75t_L g3597 ( 
.A(n_3324),
.B(n_3067),
.Y(n_3597)
);

NOR2xp33_ASAP7_75t_R g3598 ( 
.A(n_3268),
.B(n_855),
.Y(n_3598)
);

CKINVDCx20_ASAP7_75t_R g3599 ( 
.A(n_3441),
.Y(n_3599)
);

NOR2xp33_ASAP7_75t_R g3600 ( 
.A(n_3268),
.B(n_855),
.Y(n_3600)
);

BUFx24_ASAP7_75t_SL g3601 ( 
.A(n_3272),
.Y(n_3601)
);

NAND2xp33_ASAP7_75t_R g3602 ( 
.A(n_3199),
.B(n_3434),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3173),
.B(n_2863),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3240),
.Y(n_3604)
);

CKINVDCx5p33_ASAP7_75t_R g3605 ( 
.A(n_3179),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_R g3606 ( 
.A(n_3275),
.B(n_856),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3307),
.Y(n_3607)
);

BUFx3_ASAP7_75t_L g3608 ( 
.A(n_3361),
.Y(n_3608)
);

AND2x4_ASAP7_75t_L g3609 ( 
.A(n_3330),
.B(n_3345),
.Y(n_3609)
);

INVxp67_ASAP7_75t_L g3610 ( 
.A(n_3185),
.Y(n_3610)
);

NAND2xp33_ASAP7_75t_R g3611 ( 
.A(n_3199),
.B(n_856),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3263),
.B(n_2863),
.Y(n_3612)
);

OR2x6_ASAP7_75t_L g3613 ( 
.A(n_3273),
.B(n_3077),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3307),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3201),
.B(n_3063),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3308),
.Y(n_3616)
);

NAND2xp33_ASAP7_75t_R g3617 ( 
.A(n_3434),
.B(n_857),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3427),
.B(n_3074),
.Y(n_3618)
);

NAND2xp33_ASAP7_75t_R g3619 ( 
.A(n_3366),
.B(n_857),
.Y(n_3619)
);

NAND2xp33_ASAP7_75t_R g3620 ( 
.A(n_3448),
.B(n_858),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_R g3621 ( 
.A(n_3330),
.B(n_858),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3237),
.B(n_3062),
.Y(n_3622)
);

INVx1_ASAP7_75t_SL g3623 ( 
.A(n_3193),
.Y(n_3623)
);

INVxp67_ASAP7_75t_L g3624 ( 
.A(n_3331),
.Y(n_3624)
);

NAND2xp33_ASAP7_75t_R g3625 ( 
.A(n_3448),
.B(n_859),
.Y(n_3625)
);

HB1xp67_ASAP7_75t_L g3626 ( 
.A(n_3410),
.Y(n_3626)
);

XNOR2xp5_ASAP7_75t_L g3627 ( 
.A(n_3194),
.B(n_3063),
.Y(n_3627)
);

BUFx24_ASAP7_75t_SL g3628 ( 
.A(n_3372),
.Y(n_3628)
);

AND2x4_ASAP7_75t_L g3629 ( 
.A(n_3345),
.B(n_3074),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3267),
.B(n_2935),
.Y(n_3630)
);

NAND2xp33_ASAP7_75t_R g3631 ( 
.A(n_3436),
.B(n_859),
.Y(n_3631)
);

OR2x6_ASAP7_75t_L g3632 ( 
.A(n_3352),
.B(n_3087),
.Y(n_3632)
);

BUFx3_ASAP7_75t_L g3633 ( 
.A(n_3323),
.Y(n_3633)
);

AND2x4_ASAP7_75t_L g3634 ( 
.A(n_3250),
.B(n_2917),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3204),
.B(n_2807),
.Y(n_3635)
);

XNOR2xp5_ASAP7_75t_L g3636 ( 
.A(n_3380),
.B(n_2971),
.Y(n_3636)
);

XOR2xp5_ASAP7_75t_L g3637 ( 
.A(n_3156),
.B(n_2914),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_3250),
.B(n_3087),
.Y(n_3638)
);

NAND2xp33_ASAP7_75t_R g3639 ( 
.A(n_3344),
.B(n_861),
.Y(n_3639)
);

BUFx10_ASAP7_75t_L g3640 ( 
.A(n_3364),
.Y(n_3640)
);

INVxp67_ASAP7_75t_L g3641 ( 
.A(n_3306),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_SL g3642 ( 
.A(n_3209),
.B(n_3000),
.Y(n_3642)
);

NOR2xp33_ASAP7_75t_R g3643 ( 
.A(n_3418),
.B(n_3430),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3247),
.Y(n_3644)
);

CKINVDCx5p33_ASAP7_75t_R g3645 ( 
.A(n_3379),
.Y(n_3645)
);

NAND2xp33_ASAP7_75t_R g3646 ( 
.A(n_3291),
.B(n_862),
.Y(n_3646)
);

OR2x4_ASAP7_75t_L g3647 ( 
.A(n_3266),
.B(n_3126),
.Y(n_3647)
);

AND2x4_ASAP7_75t_L g3648 ( 
.A(n_3420),
.B(n_2807),
.Y(n_3648)
);

INVxp67_ASAP7_75t_L g3649 ( 
.A(n_3437),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3308),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_R g3651 ( 
.A(n_3418),
.B(n_863),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_R g3652 ( 
.A(n_3430),
.B(n_3435),
.Y(n_3652)
);

AND2x4_ASAP7_75t_L g3653 ( 
.A(n_3435),
.B(n_2814),
.Y(n_3653)
);

INVxp67_ASAP7_75t_L g3654 ( 
.A(n_3440),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3248),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3207),
.B(n_2814),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3150),
.B(n_3110),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_R g3658 ( 
.A(n_3378),
.B(n_863),
.Y(n_3658)
);

NAND2xp33_ASAP7_75t_SL g3659 ( 
.A(n_3439),
.B(n_2969),
.Y(n_3659)
);

OR2x6_ASAP7_75t_L g3660 ( 
.A(n_3243),
.B(n_2910),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3195),
.B(n_3005),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3310),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3428),
.B(n_2935),
.Y(n_3663)
);

BUFx10_ASAP7_75t_L g3664 ( 
.A(n_3364),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3310),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3311),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3442),
.B(n_2935),
.Y(n_3667)
);

INVxp67_ASAP7_75t_L g3668 ( 
.A(n_3386),
.Y(n_3668)
);

AND2x4_ASAP7_75t_L g3669 ( 
.A(n_3209),
.B(n_2789),
.Y(n_3669)
);

OR2x6_ASAP7_75t_L g3670 ( 
.A(n_3371),
.B(n_2851),
.Y(n_3670)
);

INVxp67_ASAP7_75t_L g3671 ( 
.A(n_3387),
.Y(n_3671)
);

AND2x4_ASAP7_75t_L g3672 ( 
.A(n_3404),
.B(n_3135),
.Y(n_3672)
);

BUFx12f_ASAP7_75t_L g3673 ( 
.A(n_3349),
.Y(n_3673)
);

NAND2xp33_ASAP7_75t_R g3674 ( 
.A(n_3291),
.B(n_865),
.Y(n_3674)
);

AND2x4_ASAP7_75t_L g3675 ( 
.A(n_3429),
.B(n_3135),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_3406),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3249),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3311),
.Y(n_3678)
);

OR2x6_ASAP7_75t_L g3679 ( 
.A(n_3332),
.B(n_2941),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3312),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_3346),
.B(n_3079),
.Y(n_3681)
);

NAND2xp33_ASAP7_75t_R g3682 ( 
.A(n_3423),
.B(n_865),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3405),
.B(n_2801),
.Y(n_3683)
);

NAND2xp33_ASAP7_75t_R g3684 ( 
.A(n_3350),
.B(n_866),
.Y(n_3684)
);

OR2x4_ASAP7_75t_L g3685 ( 
.A(n_3289),
.B(n_3126),
.Y(n_3685)
);

OR2x6_ASAP7_75t_L g3686 ( 
.A(n_3251),
.B(n_2889),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_R g3687 ( 
.A(n_3378),
.B(n_869),
.Y(n_3687)
);

AND2x4_ASAP7_75t_L g3688 ( 
.A(n_3424),
.B(n_2803),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3421),
.B(n_3005),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3253),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3444),
.B(n_3449),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_R g3692 ( 
.A(n_3389),
.B(n_870),
.Y(n_3692)
);

INVxp67_ASAP7_75t_L g3693 ( 
.A(n_3431),
.Y(n_3693)
);

XOR2xp5_ASAP7_75t_L g3694 ( 
.A(n_3223),
.B(n_2879),
.Y(n_3694)
);

AND2x4_ASAP7_75t_L g3695 ( 
.A(n_3358),
.B(n_3381),
.Y(n_3695)
);

AND2x4_ASAP7_75t_L g3696 ( 
.A(n_3390),
.B(n_2804),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_R g3697 ( 
.A(n_3389),
.B(n_870),
.Y(n_3697)
);

INVx3_ASAP7_75t_L g3698 ( 
.A(n_3251),
.Y(n_3698)
);

INVxp67_ASAP7_75t_L g3699 ( 
.A(n_3321),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_R g3700 ( 
.A(n_3333),
.B(n_871),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_R g3701 ( 
.A(n_3231),
.B(n_871),
.Y(n_3701)
);

AND2x4_ASAP7_75t_L g3702 ( 
.A(n_3433),
.B(n_2806),
.Y(n_3702)
);

NAND2xp33_ASAP7_75t_R g3703 ( 
.A(n_3290),
.B(n_872),
.Y(n_3703)
);

NAND2xp33_ASAP7_75t_R g3704 ( 
.A(n_3341),
.B(n_872),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_L g3705 ( 
.A(n_3246),
.B(n_3088),
.Y(n_3705)
);

CKINVDCx11_ASAP7_75t_R g3706 ( 
.A(n_3302),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3210),
.B(n_3214),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_R g3708 ( 
.A(n_3302),
.B(n_873),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3312),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3220),
.B(n_3044),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3222),
.B(n_3044),
.Y(n_3711)
);

NOR2xp33_ASAP7_75t_R g3712 ( 
.A(n_3302),
.B(n_874),
.Y(n_3712)
);

NAND2xp33_ASAP7_75t_R g3713 ( 
.A(n_3341),
.B(n_874),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3255),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3227),
.B(n_2833),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_SL g3716 ( 
.A(n_3338),
.B(n_2959),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_SL g3717 ( 
.A(n_3286),
.B(n_3422),
.Y(n_3717)
);

AND2x4_ASAP7_75t_L g3718 ( 
.A(n_3368),
.B(n_2821),
.Y(n_3718)
);

AND2x4_ASAP7_75t_L g3719 ( 
.A(n_3375),
.B(n_2821),
.Y(n_3719)
);

INVxp67_ASAP7_75t_L g3720 ( 
.A(n_3296),
.Y(n_3720)
);

AND2x4_ASAP7_75t_L g3721 ( 
.A(n_3385),
.B(n_3229),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3233),
.B(n_2782),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3235),
.B(n_2960),
.Y(n_3723)
);

AND2x4_ASAP7_75t_L g3724 ( 
.A(n_3365),
.B(n_3367),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_3374),
.B(n_2782),
.Y(n_3725)
);

OR2x4_ASAP7_75t_L g3726 ( 
.A(n_3438),
.B(n_2983),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_R g3727 ( 
.A(n_3373),
.B(n_875),
.Y(n_3727)
);

OR2x6_ASAP7_75t_L g3728 ( 
.A(n_3452),
.B(n_2898),
.Y(n_3728)
);

INVxp67_ASAP7_75t_L g3729 ( 
.A(n_3432),
.Y(n_3729)
);

OAI22xp5_ASAP7_75t_L g3730 ( 
.A1(n_3590),
.A2(n_3451),
.B1(n_3319),
.B2(n_2915),
.Y(n_3730)
);

INVx3_ASAP7_75t_L g3731 ( 
.A(n_3464),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3556),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3504),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3571),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3538),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3607),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3614),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3616),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3630),
.B(n_3316),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3650),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3662),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3496),
.B(n_3316),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3544),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_SL g3744 ( 
.A1(n_3469),
.A2(n_3369),
.B1(n_3359),
.B2(n_3443),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3583),
.Y(n_3745)
);

BUFx2_ASAP7_75t_L g3746 ( 
.A(n_3464),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3456),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3604),
.Y(n_3748)
);

AND2x4_ASAP7_75t_L g3749 ( 
.A(n_3724),
.B(n_3164),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3482),
.B(n_3408),
.Y(n_3750)
);

OR2x2_ASAP7_75t_L g3751 ( 
.A(n_3626),
.B(n_3408),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3509),
.B(n_3409),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3691),
.B(n_3409),
.Y(n_3753)
);

OR2x2_ASAP7_75t_L g3754 ( 
.A(n_3511),
.B(n_3412),
.Y(n_3754)
);

NOR2x1_ASAP7_75t_L g3755 ( 
.A(n_3470),
.B(n_3398),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3564),
.B(n_3412),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3505),
.B(n_3413),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3514),
.B(n_3489),
.Y(n_3758)
);

BUFx3_ASAP7_75t_L g3759 ( 
.A(n_3508),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_3534),
.B(n_3422),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_3580),
.B(n_3353),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_3517),
.B(n_3413),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3462),
.B(n_3414),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3644),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3455),
.B(n_3414),
.Y(n_3765)
);

BUFx3_ASAP7_75t_L g3766 ( 
.A(n_3491),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3550),
.Y(n_3767)
);

OR2x2_ASAP7_75t_L g3768 ( 
.A(n_3535),
.B(n_3314),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3524),
.Y(n_3769)
);

OR2x2_ASAP7_75t_L g3770 ( 
.A(n_3649),
.B(n_3314),
.Y(n_3770)
);

AND2x4_ASAP7_75t_L g3771 ( 
.A(n_3653),
.B(n_3698),
.Y(n_3771)
);

INVx2_ASAP7_75t_SL g3772 ( 
.A(n_3512),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3655),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3529),
.Y(n_3774)
);

INVxp67_ASAP7_75t_SL g3775 ( 
.A(n_3526),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3603),
.B(n_3315),
.Y(n_3776)
);

OR2x2_ASAP7_75t_L g3777 ( 
.A(n_3654),
.B(n_3315),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3623),
.B(n_3370),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3677),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3539),
.Y(n_3780)
);

NOR2xp33_ASAP7_75t_L g3781 ( 
.A(n_3580),
.B(n_3445),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3485),
.B(n_3370),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_3471),
.B(n_3426),
.Y(n_3783)
);

INVxp67_ASAP7_75t_SL g3784 ( 
.A(n_3500),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3725),
.B(n_3382),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3690),
.Y(n_3786)
);

AND2x4_ASAP7_75t_L g3787 ( 
.A(n_3648),
.B(n_3164),
.Y(n_3787)
);

INVx2_ASAP7_75t_SL g3788 ( 
.A(n_3596),
.Y(n_3788)
);

INVxp67_ASAP7_75t_L g3789 ( 
.A(n_3520),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3714),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3541),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3490),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3707),
.B(n_3588),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3612),
.B(n_3165),
.Y(n_3794)
);

NOR2x1_ASAP7_75t_L g3795 ( 
.A(n_3470),
.B(n_3447),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3665),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3510),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3513),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3495),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3641),
.B(n_3384),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3492),
.B(n_3392),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3594),
.B(n_3393),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3666),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3530),
.B(n_3165),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3474),
.Y(n_3805)
);

INVx3_ASAP7_75t_L g3806 ( 
.A(n_3525),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3678),
.Y(n_3807)
);

HB1xp67_ASAP7_75t_L g3808 ( 
.A(n_3633),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3475),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3610),
.B(n_3394),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3536),
.B(n_3170),
.Y(n_3811)
);

INVx1_ASAP7_75t_SL g3812 ( 
.A(n_3596),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3680),
.Y(n_3813)
);

HB1xp67_ASAP7_75t_L g3814 ( 
.A(n_3481),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3590),
.A2(n_3069),
.B1(n_3245),
.B2(n_3161),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3709),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3668),
.B(n_3395),
.Y(n_3817)
);

INVx2_ASAP7_75t_SL g3818 ( 
.A(n_3527),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3694),
.A2(n_3060),
.B1(n_3131),
.B2(n_3119),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3459),
.Y(n_3820)
);

AND2x4_ASAP7_75t_L g3821 ( 
.A(n_3722),
.B(n_3669),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3671),
.B(n_3416),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3547),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3693),
.B(n_3170),
.Y(n_3824)
);

AND2x4_ASAP7_75t_SL g3825 ( 
.A(n_3502),
.B(n_3426),
.Y(n_3825)
);

CKINVDCx14_ASAP7_75t_R g3826 ( 
.A(n_3519),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3484),
.B(n_3171),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3721),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3695),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3552),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3663),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3577),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3503),
.Y(n_3833)
);

OR2x2_ASAP7_75t_L g3834 ( 
.A(n_3656),
.B(n_3171),
.Y(n_3834)
);

BUFx2_ASAP7_75t_L g3835 ( 
.A(n_3643),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3569),
.B(n_3172),
.Y(n_3836)
);

AND2x4_ASAP7_75t_L g3837 ( 
.A(n_3507),
.B(n_3172),
.Y(n_3837)
);

OR2x2_ASAP7_75t_L g3838 ( 
.A(n_3551),
.B(n_3174),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3635),
.Y(n_3839)
);

AND2x2_ASAP7_75t_L g3840 ( 
.A(n_3609),
.B(n_3174),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3710),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3574),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3521),
.B(n_3178),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3718),
.B(n_3178),
.Y(n_3844)
);

OR2x2_ASAP7_75t_L g3845 ( 
.A(n_3543),
.B(n_3181),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3608),
.Y(n_3846)
);

INVx2_ASAP7_75t_SL g3847 ( 
.A(n_3566),
.Y(n_3847)
);

AND2x4_ASAP7_75t_L g3848 ( 
.A(n_3719),
.B(n_3181),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3729),
.B(n_3182),
.Y(n_3849)
);

INVx2_ASAP7_75t_SL g3850 ( 
.A(n_3565),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3661),
.B(n_3182),
.Y(n_3851)
);

AND2x4_ASAP7_75t_L g3852 ( 
.A(n_3634),
.B(n_3183),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3553),
.B(n_3183),
.Y(n_3853)
);

HB1xp67_ASAP7_75t_L g3854 ( 
.A(n_3558),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3624),
.B(n_3188),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3711),
.Y(n_3856)
);

HB1xp67_ASAP7_75t_L g3857 ( 
.A(n_3602),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3667),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3589),
.B(n_3188),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3615),
.B(n_3190),
.Y(n_3860)
);

OR2x2_ASAP7_75t_SL g3861 ( 
.A(n_3523),
.B(n_3359),
.Y(n_3861)
);

OR2x2_ASAP7_75t_L g3862 ( 
.A(n_3689),
.B(n_3190),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3793),
.B(n_3537),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3829),
.B(n_3533),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3814),
.B(n_3696),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3792),
.Y(n_3866)
);

AOI31xp33_ASAP7_75t_L g3867 ( 
.A1(n_3854),
.A2(n_3857),
.A3(n_3755),
.B(n_3593),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3767),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3828),
.B(n_3717),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3797),
.Y(n_3870)
);

INVxp67_ASAP7_75t_SL g3871 ( 
.A(n_3846),
.Y(n_3871)
);

OAI221xp5_ASAP7_75t_SL g3872 ( 
.A1(n_3815),
.A2(n_3582),
.B1(n_3627),
.B2(n_3637),
.C(n_3699),
.Y(n_3872)
);

BUFx6f_ASAP7_75t_L g3873 ( 
.A(n_3759),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3798),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3750),
.B(n_3672),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3778),
.B(n_3675),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3821),
.B(n_3652),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3747),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3733),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3751),
.Y(n_3880)
);

AND2x4_ASAP7_75t_SL g3881 ( 
.A(n_3808),
.B(n_3531),
.Y(n_3881)
);

BUFx2_ASAP7_75t_L g3882 ( 
.A(n_3835),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3752),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3821),
.B(n_3756),
.Y(n_3884)
);

BUFx3_ASAP7_75t_L g3885 ( 
.A(n_3766),
.Y(n_3885)
);

OAI221xp5_ASAP7_75t_L g3886 ( 
.A1(n_3760),
.A2(n_3625),
.B1(n_3620),
.B2(n_3617),
.C(n_3611),
.Y(n_3886)
);

AOI221xp5_ASAP7_75t_L g3887 ( 
.A1(n_3823),
.A2(n_3830),
.B1(n_3705),
.B2(n_3820),
.C(n_3746),
.Y(n_3887)
);

OAI222xp33_ASAP7_75t_L g3888 ( 
.A1(n_3783),
.A2(n_3731),
.B1(n_3795),
.B2(n_3845),
.C1(n_3806),
.C2(n_3546),
.Y(n_3888)
);

OAI221xp5_ASAP7_75t_L g3889 ( 
.A1(n_3819),
.A2(n_3619),
.B1(n_3595),
.B2(n_3631),
.C(n_3684),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3754),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3757),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3840),
.B(n_3673),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3763),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3753),
.B(n_3683),
.Y(n_3894)
);

BUFx3_ASAP7_75t_L g3895 ( 
.A(n_3818),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3735),
.Y(n_3896)
);

INVx3_ASAP7_75t_L g3897 ( 
.A(n_3731),
.Y(n_3897)
);

OAI22xp5_ASAP7_75t_L g3898 ( 
.A1(n_3861),
.A2(n_3685),
.B1(n_3647),
.B2(n_3525),
.Y(n_3898)
);

INVxp67_ASAP7_75t_L g3899 ( 
.A(n_3847),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_R g3900 ( 
.A(n_3826),
.B(n_3515),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3782),
.B(n_3144),
.Y(n_3901)
);

BUFx3_ASAP7_75t_L g3902 ( 
.A(n_3850),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3743),
.Y(n_3903)
);

OAI33xp33_ASAP7_75t_L g3904 ( 
.A1(n_3838),
.A2(n_3460),
.A3(n_3720),
.B1(n_3723),
.B2(n_3716),
.B3(n_3657),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3817),
.B(n_3688),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3745),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3837),
.Y(n_3907)
);

OR2x2_ASAP7_75t_L g3908 ( 
.A(n_3762),
.B(n_3144),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3748),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3822),
.B(n_3802),
.Y(n_3910)
);

AOI21xp33_ASAP7_75t_SL g3911 ( 
.A1(n_3772),
.A2(n_3458),
.B(n_3463),
.Y(n_3911)
);

INVx2_ASAP7_75t_SL g3912 ( 
.A(n_3788),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3768),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3805),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3730),
.A2(n_3679),
.B1(n_3670),
.B2(n_3686),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3841),
.B(n_3383),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_SL g3917 ( 
.A1(n_3806),
.A2(n_3581),
.B(n_3461),
.Y(n_3917)
);

BUFx3_ASAP7_75t_L g3918 ( 
.A(n_3812),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3841),
.B(n_3388),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3856),
.B(n_3397),
.Y(n_3920)
);

BUFx3_ASAP7_75t_L g3921 ( 
.A(n_3825),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3809),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3810),
.B(n_3702),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3770),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3764),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3777),
.Y(n_3926)
);

OR2x2_ASAP7_75t_L g3927 ( 
.A(n_3831),
.B(n_3148),
.Y(n_3927)
);

OAI221xp5_ASAP7_75t_L g3928 ( 
.A1(n_3744),
.A2(n_3703),
.B1(n_3682),
.B2(n_3506),
.C(n_3639),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3773),
.Y(n_3929)
);

AOI222xp33_ASAP7_75t_L g3930 ( 
.A1(n_3789),
.A2(n_3586),
.B1(n_3498),
.B2(n_3601),
.C1(n_3479),
.C2(n_3622),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3799),
.Y(n_3931)
);

OR2x2_ASAP7_75t_L g3932 ( 
.A(n_3862),
.B(n_3148),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3749),
.A2(n_3679),
.B1(n_3670),
.B2(n_3686),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3758),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3779),
.Y(n_3935)
);

AOI221xp5_ASAP7_75t_SL g3936 ( 
.A1(n_3784),
.A2(n_3599),
.B1(n_3591),
.B2(n_3501),
.C(n_3636),
.Y(n_3936)
);

BUFx2_ASAP7_75t_L g3937 ( 
.A(n_3775),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3855),
.Y(n_3938)
);

HB1xp67_ASAP7_75t_L g3939 ( 
.A(n_3837),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3785),
.B(n_3645),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3800),
.B(n_3676),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3732),
.Y(n_3942)
);

HB1xp67_ASAP7_75t_L g3943 ( 
.A(n_3786),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3790),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3849),
.B(n_3557),
.Y(n_3945)
);

AND2x4_ASAP7_75t_L g3946 ( 
.A(n_3852),
.B(n_3149),
.Y(n_3946)
);

HB1xp67_ASAP7_75t_L g3947 ( 
.A(n_3765),
.Y(n_3947)
);

AND2x2_ASAP7_75t_L g3948 ( 
.A(n_3832),
.B(n_3476),
.Y(n_3948)
);

INVx4_ASAP7_75t_L g3949 ( 
.A(n_3749),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3732),
.Y(n_3950)
);

BUFx3_ASAP7_75t_L g3951 ( 
.A(n_3781),
.Y(n_3951)
);

HB1xp67_ASAP7_75t_L g3952 ( 
.A(n_3801),
.Y(n_3952)
);

AND2x4_ASAP7_75t_L g3953 ( 
.A(n_3852),
.B(n_3149),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3824),
.B(n_3629),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3734),
.Y(n_3955)
);

OR2x2_ASAP7_75t_L g3956 ( 
.A(n_3843),
.B(n_3153),
.Y(n_3956)
);

HB1xp67_ASAP7_75t_L g3957 ( 
.A(n_3827),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3853),
.B(n_3632),
.Y(n_3958)
);

INVx1_ASAP7_75t_SL g3959 ( 
.A(n_3771),
.Y(n_3959)
);

OAI222xp33_ASAP7_75t_L g3960 ( 
.A1(n_3860),
.A2(n_3632),
.B1(n_3660),
.B2(n_3613),
.C1(n_3563),
.C2(n_3642),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3959),
.B(n_3771),
.Y(n_3961)
);

AND3x2_ASAP7_75t_L g3962 ( 
.A(n_3882),
.B(n_3761),
.C(n_3540),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3959),
.B(n_3836),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3949),
.B(n_3842),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3901),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3943),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3952),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3957),
.B(n_3856),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3949),
.B(n_3742),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3865),
.B(n_3858),
.Y(n_3970)
);

OR2x2_ASAP7_75t_L g3971 ( 
.A(n_3880),
.B(n_3839),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3950),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3876),
.B(n_3844),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3897),
.B(n_3844),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3908),
.B(n_3839),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3884),
.B(n_3848),
.Y(n_3976)
);

INVx1_ASAP7_75t_SL g3977 ( 
.A(n_3873),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3907),
.B(n_3848),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3887),
.B(n_3833),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3939),
.B(n_3787),
.Y(n_3980)
);

OR2x2_ASAP7_75t_L g3981 ( 
.A(n_3913),
.B(n_3776),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3914),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3887),
.B(n_3833),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3922),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3937),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3866),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3924),
.B(n_3739),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3905),
.B(n_3787),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3870),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3897),
.B(n_3834),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3926),
.B(n_3794),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3923),
.B(n_3859),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3931),
.Y(n_3993)
);

NOR2xp33_ASAP7_75t_L g3994 ( 
.A(n_3917),
.B(n_3726),
.Y(n_3994)
);

OR2x2_ASAP7_75t_L g3995 ( 
.A(n_3893),
.B(n_3934),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3942),
.Y(n_3996)
);

INVxp67_ASAP7_75t_SL g3997 ( 
.A(n_3871),
.Y(n_3997)
);

OR2x2_ASAP7_75t_L g3998 ( 
.A(n_3932),
.B(n_3891),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3910),
.B(n_3851),
.Y(n_3999)
);

NOR2xp33_ASAP7_75t_L g4000 ( 
.A(n_3917),
.B(n_3605),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3955),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3894),
.B(n_3816),
.Y(n_4002)
);

OR2x2_ASAP7_75t_L g4003 ( 
.A(n_3883),
.B(n_3804),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3874),
.Y(n_4004)
);

OR2x2_ASAP7_75t_L g4005 ( 
.A(n_3890),
.B(n_3811),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3938),
.B(n_3769),
.Y(n_4006)
);

OR2x2_ASAP7_75t_L g4007 ( 
.A(n_3947),
.B(n_3774),
.Y(n_4007)
);

OR2x2_ASAP7_75t_L g4008 ( 
.A(n_3956),
.B(n_3780),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3945),
.B(n_3813),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3879),
.B(n_3791),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3875),
.B(n_3807),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_3873),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3896),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3868),
.B(n_3878),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3903),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3906),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3954),
.B(n_3803),
.Y(n_4017)
);

AND2x2_ASAP7_75t_L g4018 ( 
.A(n_3877),
.B(n_3734),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3916),
.B(n_3736),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3958),
.B(n_3948),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3909),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3925),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3929),
.Y(n_4023)
);

OR2x2_ASAP7_75t_L g4024 ( 
.A(n_3927),
.B(n_3736),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_3864),
.B(n_3737),
.Y(n_4025)
);

AND2x4_ASAP7_75t_SL g4026 ( 
.A(n_3873),
.B(n_3640),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3935),
.Y(n_4027)
);

BUFx2_ASAP7_75t_SL g4028 ( 
.A(n_3885),
.Y(n_4028)
);

INVxp67_ASAP7_75t_L g4029 ( 
.A(n_3918),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3863),
.B(n_3737),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3944),
.Y(n_4031)
);

OR2x2_ASAP7_75t_L g4032 ( 
.A(n_3916),
.B(n_3738),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_3869),
.B(n_3738),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3912),
.B(n_3740),
.Y(n_4034)
);

OR2x2_ASAP7_75t_L g4035 ( 
.A(n_3919),
.B(n_3740),
.Y(n_4035)
);

BUFx3_ASAP7_75t_L g4036 ( 
.A(n_3881),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3946),
.Y(n_4037)
);

NOR2xp33_ASAP7_75t_L g4038 ( 
.A(n_3889),
.B(n_3872),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3940),
.B(n_3741),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3919),
.Y(n_4040)
);

NAND2xp33_ASAP7_75t_SL g4041 ( 
.A(n_3969),
.B(n_3900),
.Y(n_4041)
);

AOI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_4038),
.A2(n_3928),
.B1(n_3915),
.B2(n_3936),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3979),
.B(n_3867),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_4036),
.B(n_3921),
.Y(n_4044)
);

NAND2xp33_ASAP7_75t_R g4045 ( 
.A(n_3962),
.B(n_3911),
.Y(n_4045)
);

AO221x2_ASAP7_75t_L g4046 ( 
.A1(n_4028),
.A2(n_3888),
.B1(n_3898),
.B2(n_3960),
.C(n_3867),
.Y(n_4046)
);

NOR2x1_ASAP7_75t_L g4047 ( 
.A(n_4012),
.B(n_3886),
.Y(n_4047)
);

NAND2xp33_ASAP7_75t_SL g4048 ( 
.A(n_3961),
.B(n_3898),
.Y(n_4048)
);

INVx4_ASAP7_75t_L g4049 ( 
.A(n_4026),
.Y(n_4049)
);

OAI22xp33_ASAP7_75t_L g4050 ( 
.A1(n_3997),
.A2(n_3928),
.B1(n_3886),
.B2(n_3911),
.Y(n_4050)
);

AOI22xp5_ASAP7_75t_L g4051 ( 
.A1(n_3994),
.A2(n_3936),
.B1(n_3889),
.B2(n_3930),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3983),
.B(n_3946),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_4040),
.B(n_3953),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_4040),
.B(n_3953),
.Y(n_4054)
);

AND2x4_ASAP7_75t_L g4055 ( 
.A(n_4029),
.B(n_3895),
.Y(n_4055)
);

AND2x4_ASAP7_75t_SL g4056 ( 
.A(n_3964),
.B(n_3941),
.Y(n_4056)
);

CKINVDCx5p33_ASAP7_75t_R g4057 ( 
.A(n_3977),
.Y(n_4057)
);

AO221x2_ASAP7_75t_L g4058 ( 
.A1(n_4000),
.A2(n_3888),
.B1(n_3960),
.B2(n_3967),
.C(n_3985),
.Y(n_4058)
);

OAI221xp5_ASAP7_75t_L g4059 ( 
.A1(n_3968),
.A2(n_3872),
.B1(n_3933),
.B2(n_3930),
.C(n_3522),
.Y(n_4059)
);

AO221x2_ASAP7_75t_L g4060 ( 
.A1(n_4037),
.A2(n_3542),
.B1(n_3902),
.B2(n_3904),
.C(n_3899),
.Y(n_4060)
);

INVxp67_ASAP7_75t_L g4061 ( 
.A(n_4014),
.Y(n_4061)
);

NOR2xp33_ASAP7_75t_L g4062 ( 
.A(n_4018),
.B(n_3951),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_4032),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3965),
.B(n_3920),
.Y(n_4064)
);

OAI22xp5_ASAP7_75t_SL g4065 ( 
.A1(n_3974),
.A2(n_3453),
.B1(n_3454),
.B2(n_3613),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3965),
.B(n_3920),
.Y(n_4066)
);

NAND2xp33_ASAP7_75t_SL g4067 ( 
.A(n_3980),
.B(n_3560),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3999),
.B(n_3741),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3990),
.A2(n_3904),
.B1(n_3555),
.B2(n_3567),
.Y(n_4069)
);

NOR2x1_ASAP7_75t_L g4070 ( 
.A(n_3974),
.B(n_3478),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_4033),
.B(n_3796),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_4030),
.B(n_3796),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_4039),
.Y(n_4073)
);

NOR2x1_ASAP7_75t_L g4074 ( 
.A(n_3966),
.B(n_3576),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_3975),
.B(n_3327),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4035),
.Y(n_4076)
);

NOR2xp33_ASAP7_75t_L g4077 ( 
.A(n_4006),
.B(n_3892),
.Y(n_4077)
);

NOR2xp33_ASAP7_75t_L g4078 ( 
.A(n_4020),
.B(n_3618),
.Y(n_4078)
);

OAI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3998),
.A2(n_3554),
.B1(n_3545),
.B2(n_3549),
.Y(n_4079)
);

AOI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3990),
.A2(n_3497),
.B1(n_3559),
.B2(n_3681),
.Y(n_4080)
);

AO221x2_ASAP7_75t_L g4081 ( 
.A1(n_3987),
.A2(n_3516),
.B1(n_3518),
.B2(n_3575),
.C(n_3568),
.Y(n_4081)
);

AOI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_4034),
.A2(n_3473),
.B1(n_3659),
.B2(n_3573),
.Y(n_4082)
);

NOR2xp33_ASAP7_75t_L g4083 ( 
.A(n_4003),
.B(n_4005),
.Y(n_4083)
);

NAND2xp33_ASAP7_75t_SL g4084 ( 
.A(n_3978),
.B(n_3598),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3976),
.B(n_3465),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3971),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_R g4087 ( 
.A(n_3973),
.B(n_3706),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_4007),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3982),
.B(n_3347),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3984),
.B(n_3348),
.Y(n_4090)
);

OR2x2_ASAP7_75t_L g4091 ( 
.A(n_3981),
.B(n_3334),
.Y(n_4091)
);

AOI22xp5_ASAP7_75t_L g4092 ( 
.A1(n_4025),
.A2(n_3472),
.B1(n_3494),
.B2(n_3493),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_3991),
.B(n_4008),
.Y(n_4093)
);

AO221x2_ASAP7_75t_L g4094 ( 
.A1(n_3993),
.A2(n_3579),
.B1(n_3562),
.B2(n_3606),
.C(n_3600),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_4009),
.B(n_3664),
.Y(n_4095)
);

NOR2xp67_ASAP7_75t_L g4096 ( 
.A(n_4013),
.B(n_3532),
.Y(n_4096)
);

OAI22xp33_ASAP7_75t_L g4097 ( 
.A1(n_3995),
.A2(n_3528),
.B1(n_3674),
.B2(n_3646),
.Y(n_4097)
);

NOR2xp33_ASAP7_75t_L g4098 ( 
.A(n_3988),
.B(n_3660),
.Y(n_4098)
);

NAND2xp33_ASAP7_75t_SL g4099 ( 
.A(n_3963),
.B(n_3621),
.Y(n_4099)
);

AND2x4_ASAP7_75t_L g4100 ( 
.A(n_4044),
.B(n_4017),
.Y(n_4100)
);

NOR2xp33_ASAP7_75t_L g4101 ( 
.A(n_4049),
.B(n_4011),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_4046),
.B(n_3992),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_SL g4103 ( 
.A(n_4050),
.B(n_4013),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_4065),
.B(n_4024),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4046),
.B(n_3970),
.Y(n_4105)
);

CKINVDCx20_ASAP7_75t_R g4106 ( 
.A(n_4041),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_4063),
.B(n_3996),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_4093),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4076),
.B(n_3996),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_4088),
.Y(n_4110)
);

NOR2xp33_ASAP7_75t_L g4111 ( 
.A(n_4042),
.B(n_4002),
.Y(n_4111)
);

NOR2xp33_ASAP7_75t_L g4112 ( 
.A(n_4051),
.B(n_4010),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_4047),
.B(n_4001),
.Y(n_4113)
);

BUFx3_ASAP7_75t_L g4114 ( 
.A(n_4057),
.Y(n_4114)
);

INVx2_ASAP7_75t_SL g4115 ( 
.A(n_4056),
.Y(n_4115)
);

INVx1_ASAP7_75t_SL g4116 ( 
.A(n_4067),
.Y(n_4116)
);

INVx1_ASAP7_75t_SL g4117 ( 
.A(n_4055),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_4086),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4058),
.B(n_4001),
.Y(n_4119)
);

INVx1_ASAP7_75t_SL g4120 ( 
.A(n_4099),
.Y(n_4120)
);

INVx1_ASAP7_75t_SL g4121 ( 
.A(n_4084),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_4058),
.B(n_3986),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4064),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_4066),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_4096),
.B(n_3989),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_4080),
.B(n_4004),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4075),
.Y(n_4127)
);

INVx1_ASAP7_75t_SL g4128 ( 
.A(n_4087),
.Y(n_4128)
);

BUFx2_ASAP7_75t_L g4129 ( 
.A(n_4070),
.Y(n_4129)
);

INVxp67_ASAP7_75t_L g4130 ( 
.A(n_4045),
.Y(n_4130)
);

HB1xp67_ASAP7_75t_L g4131 ( 
.A(n_4061),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_4053),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_4054),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4091),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_4089),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_4043),
.B(n_4019),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_4052),
.B(n_3972),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4090),
.Y(n_4138)
);

INVx2_ASAP7_75t_L g4139 ( 
.A(n_4071),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_4083),
.B(n_3972),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_4059),
.A2(n_4060),
.B1(n_4048),
.B2(n_4094),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_4072),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4068),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_4098),
.B(n_4023),
.Y(n_4144)
);

OAI22xp5_ASAP7_75t_L g4145 ( 
.A1(n_4069),
.A2(n_3480),
.B1(n_4016),
.B2(n_4015),
.Y(n_4145)
);

INVx3_ASAP7_75t_L g4146 ( 
.A(n_4060),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4097),
.B(n_4015),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_4073),
.Y(n_4148)
);

AOI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_4081),
.A2(n_4021),
.B1(n_4022),
.B2(n_4016),
.Y(n_4149)
);

NOR2xp33_ASAP7_75t_L g4150 ( 
.A(n_4077),
.B(n_4021),
.Y(n_4150)
);

INVx3_ASAP7_75t_SL g4151 ( 
.A(n_4085),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4074),
.Y(n_4152)
);

INVx1_ASAP7_75t_SL g4153 ( 
.A(n_4062),
.Y(n_4153)
);

OR2x2_ASAP7_75t_L g4154 ( 
.A(n_4092),
.B(n_4022),
.Y(n_4154)
);

OR2x2_ASAP7_75t_L g4155 ( 
.A(n_4079),
.B(n_4031),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4078),
.B(n_4027),
.Y(n_4156)
);

BUFx3_ASAP7_75t_L g4157 ( 
.A(n_4081),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4095),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_4082),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4112),
.B(n_4027),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_4146),
.B(n_4141),
.Y(n_4161)
);

INVxp67_ASAP7_75t_SL g4162 ( 
.A(n_4114),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4108),
.Y(n_4163)
);

O2A1O1Ixp33_ASAP7_75t_L g4164 ( 
.A1(n_4130),
.A2(n_3425),
.B(n_3108),
.C(n_3090),
.Y(n_4164)
);

AOI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_4157),
.A2(n_3713),
.B1(n_3704),
.B2(n_3584),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_4128),
.B(n_4031),
.Y(n_4166)
);

AOI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_4121),
.A2(n_3572),
.B1(n_3638),
.B2(n_3570),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_4131),
.B(n_3561),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4140),
.Y(n_4169)
);

AO22x1_ASAP7_75t_L g4170 ( 
.A1(n_4121),
.A2(n_3548),
.B1(n_3466),
.B2(n_3468),
.Y(n_4170)
);

OR2x2_ASAP7_75t_L g4171 ( 
.A(n_4123),
.B(n_3335),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_4117),
.B(n_3578),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4140),
.Y(n_4173)
);

BUFx3_ASAP7_75t_L g4174 ( 
.A(n_4148),
.Y(n_4174)
);

NAND4xp25_ASAP7_75t_SL g4175 ( 
.A(n_4116),
.B(n_3457),
.C(n_3651),
.D(n_3411),
.Y(n_4175)
);

AOI22xp5_ASAP7_75t_L g4176 ( 
.A1(n_4120),
.A2(n_3728),
.B1(n_3715),
.B2(n_3355),
.Y(n_4176)
);

AND2x4_ASAP7_75t_SL g4177 ( 
.A(n_4115),
.B(n_3587),
.Y(n_4177)
);

AOI221xp5_ASAP7_75t_L g4178 ( 
.A1(n_4119),
.A2(n_3488),
.B1(n_3592),
.B2(n_3585),
.C(n_3467),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4143),
.B(n_3700),
.Y(n_4179)
);

OAI32xp33_ASAP7_75t_L g4180 ( 
.A1(n_4146),
.A2(n_3687),
.A3(n_3697),
.B1(n_3692),
.B2(n_3658),
.Y(n_4180)
);

INVx1_ASAP7_75t_SL g4181 ( 
.A(n_4128),
.Y(n_4181)
);

NAND4xp25_ASAP7_75t_L g4182 ( 
.A(n_4116),
.B(n_4120),
.C(n_4104),
.D(n_4117),
.Y(n_4182)
);

AOI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_4102),
.A2(n_4111),
.B1(n_4105),
.B2(n_4106),
.Y(n_4183)
);

OAI21xp33_ASAP7_75t_L g4184 ( 
.A1(n_4122),
.A2(n_3708),
.B(n_3701),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4107),
.Y(n_4185)
);

OR2x2_ASAP7_75t_L g4186 ( 
.A(n_4124),
.B(n_3336),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_4138),
.B(n_3354),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4136),
.B(n_4132),
.Y(n_4188)
);

OR2x2_ASAP7_75t_L g4189 ( 
.A(n_4137),
.B(n_3340),
.Y(n_4189)
);

OAI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_4153),
.A2(n_4149),
.B1(n_4151),
.B2(n_4159),
.Y(n_4190)
);

AOI22xp5_ASAP7_75t_SL g4191 ( 
.A1(n_4153),
.A2(n_3727),
.B1(n_3712),
.B2(n_3597),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_4101),
.B(n_3477),
.Y(n_4192)
);

AOI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_4103),
.A2(n_3342),
.B(n_2986),
.Y(n_4193)
);

AOI31xp33_ASAP7_75t_SL g4194 ( 
.A1(n_4147),
.A2(n_3040),
.A3(n_2839),
.B(n_2933),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4136),
.B(n_3343),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_SL g4196 ( 
.A(n_4129),
.B(n_3483),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4107),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4181),
.B(n_4135),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_4174),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4163),
.Y(n_4200)
);

AND2x4_ASAP7_75t_L g4201 ( 
.A(n_4162),
.B(n_4100),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_4169),
.B(n_4118),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4166),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4172),
.B(n_4113),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4173),
.B(n_4134),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4188),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_4183),
.B(n_4133),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4185),
.B(n_4139),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4177),
.B(n_4126),
.Y(n_4209)
);

NAND2xp33_ASAP7_75t_SL g4210 ( 
.A(n_4161),
.B(n_4155),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4187),
.Y(n_4211)
);

AOI31xp33_ASAP7_75t_L g4212 ( 
.A1(n_4178),
.A2(n_4145),
.A3(n_4158),
.B(n_4152),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4197),
.B(n_4142),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4168),
.Y(n_4214)
);

INVxp67_ASAP7_75t_L g4215 ( 
.A(n_4182),
.Y(n_4215)
);

INVx1_ASAP7_75t_SL g4216 ( 
.A(n_4191),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4192),
.B(n_4100),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_4160),
.B(n_4127),
.Y(n_4218)
);

AOI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_4190),
.A2(n_4145),
.B1(n_4154),
.B2(n_4156),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4193),
.B(n_4150),
.Y(n_4220)
);

AND2x4_ASAP7_75t_L g4221 ( 
.A(n_4196),
.B(n_4144),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4189),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4176),
.B(n_4137),
.Y(n_4223)
);

NOR2x1_ASAP7_75t_L g4224 ( 
.A(n_4175),
.B(n_4156),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_4184),
.B(n_4109),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4179),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_SL g4227 ( 
.A(n_4167),
.B(n_4110),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4199),
.B(n_4195),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_4215),
.B(n_4170),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4198),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4202),
.Y(n_4231)
);

HB1xp67_ASAP7_75t_L g4232 ( 
.A(n_4200),
.Y(n_4232)
);

INVxp33_ASAP7_75t_SL g4233 ( 
.A(n_4216),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4218),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4201),
.Y(n_4235)
);

INVxp67_ASAP7_75t_L g4236 ( 
.A(n_4201),
.Y(n_4236)
);

INVx1_ASAP7_75t_SL g4237 ( 
.A(n_4226),
.Y(n_4237)
);

BUFx12f_ASAP7_75t_L g4238 ( 
.A(n_4221),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4208),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4213),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4205),
.Y(n_4241)
);

INVxp67_ASAP7_75t_L g4242 ( 
.A(n_4203),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4206),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_4212),
.B(n_4165),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4222),
.Y(n_4245)
);

INVxp67_ASAP7_75t_L g4246 ( 
.A(n_4207),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4204),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4221),
.Y(n_4248)
);

NOR2xp33_ASAP7_75t_L g4249 ( 
.A(n_4209),
.B(n_4171),
.Y(n_4249)
);

BUFx6f_ASAP7_75t_L g4250 ( 
.A(n_4217),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4211),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4214),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4220),
.B(n_4109),
.Y(n_4253)
);

AOI211x1_ASAP7_75t_SL g4254 ( 
.A1(n_4244),
.A2(n_4223),
.B(n_4227),
.C(n_4210),
.Y(n_4254)
);

AOI211xp5_ASAP7_75t_L g4255 ( 
.A1(n_4236),
.A2(n_4180),
.B(n_4225),
.C(n_4194),
.Y(n_4255)
);

OAI211xp5_ASAP7_75t_SL g4256 ( 
.A1(n_4246),
.A2(n_4224),
.B(n_4219),
.C(n_4165),
.Y(n_4256)
);

NAND4xp25_ASAP7_75t_L g4257 ( 
.A(n_4229),
.B(n_4164),
.C(n_2904),
.D(n_2835),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_SL g4258 ( 
.A(n_4233),
.B(n_4186),
.Y(n_4258)
);

NAND4xp25_ASAP7_75t_L g4259 ( 
.A(n_4235),
.B(n_3021),
.C(n_3004),
.D(n_3123),
.Y(n_4259)
);

AOI222xp33_ASAP7_75t_L g4260 ( 
.A1(n_4230),
.A2(n_4125),
.B1(n_2926),
.B2(n_3061),
.C1(n_2817),
.C2(n_2785),
.Y(n_4260)
);

NOR3xp33_ASAP7_75t_L g4261 ( 
.A(n_4242),
.B(n_4237),
.C(n_4248),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4231),
.Y(n_4262)
);

NOR2x1_ASAP7_75t_L g4263 ( 
.A(n_4243),
.B(n_3339),
.Y(n_4263)
);

NOR3xp33_ASAP7_75t_L g4264 ( 
.A(n_4239),
.B(n_4240),
.C(n_4234),
.Y(n_4264)
);

OAI32xp33_ASAP7_75t_L g4265 ( 
.A1(n_4247),
.A2(n_4241),
.A3(n_4253),
.B1(n_4245),
.B2(n_4252),
.Y(n_4265)
);

AND3x1_ASAP7_75t_L g4266 ( 
.A(n_4249),
.B(n_2913),
.C(n_3278),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4232),
.B(n_3351),
.Y(n_4267)
);

A2O1A1Ixp33_ASAP7_75t_SL g4268 ( 
.A1(n_4251),
.A2(n_2965),
.B(n_2991),
.C(n_3028),
.Y(n_4268)
);

AOI211xp5_ASAP7_75t_SL g4269 ( 
.A1(n_4228),
.A2(n_3058),
.B(n_2882),
.C(n_3140),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_L g4270 ( 
.A(n_4238),
.B(n_875),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4250),
.B(n_876),
.Y(n_4271)
);

OAI211xp5_ASAP7_75t_L g4272 ( 
.A1(n_4255),
.A2(n_4250),
.B(n_2836),
.C(n_2878),
.Y(n_4272)
);

OAI22xp5_ASAP7_75t_L g4273 ( 
.A1(n_4270),
.A2(n_4250),
.B1(n_3728),
.B2(n_3030),
.Y(n_4273)
);

NAND3xp33_ASAP7_75t_L g4274 ( 
.A(n_4261),
.B(n_3091),
.C(n_3072),
.Y(n_4274)
);

OAI211xp5_ASAP7_75t_SL g4275 ( 
.A1(n_4254),
.A2(n_2927),
.B(n_3111),
.C(n_2964),
.Y(n_4275)
);

OAI22xp5_ASAP7_75t_L g4276 ( 
.A1(n_4262),
.A2(n_3046),
.B1(n_3317),
.B2(n_3068),
.Y(n_4276)
);

OAI22xp33_ASAP7_75t_L g4277 ( 
.A1(n_4257),
.A2(n_3057),
.B1(n_2865),
.B2(n_2871),
.Y(n_4277)
);

A2O1A1Ixp33_ASAP7_75t_SL g4278 ( 
.A1(n_4264),
.A2(n_4256),
.B(n_4271),
.C(n_4265),
.Y(n_4278)
);

AOI22xp5_ASAP7_75t_L g4279 ( 
.A1(n_4258),
.A2(n_3487),
.B1(n_3499),
.B2(n_3486),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4263),
.Y(n_4280)
);

BUFx2_ASAP7_75t_L g4281 ( 
.A(n_4267),
.Y(n_4281)
);

CKINVDCx5p33_ASAP7_75t_R g4282 ( 
.A(n_4266),
.Y(n_4282)
);

OR2x2_ASAP7_75t_L g4283 ( 
.A(n_4268),
.B(n_876),
.Y(n_4283)
);

AOI221xp5_ASAP7_75t_L g4284 ( 
.A1(n_4259),
.A2(n_3097),
.B1(n_3013),
.B2(n_3075),
.C(n_2776),
.Y(n_4284)
);

NOR2x1_ASAP7_75t_L g4285 ( 
.A(n_4283),
.B(n_3008),
.Y(n_4285)
);

OR2x2_ASAP7_75t_L g4286 ( 
.A(n_4281),
.B(n_877),
.Y(n_4286)
);

HB1xp67_ASAP7_75t_L g4287 ( 
.A(n_4280),
.Y(n_4287)
);

NAND4xp75_ASAP7_75t_L g4288 ( 
.A(n_4278),
.B(n_2887),
.C(n_4260),
.D(n_3133),
.Y(n_4288)
);

NAND2xp33_ASAP7_75t_L g4289 ( 
.A(n_4282),
.B(n_4269),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_4279),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4274),
.Y(n_4291)
);

NAND4xp75_ASAP7_75t_L g4292 ( 
.A(n_4272),
.B(n_2963),
.C(n_2942),
.D(n_2956),
.Y(n_4292)
);

NOR2xp33_ASAP7_75t_R g4293 ( 
.A(n_4289),
.B(n_877),
.Y(n_4293)
);

NOR2xp33_ASAP7_75t_R g4294 ( 
.A(n_4286),
.B(n_878),
.Y(n_4294)
);

NAND2xp33_ASAP7_75t_SL g4295 ( 
.A(n_4287),
.B(n_4273),
.Y(n_4295)
);

OAI22xp5_ASAP7_75t_SL g4296 ( 
.A1(n_4293),
.A2(n_4291),
.B1(n_4290),
.B2(n_4285),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4295),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4294),
.B(n_4288),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4297),
.Y(n_4299)
);

AOI22xp33_ASAP7_75t_L g4300 ( 
.A1(n_4299),
.A2(n_4296),
.B1(n_4298),
.B2(n_4277),
.Y(n_4300)
);

OAI22xp5_ASAP7_75t_SL g4301 ( 
.A1(n_4300),
.A2(n_4276),
.B1(n_4275),
.B2(n_4292),
.Y(n_4301)
);

OAI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4301),
.A2(n_4284),
.B(n_2932),
.Y(n_4302)
);

AOI222xp33_ASAP7_75t_SL g4303 ( 
.A1(n_4302),
.A2(n_3628),
.B1(n_2939),
.B2(n_2853),
.C1(n_3114),
.C2(n_880),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4303),
.Y(n_4304)
);

OAI221xp5_ASAP7_75t_L g4305 ( 
.A1(n_4304),
.A2(n_3134),
.B1(n_2874),
.B2(n_3139),
.C(n_3070),
.Y(n_4305)
);

AOI211xp5_ASAP7_75t_L g4306 ( 
.A1(n_4305),
.A2(n_3105),
.B(n_3106),
.C(n_3093),
.Y(n_4306)
);


endmodule