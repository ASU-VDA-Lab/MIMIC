module fake_netlist_5_340_n_1803 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1803);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1803;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_62),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_11),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_45),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_25),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_67),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_30),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_83),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_58),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_24),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_63),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_66),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_116),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_101),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_16),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_64),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_50),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_19),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_54),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_76),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_21),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_73),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_59),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_77),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_35),
.Y(n_193)
);

BUFx8_ASAP7_75t_SL g194 ( 
.A(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_85),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_107),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_44),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_115),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_48),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_20),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_78),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

BUFx2_ASAP7_75t_SL g208 ( 
.A(n_36),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_53),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_95),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_105),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_42),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_146),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_61),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_16),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_46),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_33),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_22),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_3),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_49),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_10),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_6),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_148),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_75),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_144),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_25),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_80),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_70),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_11),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_135),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_36),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_41),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_151),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_9),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_120),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_84),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_137),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_145),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_119),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_24),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_91),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_140),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_79),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_0),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_153),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_154),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_41),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_4),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_52),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_89),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_114),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_5),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_69),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_51),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_17),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_55),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_50),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_86),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_26),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_100),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_46),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_26),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_7),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_136),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_65),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_134),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_150),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_99),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_96),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_139),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_124),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_131),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_60),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_194),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_199),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_156),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_168),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_203),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_168),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_183),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_207),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_183),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_157),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_189),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_163),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_204),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_267),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_271),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_182),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_160),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_221),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_165),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_167),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_170),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_176),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_221),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_184),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_248),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_169),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_288),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_179),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_169),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_180),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_186),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_188),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_166),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_171),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_175),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_190),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_175),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_171),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_270),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_279),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_289),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_234),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_158),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_234),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_192),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_274),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_261),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_207),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_196),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_259),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_R g395 ( 
.A(n_312),
.B(n_198),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_370),
.B(n_171),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_314),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_322),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_R g401 ( 
.A(n_317),
.B(n_162),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_324),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_247),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_161),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_285),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_247),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_159),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_316),
.B(n_161),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_159),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_209),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_323),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_313),
.B(n_315),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_313),
.B(n_173),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_327),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_334),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_344),
.B(n_172),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_323),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_334),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

AND3x2_ASAP7_75t_L g435 ( 
.A(n_350),
.B(n_191),
.C(n_172),
.Y(n_435)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_191),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_325),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_325),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_319),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_315),
.B(n_173),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_326),
.B(n_174),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_336),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_337),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_386),
.B(n_303),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_334),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_386),
.B(n_303),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_174),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_326),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_385),
.B(n_329),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_328),
.B(n_332),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_328),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_332),
.B(n_185),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_335),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_338),
.B(n_185),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_335),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_339),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_340),
.B(n_212),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_421),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_449),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_400),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_427),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_408),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_417),
.B(n_331),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_427),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_402),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_417),
.A2(n_447),
.B1(n_415),
.B2(n_408),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_417),
.B(n_207),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_420),
.B(n_370),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

OAI22xp33_ASAP7_75t_L g484 ( 
.A1(n_394),
.A2(n_343),
.B1(n_377),
.B2(n_333),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_389),
.B(n_348),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_434),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_389),
.B(n_354),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_356),
.Y(n_493)
);

BUFx4f_ASAP7_75t_L g494 ( 
.A(n_430),
.Y(n_494)
);

AND3x2_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_379),
.C(n_205),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_423),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_408),
.A2(n_254),
.B1(n_208),
.B2(n_193),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_454),
.B(n_207),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_376),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_413),
.B(n_357),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_413),
.B(n_359),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_423),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_396),
.B(n_208),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_423),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_187),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_401),
.A2(n_384),
.B1(n_378),
.B2(n_377),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_430),
.B(n_187),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_429),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_421),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_401),
.A2(n_378),
.B1(n_343),
.B2(n_333),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_422),
.B(n_376),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_422),
.B(n_376),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_415),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_415),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_444),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_400),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_458),
.B(n_261),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_449),
.B(n_330),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_420),
.B(n_342),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_444),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_396),
.B(n_342),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_407),
.B(n_341),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_444),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_446),
.A2(n_452),
.B1(n_441),
.B2(n_426),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_436),
.B(n_446),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_436),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_397),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_428),
.B(n_215),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_428),
.B(n_254),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_441),
.B(n_195),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_429),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_429),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_446),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_442),
.B(n_164),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_450),
.B(n_346),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_R g555 ( 
.A(n_402),
.B(n_214),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_421),
.B(n_217),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_432),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_421),
.B(n_233),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_432),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_449),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_421),
.B(n_235),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_391),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_391),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_445),
.B(n_236),
.Y(n_570)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_390),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_393),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_441),
.B(n_195),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_445),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_426),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_442),
.B(n_178),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_445),
.B(n_452),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_445),
.B(n_238),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_443),
.B(n_215),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_443),
.B(n_215),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_445),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_435),
.Y(n_582)
);

AND3x1_ASAP7_75t_L g583 ( 
.A(n_452),
.B(n_347),
.C(n_346),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_445),
.B(n_239),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_445),
.B(n_243),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_440),
.A2(n_200),
.B1(n_201),
.B2(n_206),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_456),
.A2(n_256),
.B1(n_246),
.B2(n_252),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_414),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_448),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_448),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_450),
.B(n_347),
.Y(n_591)
);

BUFx6f_ASAP7_75t_SL g592 ( 
.A(n_393),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_448),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_435),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_403),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_409),
.B(n_255),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_403),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_456),
.B(n_395),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_404),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_395),
.B(n_222),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g603 ( 
.A(n_390),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_451),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_404),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_406),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_451),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_409),
.B(n_257),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_478),
.B(n_197),
.C(n_181),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_485),
.B(n_418),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_261),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_499),
.A2(n_440),
.B1(n_310),
.B2(n_211),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_496),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_467),
.B(n_260),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_467),
.B(n_202),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_499),
.A2(n_539),
.B1(n_527),
.B2(n_528),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_499),
.A2(n_527),
.B1(n_528),
.B2(n_559),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_506),
.B(n_266),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_490),
.B(n_275),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_493),
.B(n_210),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_567),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_586),
.A2(n_440),
.B1(n_310),
.B2(n_211),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_559),
.B(n_575),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_462),
.B(n_390),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_567),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_575),
.B(n_418),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_536),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_568),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_496),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_475),
.B(n_277),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_468),
.B(n_425),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_542),
.B(n_451),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_542),
.B(n_457),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_468),
.B(n_425),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_457),
.Y(n_635)
);

AND2x6_ASAP7_75t_SL g636 ( 
.A(n_537),
.B(n_349),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_475),
.B(n_280),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_484),
.B(n_201),
.C(n_200),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_586),
.A2(n_206),
.B1(n_283),
.B2(n_273),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_525),
.B(n_457),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_482),
.B(n_457),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_482),
.B(n_409),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_500),
.B(n_409),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_475),
.B(n_287),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_469),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_568),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_500),
.B(n_425),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_572),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_536),
.A2(n_249),
.B(n_300),
.C(n_283),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_469),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_573),
.B(n_261),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_573),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_494),
.A2(n_213),
.B1(n_218),
.B2(n_242),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_583),
.A2(n_305),
.B1(n_291),
.B2(n_298),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_592),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_573),
.B(n_304),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_516),
.B(n_306),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_572),
.Y(n_659)
);

O2A1O1Ixp5_ASAP7_75t_L g660 ( 
.A1(n_547),
.A2(n_455),
.B(n_453),
.C(n_438),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_533),
.B(n_597),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_533),
.B(n_409),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_597),
.B(n_213),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_505),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_546),
.B(n_307),
.Y(n_665)
);

NAND2x1_ASAP7_75t_L g666 ( 
.A(n_588),
.B(n_463),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_599),
.B(n_218),
.Y(n_667)
);

INVx8_ASAP7_75t_L g668 ( 
.A(n_592),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_599),
.B(n_242),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_586),
.A2(n_573),
.B1(n_547),
.B2(n_479),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_494),
.B(n_309),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_494),
.A2(n_249),
.B1(n_253),
.B2(n_262),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_487),
.A2(n_253),
.B1(n_262),
.B2(n_273),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_509),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_502),
.B(n_554),
.Y(n_675)
);

O2A1O1Ixp5_ASAP7_75t_L g676 ( 
.A1(n_547),
.A2(n_577),
.B(n_605),
.C(n_601),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_512),
.A2(n_300),
.B1(n_453),
.B2(n_411),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_605),
.Y(n_678)
);

BUFx8_ASAP7_75t_L g679 ( 
.A(n_565),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_606),
.B(n_487),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_606),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_489),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_489),
.B(n_501),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_554),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_586),
.A2(n_455),
.B1(n_438),
.B2(n_437),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_591),
.B(n_222),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_406),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_512),
.B(n_216),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_503),
.B(n_411),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_512),
.B(n_553),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_503),
.B(n_424),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_508),
.B(n_424),
.Y(n_692)
);

AO22x2_ASAP7_75t_L g693 ( 
.A1(n_582),
.A2(n_363),
.B1(n_349),
.B2(n_352),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_591),
.B(n_222),
.Y(n_694)
);

BUFx6f_ASAP7_75t_SL g695 ( 
.A(n_510),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_508),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_513),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_513),
.B(n_431),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_587),
.B(n_431),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_543),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_565),
.B(n_512),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_519),
.B(n_437),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_576),
.B(n_219),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_519),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_509),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_520),
.B(n_388),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_481),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_520),
.B(n_388),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_521),
.B(n_388),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_531),
.A2(n_369),
.B(n_353),
.C(n_358),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_521),
.Y(n_711)
);

O2A1O1Ixp5_ASAP7_75t_L g712 ( 
.A1(n_526),
.A2(n_388),
.B(n_392),
.C(n_416),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_526),
.B(n_529),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_529),
.B(n_534),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_481),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_534),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_523),
.B(n_220),
.Y(n_717)
);

INVx8_ASAP7_75t_L g718 ( 
.A(n_592),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_573),
.B(n_223),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_573),
.A2(n_439),
.B1(n_397),
.B2(n_229),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_538),
.B(n_392),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_538),
.A2(n_228),
.B1(n_224),
.B2(n_225),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_540),
.B(n_392),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_545),
.B(n_226),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_498),
.B(n_227),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_549),
.B(n_352),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_540),
.Y(n_727)
);

BUFx4_ASAP7_75t_L g728 ( 
.A(n_603),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_544),
.B(n_392),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_230),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_549),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_544),
.B(n_398),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_479),
.A2(n_353),
.B1(n_358),
.B2(n_360),
.Y(n_733)
);

BUFx8_ASAP7_75t_L g734 ( 
.A(n_582),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_531),
.A2(n_369),
.B(n_361),
.C(n_362),
.Y(n_735)
);

BUFx6f_ASAP7_75t_SL g736 ( 
.A(n_510),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_551),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_551),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_511),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_555),
.B(n_231),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_290),
.C(n_237),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_600),
.B(n_56),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_460),
.B(n_398),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_580),
.B(n_232),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_594),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_541),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_594),
.B(n_240),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_510),
.B(n_241),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_571),
.B(n_360),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_460),
.B(n_398),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_470),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_470),
.B(n_244),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_495),
.B(n_245),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_SL g754 ( 
.A(n_473),
.B(n_439),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_511),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_474),
.B(n_414),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_474),
.B(n_477),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_477),
.B(n_250),
.Y(n_758)
);

NOR2xp67_ASAP7_75t_L g759 ( 
.A(n_473),
.B(n_57),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_461),
.B(n_398),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_522),
.B(n_399),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_532),
.B(n_363),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_532),
.B(n_365),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_557),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_598),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_557),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_589),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_589),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_479),
.B(n_399),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_515),
.B(n_366),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_608),
.B(n_558),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_479),
.B(n_399),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_562),
.B(n_566),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_570),
.A2(n_292),
.B1(n_258),
.B2(n_263),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_514),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_578),
.B(n_251),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_514),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_584),
.B(n_264),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_684),
.B(n_620),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_682),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_696),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_620),
.B(n_479),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_697),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_695),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_749),
.B(n_367),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_627),
.Y(n_786)
);

AOI221xp5_ASAP7_75t_L g787 ( 
.A1(n_638),
.A2(n_684),
.B1(n_688),
.B2(n_730),
.C(n_724),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_704),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_653),
.B(n_616),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_612),
.A2(n_603),
.B1(n_585),
.B2(n_581),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_612),
.A2(n_479),
.B1(n_517),
.B2(n_515),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_653),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_746),
.B(n_564),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_675),
.B(n_745),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_711),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_656),
.B(n_367),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_648),
.B(n_623),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_631),
.B(n_368),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_716),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_SL g800 ( 
.A(n_638),
.B(n_286),
.C(n_265),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_727),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_651),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_653),
.B(n_564),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_690),
.A2(n_372),
.B(n_375),
.C(n_596),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_653),
.Y(n_805)
);

CKINVDCx14_ASAP7_75t_R g806 ( 
.A(n_624),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_651),
.B(n_569),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_634),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_651),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_661),
.B(n_569),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_621),
.B(n_574),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_762),
.B(n_372),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_763),
.B(n_272),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_737),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_656),
.B(n_574),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_625),
.B(n_581),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_690),
.A2(n_617),
.B1(n_765),
.B2(n_699),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_726),
.B(n_515),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_738),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_651),
.B(n_731),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_726),
.B(n_515),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_701),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_764),
.Y(n_823)
);

O2A1O1Ixp5_ASAP7_75t_L g824 ( 
.A1(n_660),
.A2(n_607),
.B(n_604),
.C(n_596),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_700),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_695),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_628),
.B(n_515),
.Y(n_827)
);

BUFx2_ASAP7_75t_SL g828 ( 
.A(n_736),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_766),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_731),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_728),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_660),
.A2(n_607),
.B(n_604),
.C(n_595),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_751),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_613),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_731),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_647),
.B(n_649),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_715),
.B(n_515),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_515),
.Y(n_838)
);

CKINVDCx11_ASAP7_75t_R g839 ( 
.A(n_636),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_629),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

AND2x4_ASAP7_75t_SL g842 ( 
.A(n_731),
.B(n_588),
.Y(n_842)
);

AND2x4_ASAP7_75t_SL g843 ( 
.A(n_715),
.B(n_588),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_670),
.B(n_483),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_745),
.B(n_276),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_615),
.B(n_724),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_615),
.B(n_278),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_664),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_646),
.B(n_517),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_646),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_734),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_707),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_678),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_674),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_670),
.B(n_707),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_776),
.A2(n_778),
.B1(n_714),
.B2(n_713),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_681),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_734),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_686),
.B(n_466),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_705),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_730),
.B(n_281),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_739),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_610),
.B(n_517),
.Y(n_863)
);

BUFx4f_ASAP7_75t_L g864 ( 
.A(n_656),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_668),
.B(n_518),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_770),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_770),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_741),
.B(n_518),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_747),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_755),
.Y(n_870)
);

AND3x2_ASAP7_75t_SL g871 ( 
.A(n_640),
.B(n_1),
.C(n_2),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_736),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_683),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_668),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_759),
.B(n_517),
.Y(n_875)
);

AND2x4_ASAP7_75t_SL g876 ( 
.A(n_720),
.B(n_466),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_694),
.B(n_466),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_668),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_622),
.B(n_483),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_718),
.B(n_535),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_666),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_775),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_754),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_642),
.B(n_517),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_609),
.B(n_463),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_679),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_622),
.B(n_483),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_718),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_676),
.B(n_483),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_SL g890 ( 
.A(n_640),
.B(n_483),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_777),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_679),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_662),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_767),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_635),
.B(n_517),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_742),
.B(n_643),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_768),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_641),
.B(n_517),
.Y(n_898)
);

OR2x6_ASAP7_75t_L g899 ( 
.A(n_718),
.B(n_693),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_644),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_757),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_743),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_R g903 ( 
.A(n_719),
.B(n_282),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_687),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_676),
.B(n_680),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_752),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_632),
.B(n_463),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_688),
.B(n_464),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_693),
.Y(n_909)
);

INVx8_ASAP7_75t_L g910 ( 
.A(n_693),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_740),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_692),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_633),
.B(n_464),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_750),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_706),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_744),
.A2(n_550),
.B1(n_535),
.B2(n_548),
.Y(n_916)
);

INVxp33_ASAP7_75t_L g917 ( 
.A(n_744),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_771),
.B(n_530),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_771),
.B(n_530),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_758),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_689),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_708),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_773),
.B(n_464),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_733),
.B(n_530),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_698),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_677),
.B(n_548),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_691),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_703),
.B(n_284),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_626),
.A2(n_491),
.B1(n_497),
.B2(n_480),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_733),
.B(n_530),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_769),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_773),
.B(n_480),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_654),
.A2(n_672),
.B1(n_611),
.B2(n_652),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_753),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_619),
.B(n_480),
.Y(n_935)
);

AND2x4_ASAP7_75t_SL g936 ( 
.A(n_685),
.B(n_655),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_614),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_663),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_709),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_671),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_721),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_748),
.B(n_550),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_725),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_702),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_685),
.B(n_491),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_667),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_669),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_723),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_618),
.B(n_491),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_772),
.B(n_729),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_717),
.B(n_630),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_658),
.B(n_552),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_732),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_650),
.B(n_497),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_756),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_673),
.A2(n_593),
.B1(n_590),
.B2(n_595),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_760),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_761),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_665),
.B(n_497),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_774),
.B(n_507),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_637),
.B(n_507),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_712),
.Y(n_962)
);

AND2x6_ASAP7_75t_L g963 ( 
.A(n_753),
.B(n_507),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_671),
.B(n_530),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_645),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_722),
.B(n_552),
.Y(n_966)
);

AND2x2_ASAP7_75t_SL g967 ( 
.A(n_657),
.B(n_590),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_710),
.B(n_299),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_712),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_735),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_779),
.B(n_593),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_812),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_792),
.A2(n_805),
.B(n_923),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_933),
.A2(n_302),
.B1(n_311),
.B2(n_471),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_846),
.A2(n_563),
.B(n_561),
.C(n_560),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_779),
.A2(n_472),
.B(n_459),
.C(n_465),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_917),
.A2(n_563),
.B(n_561),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_794),
.A2(n_560),
.B(n_556),
.C(n_471),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_830),
.Y(n_979)
);

BUFx12f_ASAP7_75t_L g980 ( 
.A(n_886),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_783),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_917),
.B(n_556),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_933),
.A2(n_459),
.B1(n_492),
.B2(n_488),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_792),
.A2(n_504),
.B(n_414),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_921),
.B(n_472),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_788),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_792),
.A2(n_504),
.B(n_419),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_792),
.A2(n_504),
.B(n_419),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_800),
.A2(n_476),
.B1(n_492),
.B2(n_488),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_805),
.A2(n_504),
.B(n_419),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_780),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_861),
.A2(n_465),
.B(n_476),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_SL g993 ( 
.A(n_878),
.B(n_504),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_794),
.A2(n_486),
.B(n_399),
.C(n_405),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_873),
.A2(n_486),
.B1(n_504),
.B2(n_416),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_937),
.A2(n_416),
.B1(n_412),
.B2(n_405),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_808),
.B(n_414),
.Y(n_997)
);

CKINVDCx10_ASAP7_75t_R g998 ( 
.A(n_839),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_912),
.B(n_416),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_806),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_809),
.B(n_419),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_825),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_795),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_889),
.A2(n_412),
.B(n_405),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_808),
.B(n_419),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_805),
.A2(n_419),
.B(n_414),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_805),
.A2(n_419),
.B(n_414),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_932),
.A2(n_419),
.B(n_414),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_781),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_799),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_921),
.B(n_405),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_925),
.A2(n_412),
.B(n_414),
.C(n_13),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_927),
.B(n_412),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_800),
.A2(n_804),
.B(n_927),
.C(n_797),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_944),
.B(n_8),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_804),
.A2(n_8),
.B(n_12),
.C(n_14),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_786),
.B(n_12),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_817),
.B(n_87),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_SL g1019 ( 
.A1(n_964),
.A2(n_905),
.B(n_889),
.C(n_918),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_904),
.B(n_15),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_855),
.A2(n_791),
.B1(n_844),
.B2(n_936),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_855),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_786),
.B(n_18),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_785),
.B(n_22),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_918),
.A2(n_919),
.B(n_964),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_937),
.B(n_23),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_919),
.A2(n_102),
.B(n_143),
.Y(n_1027)
);

OA21x2_ASAP7_75t_L g1028 ( 
.A1(n_905),
.A2(n_98),
.B(n_133),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_SL g1029 ( 
.A(n_784),
.B(n_27),
.C(n_28),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_807),
.A2(n_92),
.B(n_130),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_888),
.B(n_81),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_884),
.A2(n_72),
.B(n_127),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_782),
.A2(n_155),
.B(n_125),
.C(n_123),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_847),
.B(n_27),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_822),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_904),
.B(n_28),
.Y(n_1036)
);

AO22x1_ASAP7_75t_L g1037 ( 
.A1(n_883),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_842),
.A2(n_106),
.B(n_113),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_798),
.B(n_32),
.Y(n_1039)
);

OR2x6_ASAP7_75t_SL g1040 ( 
.A(n_826),
.B(n_35),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_938),
.B(n_38),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_818),
.B(n_109),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_789),
.A2(n_110),
.B(n_111),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_801),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_869),
.A2(n_121),
.B1(n_40),
.B2(n_42),
.Y(n_1045)
);

AO31x2_ASAP7_75t_L g1046 ( 
.A1(n_885),
.A2(n_38),
.A3(n_40),
.B(n_43),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_SL g1047 ( 
.A1(n_789),
.A2(n_844),
.B(n_879),
.C(n_887),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_814),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_830),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_813),
.B(n_806),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_893),
.B(n_900),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_833),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_824),
.A2(n_832),
.B(n_950),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_798),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_895),
.A2(n_898),
.B(n_863),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_899),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_894),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_943),
.A2(n_946),
.B(n_790),
.C(n_920),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_908),
.A2(n_856),
.B(n_890),
.C(n_885),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_901),
.B(n_958),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_824),
.A2(n_832),
.B(n_929),
.Y(n_1061)
);

BUFx8_ASAP7_75t_L g1062 ( 
.A(n_851),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_874),
.Y(n_1063)
);

AND2x4_ASAP7_75t_SL g1064 ( 
.A(n_888),
.B(n_809),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_SL g1065 ( 
.A1(n_911),
.A2(n_892),
.B1(n_831),
.B2(n_934),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_819),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_796),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_901),
.B(n_957),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_830),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_897),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_915),
.B(n_922),
.Y(n_1071)
);

BUFx8_ASAP7_75t_SL g1072 ( 
.A(n_872),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_920),
.B(n_951),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_864),
.B(n_878),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_939),
.B(n_941),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_807),
.A2(n_820),
.B(n_950),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_791),
.A2(n_909),
.B1(n_879),
.B2(n_887),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_796),
.Y(n_1078)
);

INVx6_ASAP7_75t_L g1079 ( 
.A(n_878),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_890),
.A2(n_943),
.B(n_966),
.C(n_859),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_948),
.B(n_902),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_874),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_967),
.A2(n_843),
.B(n_810),
.Y(n_1083)
);

INVx11_ASAP7_75t_L g1084 ( 
.A(n_963),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_909),
.A2(n_910),
.B1(n_947),
.B2(n_926),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_965),
.B(n_818),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_830),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_947),
.B(n_914),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_845),
.B(n_965),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_859),
.A2(n_877),
.B(n_961),
.C(n_966),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_853),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_836),
.B(n_857),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_910),
.A2(n_926),
.B1(n_821),
.B2(n_963),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_965),
.B(n_906),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_823),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_965),
.B(n_821),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_877),
.A2(n_961),
.B(n_829),
.C(n_970),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_953),
.B(n_850),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_953),
.B(n_850),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_852),
.B(n_945),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_834),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_849),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_967),
.A2(n_793),
.B(n_907),
.Y(n_1103)
);

AND2x4_ASAP7_75t_SL g1104 ( 
.A(n_867),
.B(n_865),
.Y(n_1104)
);

OR2x6_ASAP7_75t_L g1105 ( 
.A(n_828),
.B(n_910),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_913),
.A2(n_803),
.B(n_935),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_849),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_SL g1108 ( 
.A1(n_820),
.A2(n_891),
.B(n_960),
.C(n_802),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_968),
.A2(n_928),
.B(n_954),
.C(n_899),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_SL g1110 ( 
.A1(n_924),
.A2(n_930),
.B(n_955),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_SL g1111 ( 
.A(n_903),
.B(n_940),
.C(n_838),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_899),
.A2(n_924),
.B1(n_930),
.B2(n_871),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_L g1113 ( 
.A(n_878),
.B(n_858),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_SL g1114 ( 
.A1(n_796),
.A2(n_871),
.B1(n_839),
.B2(n_880),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_811),
.A2(n_816),
.B(n_942),
.C(n_827),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_864),
.B(n_866),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_852),
.B(n_802),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_962),
.A2(n_969),
.B(n_956),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_867),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_840),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_SL g1121 ( 
.A(n_949),
.B(n_959),
.C(n_803),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1059),
.A2(n_896),
.B(n_875),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_972),
.B(n_942),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1051),
.B(n_931),
.Y(n_1124)
);

AOI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_1109),
.A2(n_942),
.B(n_940),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1063),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1090),
.A2(n_896),
.B(n_875),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1055),
.A2(n_876),
.B(n_837),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1051),
.B(n_931),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1004),
.A2(n_956),
.B(n_916),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1009),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1081),
.B(n_931),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_1069),
.B(n_835),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1103),
.A2(n_837),
.B(n_931),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1105),
.B(n_880),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_1079),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1010),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1019),
.A2(n_868),
.B(n_952),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1081),
.B(n_963),
.Y(n_1139)
);

AOI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_1014),
.A2(n_952),
.B(n_882),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1087),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1071),
.B(n_963),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_1098),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1080),
.A2(n_860),
.B(n_862),
.C(n_841),
.Y(n_1144)
);

OA21x2_ASAP7_75t_L g1145 ( 
.A1(n_1061),
.A2(n_870),
.B(n_854),
.Y(n_1145)
);

AO22x2_ASAP7_75t_L g1146 ( 
.A1(n_1112),
.A2(n_835),
.B1(n_866),
.B2(n_848),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1110),
.A2(n_963),
.B(n_891),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_1053),
.A2(n_903),
.B(n_881),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1022),
.A2(n_865),
.B(n_880),
.C(n_815),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1076),
.A2(n_815),
.B(n_881),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_1079),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1002),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1044),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1092),
.B(n_867),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_1082),
.B(n_867),
.Y(n_1155)
);

OAI22x1_ASAP7_75t_L g1156 ( 
.A1(n_1026),
.A2(n_865),
.B1(n_815),
.B2(n_881),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1024),
.B(n_1054),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1083),
.A2(n_1025),
.B(n_1106),
.Y(n_1158)
);

OAI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1073),
.A2(n_1034),
.B(n_1089),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1048),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1115),
.A2(n_1118),
.B(n_1047),
.Y(n_1161)
);

AOI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1018),
.A2(n_971),
.B(n_1008),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1000),
.Y(n_1163)
);

OAI22x1_ASAP7_75t_L g1164 ( 
.A1(n_1056),
.A2(n_1094),
.B1(n_1045),
.B2(n_1023),
.Y(n_1164)
);

AO22x2_ASAP7_75t_L g1165 ( 
.A1(n_1112),
.A2(n_1022),
.B1(n_1077),
.B2(n_1021),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1039),
.B(n_1050),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1075),
.B(n_1060),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_1077),
.A2(n_1021),
.B(n_1016),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1068),
.B(n_1088),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1066),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1058),
.B(n_1015),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1035),
.B(n_981),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1017),
.A2(n_974),
.B1(n_1037),
.B2(n_1114),
.C(n_1095),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1091),
.B(n_985),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1041),
.B(n_1020),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1118),
.A2(n_1111),
.B(n_973),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1053),
.A2(n_1121),
.B(n_994),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1108),
.A2(n_975),
.B(n_978),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1099),
.A2(n_1100),
.B(n_992),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1085),
.A2(n_1093),
.B1(n_1036),
.B2(n_1084),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1116),
.B(n_1096),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_986),
.B(n_1052),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1003),
.B(n_1057),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1070),
.B(n_1107),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1101),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1102),
.B(n_1107),
.Y(n_1186)
);

AO32x2_ASAP7_75t_L g1187 ( 
.A1(n_974),
.A2(n_995),
.A3(n_983),
.B1(n_1046),
.B2(n_1065),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1120),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1072),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1033),
.A2(n_1012),
.B(n_1032),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1031),
.A2(n_1043),
.B(n_1038),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1067),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1078),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1086),
.B(n_1029),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1069),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_982),
.B(n_1011),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_983),
.A2(n_1030),
.B(n_995),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_984),
.A2(n_987),
.B(n_988),
.Y(n_1198)
);

OAI21xp33_ASAP7_75t_L g1199 ( 
.A1(n_1013),
.A2(n_1105),
.B(n_999),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_976),
.A2(n_999),
.B(n_1027),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_990),
.A2(n_1006),
.B(n_1007),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1001),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1069),
.A2(n_1005),
.B(n_997),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1087),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_977),
.A2(n_1117),
.B(n_1049),
.C(n_979),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1069),
.A2(n_977),
.B(n_1028),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_989),
.A2(n_1001),
.B(n_1028),
.Y(n_1207)
);

AO21x1_ASAP7_75t_L g1208 ( 
.A1(n_996),
.A2(n_1104),
.B(n_1031),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1102),
.B(n_1105),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_979),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1046),
.A2(n_1113),
.B(n_993),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1049),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1119),
.B(n_1087),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1046),
.A2(n_1042),
.A3(n_1119),
.B(n_1074),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1064),
.B(n_1119),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1042),
.A2(n_1062),
.B(n_1040),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1042),
.A2(n_1062),
.B(n_980),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1042),
.A2(n_1059),
.B(n_1090),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_998),
.A2(n_1004),
.B(n_1076),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_1098),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1059),
.A2(n_787),
.B(n_846),
.C(n_779),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1059),
.A2(n_1080),
.A3(n_1097),
.B(n_1112),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_972),
.B(n_917),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1059),
.A2(n_1019),
.B(n_1080),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_991),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1059),
.A2(n_787),
.B(n_846),
.C(n_779),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1059),
.A2(n_1019),
.B(n_1080),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1073),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_972),
.B(n_468),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1059),
.A2(n_787),
.B(n_846),
.C(n_779),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1051),
.B(n_873),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1116),
.B(n_1086),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_991),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_972),
.B(n_762),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_991),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1059),
.A2(n_805),
.B(n_792),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_972),
.B(n_762),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1051),
.A2(n_612),
.B1(n_499),
.B2(n_933),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1051),
.B(n_873),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1051),
.B(n_779),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1059),
.A2(n_787),
.B(n_846),
.C(n_779),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1051),
.B(n_779),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1059),
.A2(n_1019),
.B(n_1080),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1051),
.B(n_779),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1072),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1051),
.B(n_873),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_991),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_SL g1253 ( 
.A(n_1114),
.B(n_499),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1050),
.A2(n_620),
.B1(n_537),
.B2(n_846),
.Y(n_1254)
);

NOR2x1_ASAP7_75t_L g1255 ( 
.A(n_1063),
.B(n_888),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_991),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1002),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1059),
.A2(n_805),
.B(n_792),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_972),
.B(n_762),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1059),
.A2(n_1080),
.B(n_1097),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1004),
.A2(n_1076),
.B(n_1061),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1059),
.A2(n_787),
.B(n_846),
.C(n_779),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1059),
.A2(n_620),
.B(n_846),
.C(n_787),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1059),
.A2(n_805),
.B(n_792),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1079),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1002),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_SL g1268 ( 
.A1(n_1109),
.A2(n_909),
.B(n_1058),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1059),
.A2(n_1080),
.A3(n_1097),
.B(n_1112),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1002),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1051),
.A2(n_612),
.B1(n_499),
.B2(n_933),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1189),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1267),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_1152),
.B(n_1136),
.Y(n_1274)
);

AO21x2_ASAP7_75t_L g1275 ( 
.A1(n_1125),
.A2(n_1176),
.B(n_1178),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1168),
.A2(n_1253),
.B1(n_1165),
.B2(n_1271),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1145),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1157),
.B(n_1166),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1227),
.A2(n_1240),
.B(n_1232),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1136),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1246),
.A2(n_1256),
.B(n_1250),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1241),
.A2(n_1271),
.B(n_1231),
.C(n_1263),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1243),
.B(n_1245),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1262),
.A2(n_1201),
.B(n_1198),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1249),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1136),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1270),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1266),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1158),
.A2(n_1150),
.B(n_1197),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1248),
.B(n_1233),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1137),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1254),
.A2(n_1253),
.B1(n_1175),
.B2(n_1159),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_SL g1293 ( 
.A1(n_1241),
.A2(n_1244),
.B(n_1221),
.C(n_1226),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1125),
.A2(n_1178),
.B(n_1161),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_L g1295 ( 
.A1(n_1264),
.A2(n_1173),
.B1(n_1261),
.B2(n_1229),
.C(n_1165),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1171),
.B(n_1194),
.C(n_1223),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1130),
.A2(n_1207),
.B(n_1134),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1233),
.A2(n_1251),
.B1(n_1242),
.B2(n_1239),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1153),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1149),
.B(n_1191),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1224),
.A2(n_1228),
.B(n_1247),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_SL g1302 ( 
.A(n_1216),
.B(n_1242),
.C(n_1251),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1206),
.A2(n_1122),
.B(n_1147),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1179),
.A2(n_1127),
.A3(n_1208),
.B(n_1259),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1126),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1138),
.A2(n_1200),
.B(n_1140),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1200),
.A2(n_1140),
.B(n_1162),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1128),
.A2(n_1265),
.B(n_1238),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1219),
.A2(n_1205),
.B(n_1139),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1160),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1139),
.A2(n_1142),
.B(n_1190),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1142),
.A2(n_1190),
.B(n_1203),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1199),
.A2(n_1220),
.B(n_1143),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1129),
.A2(n_1124),
.B(n_1132),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1266),
.B(n_1195),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1167),
.B(n_1169),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1131),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1167),
.B(n_1169),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1148),
.A2(n_1144),
.B(n_1218),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1132),
.A2(n_1154),
.B(n_1174),
.C(n_1225),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1177),
.A2(n_1218),
.B(n_1180),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1266),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1235),
.A2(n_1252),
.B(n_1237),
.C(n_1257),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1236),
.A2(n_1260),
.B1(n_1180),
.B2(n_1234),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1177),
.A2(n_1146),
.B(n_1156),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_1230),
.B(n_1186),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1188),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1183),
.B(n_1182),
.C(n_1234),
.Y(n_1329)
);

CKINVDCx6p67_ASAP7_75t_R g1330 ( 
.A(n_1267),
.Y(n_1330)
);

OAI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1163),
.A2(n_1123),
.B1(n_1193),
.B2(n_1192),
.C(n_1172),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1151),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1184),
.A2(n_1181),
.B(n_1202),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1210),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1211),
.A2(n_1133),
.B(n_1209),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1211),
.A2(n_1133),
.B(n_1212),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1258),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1213),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1269),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1269),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1164),
.B(n_1217),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1155),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1269),
.Y(n_1343)
);

BUFx8_ASAP7_75t_L g1344 ( 
.A(n_1215),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1213),
.A2(n_1146),
.B(n_1204),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1217),
.B(n_1151),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1255),
.A2(n_1195),
.B(n_1215),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1222),
.B(n_1135),
.Y(n_1348)
);

NOR2x1_ASAP7_75t_SL g1349 ( 
.A(n_1135),
.B(n_1141),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1135),
.B(n_1141),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1214),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1214),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1187),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1187),
.A2(n_1168),
.A3(n_1161),
.B(n_1176),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1126),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1168),
.A2(n_787),
.B1(n_846),
.B2(n_779),
.Y(n_1356)
);

NOR3xp33_ASAP7_75t_SL g1357 ( 
.A(n_1159),
.B(n_473),
.C(n_402),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1157),
.B(n_1166),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1243),
.B(n_1245),
.Y(n_1359)
);

AOI22x1_ASAP7_75t_L g1360 ( 
.A1(n_1164),
.A2(n_846),
.B1(n_1156),
.B2(n_861),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1159),
.B(n_620),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1168),
.A2(n_787),
.B1(n_846),
.B2(n_779),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1145),
.Y(n_1364)
);

BUFx2_ASAP7_75t_SL g1365 ( 
.A(n_1136),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1227),
.A2(n_1240),
.B(n_1232),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1189),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1227),
.A2(n_1240),
.B(n_1232),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1145),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1168),
.A2(n_1161),
.A3(n_1176),
.B(n_1059),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1145),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1159),
.B(n_620),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1136),
.B(n_1266),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_SL g1375 ( 
.A1(n_1241),
.A2(n_1271),
.B(n_1226),
.C(n_1231),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1243),
.B(n_1245),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1125),
.A2(n_1176),
.B(n_1178),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1125),
.A2(n_1176),
.B(n_1178),
.Y(n_1378)
);

OAI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1254),
.A2(n_787),
.B1(n_620),
.B2(n_493),
.C(n_730),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1152),
.B(n_1136),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1137),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1227),
.A2(n_1240),
.B(n_1232),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1264),
.A2(n_620),
.B(n_846),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1137),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1268),
.A2(n_1208),
.B(n_1149),
.Y(n_1385)
);

AO31x2_ASAP7_75t_L g1386 ( 
.A1(n_1168),
.A2(n_1161),
.A3(n_1176),
.B(n_1059),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1224),
.A2(n_1247),
.B(n_1228),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1268),
.A2(n_1208),
.B(n_1149),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1254),
.A2(n_1243),
.B1(n_1248),
.B2(n_1245),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1224),
.A2(n_1247),
.B(n_1228),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1264),
.A2(n_620),
.B(n_846),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1258),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1268),
.A2(n_1208),
.B(n_1149),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1189),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1125),
.A2(n_1176),
.B(n_1178),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1137),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1243),
.B(n_1245),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1267),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1145),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_L g1401 ( 
.A(n_1264),
.B(n_620),
.C(n_787),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1159),
.B(n_620),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1224),
.A2(n_1247),
.B(n_1228),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1137),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1136),
.B(n_1266),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1168),
.A2(n_1161),
.A3(n_1176),
.B(n_1059),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1379),
.A2(n_1392),
.B(n_1383),
.C(n_1373),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_SL g1408 ( 
.A(n_1300),
.B(n_1302),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1292),
.A2(n_1363),
.B1(n_1356),
.B2(n_1401),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1278),
.B(n_1358),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1300),
.A2(n_1318),
.B(n_1316),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1356),
.A2(n_1363),
.B1(n_1296),
.B2(n_1357),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1283),
.A2(n_1376),
.B1(n_1359),
.B2(n_1398),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1362),
.A2(n_1373),
.B(n_1402),
.C(n_1295),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1361),
.B(n_1367),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1362),
.A2(n_1402),
.B1(n_1276),
.B2(n_1290),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1276),
.A2(n_1331),
.B1(n_1342),
.B2(n_1390),
.Y(n_1417)
);

BUFx4f_ASAP7_75t_L g1418 ( 
.A(n_1286),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1298),
.B(n_1388),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1327),
.B(n_1338),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1273),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1325),
.B(n_1310),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1300),
.A2(n_1293),
.B(n_1282),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1313),
.A2(n_1329),
.B(n_1321),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1293),
.A2(n_1375),
.B(n_1282),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1375),
.A2(n_1385),
.B(n_1394),
.C(n_1389),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_R g1427 ( 
.A(n_1280),
.B(n_1272),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1393),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1329),
.A2(n_1321),
.B(n_1374),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1317),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1314),
.B(n_1348),
.Y(n_1431)
);

OAI211xp5_ASAP7_75t_L g1432 ( 
.A1(n_1360),
.A2(n_1324),
.B(n_1333),
.C(n_1347),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1324),
.A2(n_1399),
.B(n_1350),
.C(n_1341),
.Y(n_1433)
);

BUFx2_ASAP7_75t_SL g1434 ( 
.A(n_1274),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1314),
.B(n_1328),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1330),
.A2(n_1353),
.B1(n_1286),
.B2(n_1323),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1349),
.B(n_1346),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1314),
.B(n_1291),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1277),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1299),
.B(n_1381),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1384),
.B(n_1397),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_R g1442 ( 
.A(n_1285),
.B(n_1395),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1374),
.A2(n_1405),
.B(n_1280),
.Y(n_1443)
);

BUFx10_ASAP7_75t_L g1444 ( 
.A(n_1305),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1285),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1404),
.B(n_1337),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1326),
.A2(n_1320),
.B(n_1339),
.C(n_1340),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1353),
.A2(n_1303),
.B(n_1343),
.C(n_1339),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1330),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1319),
.A2(n_1315),
.B(n_1355),
.C(n_1294),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1337),
.A2(n_1380),
.B1(n_1315),
.B2(n_1405),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1365),
.A2(n_1332),
.B1(n_1288),
.B2(n_1301),
.Y(n_1452)
);

O2A1O1Ixp5_ASAP7_75t_L g1453 ( 
.A1(n_1352),
.A2(n_1334),
.B(n_1372),
.C(n_1364),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1303),
.A2(n_1289),
.B(n_1312),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1308),
.A2(n_1311),
.B(n_1309),
.C(n_1312),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1371),
.B(n_1386),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1301),
.A2(n_1387),
.B1(n_1403),
.B2(n_1391),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1371),
.B(n_1406),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1345),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1294),
.A2(n_1378),
.B(n_1275),
.C(n_1396),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1371),
.B(n_1406),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1351),
.B(n_1335),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1395),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1275),
.A2(n_1378),
.B(n_1377),
.C(n_1396),
.Y(n_1465)
);

O2A1O1Ixp5_ASAP7_75t_L g1466 ( 
.A1(n_1370),
.A2(n_1400),
.B(n_1371),
.C(n_1406),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1344),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1301),
.B(n_1403),
.Y(n_1468)
);

O2A1O1Ixp5_ASAP7_75t_L g1469 ( 
.A1(n_1386),
.A2(n_1354),
.B(n_1306),
.C(n_1304),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1311),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1309),
.A2(n_1297),
.B(n_1386),
.C(n_1354),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1289),
.A2(n_1284),
.B(n_1297),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1354),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1344),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1354),
.B(n_1391),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1387),
.B(n_1322),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1307),
.A2(n_1304),
.B(n_1344),
.C(n_1287),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1307),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1279),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1272),
.A2(n_1368),
.B(n_1284),
.C(n_1281),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1279),
.B(n_1281),
.Y(n_1481)
);

CKINVDCx6p67_ASAP7_75t_R g1482 ( 
.A(n_1366),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1366),
.B(n_1369),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1382),
.B(n_1361),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1383),
.A2(n_1271),
.B(n_1241),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1383),
.A2(n_1271),
.B(n_1241),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1379),
.A2(n_1254),
.B1(n_1292),
.B2(n_1356),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1278),
.B(n_1358),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1361),
.B(n_1367),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1320),
.A2(n_1303),
.B(n_1228),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1285),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1379),
.A2(n_620),
.B(n_1392),
.C(n_1383),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1379),
.A2(n_1254),
.B1(n_1292),
.B2(n_1356),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1439),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1438),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1492),
.A2(n_1407),
.B(n_1414),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1461),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1435),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1414),
.A2(n_1493),
.B(n_1487),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1468),
.B(n_1476),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1446),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_R g1502 ( 
.A(n_1445),
.B(n_1464),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1481),
.B(n_1483),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1431),
.B(n_1475),
.Y(n_1504)
);

INVx4_ASAP7_75t_SL g1505 ( 
.A(n_1463),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1459),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1459),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1482),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1485),
.A2(n_1486),
.B(n_1455),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1454),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1411),
.B(n_1419),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1454),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1454),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1412),
.B(n_1416),
.C(n_1409),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1466),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1436),
.A2(n_1417),
.B1(n_1423),
.B2(n_1425),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1472),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1424),
.B(n_1429),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1470),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1415),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1472),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1437),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1478),
.B(n_1456),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1455),
.A2(n_1465),
.B(n_1460),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1490),
.B(n_1471),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1490),
.B(n_1471),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1478),
.B(n_1462),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1458),
.B(n_1469),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1479),
.B(n_1447),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1472),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1437),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1453),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1430),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1408),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1520),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1510),
.B(n_1491),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1537),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1494),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1537),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1502),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1500),
.B(n_1410),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1495),
.B(n_1420),
.Y(n_1546)
);

NOR2x1_ASAP7_75t_L g1547 ( 
.A(n_1521),
.B(n_1450),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1516),
.B(n_1428),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1488),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1521),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1522),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1497),
.B(n_1441),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1502),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1495),
.B(n_1489),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1521),
.B(n_1452),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1499),
.A2(n_1413),
.B1(n_1474),
.B2(n_1421),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1521),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1522),
.Y(n_1558)
);

NAND2x1_ASAP7_75t_L g1559 ( 
.A(n_1521),
.B(n_1443),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1518),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1521),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1426),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1508),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1516),
.A2(n_1432),
.B1(n_1449),
.B2(n_1433),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1503),
.B(n_1422),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1513),
.B(n_1440),
.Y(n_1567)
);

OAI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1565),
.A2(n_1499),
.B1(n_1496),
.B2(n_1513),
.C(n_1531),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1541),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1560),
.A2(n_1515),
.B(n_1512),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

NAND4xp25_ASAP7_75t_L g1573 ( 
.A(n_1548),
.B(n_1496),
.C(n_1519),
.D(n_1523),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

OAI31xp33_ASAP7_75t_L g1575 ( 
.A1(n_1565),
.A2(n_1548),
.A3(n_1556),
.B(n_1451),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1566),
.B(n_1504),
.Y(n_1576)
);

OAI33xp33_ASAP7_75t_L g1577 ( 
.A1(n_1567),
.A2(n_1504),
.A3(n_1530),
.B1(n_1526),
.B2(n_1498),
.B3(n_1506),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1556),
.B(n_1519),
.C(n_1531),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1567),
.B(n_1523),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1559),
.Y(n_1580)
);

OAI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1531),
.B1(n_1555),
.B2(n_1559),
.C(n_1563),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1551),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1554),
.B(n_1501),
.Y(n_1584)
);

AOI33xp33_ASAP7_75t_L g1585 ( 
.A1(n_1541),
.A2(n_1532),
.A3(n_1528),
.B1(n_1529),
.B2(n_1533),
.B3(n_1498),
.Y(n_1585)
);

OAI31xp33_ASAP7_75t_L g1586 ( 
.A1(n_1550),
.A2(n_1507),
.A3(n_1509),
.B(n_1528),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1546),
.A2(n_1511),
.B1(n_1518),
.B2(n_1501),
.C(n_1532),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1543),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1563),
.A2(n_1531),
.B1(n_1467),
.B2(n_1418),
.Y(n_1590)
);

OAI321xp33_ASAP7_75t_L g1591 ( 
.A1(n_1563),
.A2(n_1531),
.A3(n_1528),
.B1(n_1529),
.B2(n_1506),
.C(n_1533),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1558),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1546),
.A2(n_1511),
.B1(n_1518),
.B2(n_1532),
.C(n_1533),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1558),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1564),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_R g1599 ( 
.A(n_1544),
.B(n_1418),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1563),
.A2(n_1511),
.B1(n_1531),
.B2(n_1474),
.Y(n_1600)
);

AOI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1539),
.A2(n_1524),
.B(n_1534),
.Y(n_1601)
);

AOI33xp33_ASAP7_75t_L g1602 ( 
.A1(n_1566),
.A2(n_1529),
.A3(n_1509),
.B1(n_1507),
.B2(n_1536),
.B3(n_1517),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1564),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1504),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1542),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1563),
.A2(n_1467),
.B1(n_1525),
.B2(n_1535),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1580),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1601),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1570),
.Y(n_1609)
);

AND4x1_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1547),
.C(n_1555),
.D(n_1427),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1594),
.B(n_1553),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1574),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1571),
.A2(n_1524),
.B(n_1534),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1568),
.A2(n_1563),
.B(n_1559),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1589),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1592),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1605),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1597),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1583),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1569),
.B(n_1582),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1594),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1561),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1600),
.A2(n_1514),
.B(n_1512),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1598),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1569),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1603),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1593),
.Y(n_1627)
);

INVx4_ASAP7_75t_SL g1628 ( 
.A(n_1580),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1579),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1569),
.B(n_1505),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1588),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1599),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1604),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1582),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1581),
.B(n_1563),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1587),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1572),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1636),
.B(n_1585),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1636),
.B(n_1585),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1613),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1613),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1625),
.B(n_1602),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1629),
.B(n_1602),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1610),
.A2(n_1578),
.B(n_1573),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1609),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1629),
.B(n_1545),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1634),
.B(n_1582),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1620),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1615),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1615),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1616),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1618),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1614),
.A2(n_1511),
.B1(n_1600),
.B2(n_1557),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1632),
.B(n_1591),
.C(n_1577),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1610),
.A2(n_1590),
.B(n_1586),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1614),
.B(n_1606),
.C(n_1584),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1616),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1617),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1635),
.B(n_1557),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1617),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1608),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1624),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1624),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1608),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1637),
.B(n_1620),
.Y(n_1668)
);

NAND2x1_ASAP7_75t_L g1669 ( 
.A(n_1620),
.B(n_1580),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1645),
.A2(n_1635),
.B(n_1632),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1650),
.B(n_1620),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1645),
.A2(n_1621),
.B1(n_1630),
.B2(n_1511),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1658),
.A2(n_1621),
.B1(n_1630),
.B2(n_1620),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1650),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1638),
.B(n_1633),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

OAI32xp33_ASAP7_75t_L g1677 ( 
.A1(n_1638),
.A2(n_1619),
.A3(n_1627),
.B1(n_1622),
.B2(n_1626),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1642),
.Y(n_1678)
);

NAND2x1_ASAP7_75t_SL g1679 ( 
.A(n_1643),
.B(n_1630),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1647),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1644),
.B(n_1633),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1630),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1652),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1668),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1643),
.B(n_1630),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1639),
.B(n_1657),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1611),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1658),
.A2(n_1612),
.B(n_1627),
.C(n_1608),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1644),
.A2(n_1557),
.B1(n_1562),
.B2(n_1550),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1655),
.B(n_1607),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1434),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1655),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1668),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1653),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1668),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1653),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1549),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1646),
.Y(n_1700)
);

AOI21xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1662),
.A2(n_1623),
.B(n_1599),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1659),
.A2(n_1623),
.B(n_1612),
.C(n_1550),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1654),
.Y(n_1703)
);

AOI21xp33_ASAP7_75t_L g1704 ( 
.A1(n_1656),
.A2(n_1607),
.B(n_1623),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1662),
.B(n_1628),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1676),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1689),
.B(n_1669),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1700),
.B(n_1665),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1674),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1678),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1679),
.Y(n_1711)
);

CKINVDCx16_ASAP7_75t_R g1712 ( 
.A(n_1688),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1674),
.B(n_1671),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1671),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1689),
.B(n_1646),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1683),
.B(n_1649),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1670),
.A2(n_1646),
.B1(n_1662),
.B2(n_1527),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_L g1718 ( 
.A(n_1690),
.B(n_1664),
.C(n_1667),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1683),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1680),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1686),
.B(n_1649),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1694),
.B(n_1648),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1686),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1699),
.B(n_1665),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1705),
.B(n_1649),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1681),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1705),
.B(n_1651),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1685),
.Y(n_1729)
);

AOI222xp33_ASAP7_75t_L g1730 ( 
.A1(n_1677),
.A2(n_1702),
.B1(n_1675),
.B2(n_1692),
.C1(n_1691),
.C2(n_1698),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1712),
.B(n_1673),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1709),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1713),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1692),
.Y(n_1735)
);

AOI321xp33_ASAP7_75t_L g1736 ( 
.A1(n_1715),
.A2(n_1672),
.A3(n_1702),
.B1(n_1704),
.B2(n_1701),
.C(n_1697),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1716),
.B(n_1693),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1714),
.B(n_1685),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1716),
.B(n_1693),
.Y(n_1739)
);

OAI31xp33_ASAP7_75t_L g1740 ( 
.A1(n_1711),
.A2(n_1682),
.A3(n_1697),
.B(n_1695),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1730),
.A2(n_1662),
.B1(n_1693),
.B2(n_1695),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1708),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1717),
.A2(n_1662),
.B1(n_1607),
.B2(n_1648),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1708),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1717),
.A2(n_1662),
.B(n_1703),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1713),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1707),
.B(n_1722),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1718),
.A2(n_1442),
.B(n_1696),
.C(n_1687),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1733),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1731),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1735),
.B(n_1719),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1733),
.B(n_1719),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1738),
.B(n_1723),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1748),
.B(n_1723),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1742),
.Y(n_1757)
);

NOR2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1732),
.B(n_1725),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1731),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1742),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1741),
.B(n_1724),
.C(n_1718),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1747),
.B(n_1750),
.Y(n_1762)
);

OAI21xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1758),
.A2(n_1740),
.B(n_1739),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_L g1764 ( 
.A1(n_1753),
.A2(n_1750),
.B(n_1744),
.C(n_1749),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1759),
.B(n_1734),
.Y(n_1765)
);

NAND4xp25_ASAP7_75t_L g1766 ( 
.A(n_1756),
.B(n_1736),
.C(n_1743),
.D(n_1734),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_L g1767 ( 
.A1(n_1759),
.A2(n_1745),
.B(n_1724),
.C(n_1746),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1755),
.A2(n_1725),
.B1(n_1739),
.B2(n_1737),
.C(n_1745),
.Y(n_1768)
);

AND3x1_ASAP7_75t_L g1769 ( 
.A(n_1752),
.B(n_1737),
.C(n_1746),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1751),
.B(n_1726),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1765),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1770),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1769),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1767),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1768),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_R g1776 ( 
.A(n_1773),
.B(n_1757),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1772),
.B(n_1762),
.Y(n_1777)
);

NOR2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1771),
.B(n_1772),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1774),
.B(n_1754),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1775),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1772),
.B(n_1760),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1779),
.B(n_1777),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_L g1783 ( 
.A(n_1780),
.B(n_1763),
.C(n_1766),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1778),
.A2(n_1764),
.B1(n_1726),
.B2(n_1728),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1776),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1781),
.Y(n_1786)
);

NOR2x1_ASAP7_75t_L g1787 ( 
.A(n_1786),
.B(n_1781),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1782),
.B(n_1706),
.Y(n_1788)
);

AOI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1783),
.A2(n_1720),
.B(n_1706),
.C(n_1727),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1788),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1790),
.B(n_1784),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1785),
.B1(n_1787),
.B2(n_1789),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1791),
.Y(n_1793)
);

OAI22x1_ASAP7_75t_L g1794 ( 
.A1(n_1792),
.A2(n_1710),
.B1(n_1720),
.B2(n_1727),
.Y(n_1794)
);

OAI22x1_ASAP7_75t_L g1795 ( 
.A1(n_1793),
.A2(n_1710),
.B1(n_1729),
.B2(n_1728),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1795),
.A2(n_1664),
.B1(n_1667),
.B2(n_1721),
.C(n_1666),
.Y(n_1796)
);

AO22x2_ASAP7_75t_L g1797 ( 
.A1(n_1794),
.A2(n_1721),
.B1(n_1667),
.B2(n_1664),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_1666),
.B1(n_1654),
.B2(n_1660),
.Y(n_1798)
);

OA22x2_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1797),
.B1(n_1640),
.B2(n_1641),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1660),
.B(n_1442),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1800),
.Y(n_1801)
);

AOI31xp33_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_1444),
.A3(n_1540),
.B(n_1663),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1540),
.B(n_1663),
.C(n_1661),
.Y(n_1803)
);


endmodule