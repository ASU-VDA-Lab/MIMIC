module fake_jpeg_2790_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_49),
.B1(n_36),
.B2(n_44),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_41),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_43),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_70),
.C(n_77),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_44),
.B1(n_46),
.B2(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_46),
.C(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_80),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_6),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_4),
.Y(n_100)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_17),
.C(n_30),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_101),
.C(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_107),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_19),
.B(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_15),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_109),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_8),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_34),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.C(n_22),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_117),
.A3(n_115),
.B1(n_111),
.B2(n_118),
.C1(n_112),
.C2(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_120),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_126),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_134),
.B(n_131),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_124),
.B(n_119),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_138),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_129),
.C(n_25),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);


endmodule