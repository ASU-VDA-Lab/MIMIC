module fake_jpeg_1422_n_176 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_48),
.B1(n_50),
.B2(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_54),
.B1(n_49),
.B2(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_44),
.B(n_47),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_93),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_19),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_49),
.B1(n_55),
.B2(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_54),
.B1(n_59),
.B2(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_69),
.B1(n_46),
.B2(n_52),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_110),
.B1(n_6),
.B2(n_8),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_102),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_69),
.C(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_21),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_90),
.B(n_52),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_9),
.B(n_10),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_5),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_6),
.Y(n_126)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_131),
.B(n_23),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_126),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_132),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_28),
.B1(n_37),
.B2(n_35),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_101),
.C(n_97),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_147),
.C(n_125),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_114),
.B(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_11),
.B(n_12),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_40),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_131),
.B(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_153),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_158),
.B1(n_147),
.B2(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_164),
.B(n_156),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_166),
.B1(n_160),
.B2(n_149),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_151),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_167),
.A2(n_138),
.B(n_162),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_169),
.B1(n_161),
.B2(n_141),
.Y(n_170)
);

AOI31xp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_158),
.A3(n_144),
.B(n_141),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_15),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_16),
.C(n_18),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_33),
.Y(n_176)
);


endmodule