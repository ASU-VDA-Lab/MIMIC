module fake_jpeg_877_n_528 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_0),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_59),
.Y(n_165)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_69),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_0),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_89),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_0),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_18),
.B(n_1),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_29),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_22),
.B1(n_38),
.B2(n_29),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_35),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_96),
.B1(n_103),
.B2(n_53),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_107),
.A2(n_144),
.B1(n_26),
.B2(n_27),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_32),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_118),
.Y(n_175)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_56),
.B(n_91),
.CON(n_117),
.SN(n_117)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_117),
.A2(n_142),
.B(n_36),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_32),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_120),
.B(n_31),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_61),
.A2(n_24),
.B1(n_21),
.B2(n_45),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_129),
.B1(n_132),
.B2(n_160),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_63),
.A2(n_24),
.B1(n_45),
.B2(n_42),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_45),
.B1(n_42),
.B2(n_40),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_40),
.B(n_38),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_67),
.A2(n_17),
.B(n_46),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_33),
.CI(n_36),
.CON(n_179),
.SN(n_179)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_76),
.A2(n_79),
.B1(n_88),
.B2(n_86),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_48),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_108),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_170),
.B(n_173),
.Y(n_232)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_56),
.B1(n_87),
.B2(n_75),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_172),
.A2(n_193),
.B1(n_203),
.B2(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_179),
.A2(n_164),
.B(n_123),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_31),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_183),
.B(n_189),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_194),
.Y(n_222)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_190),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_70),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_90),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_129),
.A2(n_50),
.B1(n_71),
.B2(n_72),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_121),
.A2(n_105),
.B1(n_80),
.B2(n_78),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_198),
.Y(n_226)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_146),
.B(n_46),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_107),
.A2(n_84),
.B1(n_64),
.B2(n_26),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_208),
.B1(n_137),
.B2(n_153),
.Y(n_242)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_109),
.B(n_27),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_43),
.B1(n_36),
.B2(n_33),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_209),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_207),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_142),
.A2(n_43),
.B1(n_30),
.B2(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_138),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_211),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_135),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_125),
.B(n_43),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_216),
.Y(n_250)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_153),
.A2(n_30),
.B1(n_2),
.B2(n_5),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_114),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_220),
.B(n_231),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_165),
.B(n_117),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_221),
.A2(n_126),
.B(n_122),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g228 ( 
.A(n_170),
.B(n_161),
.C(n_137),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_187),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_133),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_179),
.A2(n_164),
.B(n_154),
.C(n_165),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_240),
.B(n_248),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_214),
.B1(n_192),
.B2(n_191),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_168),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_175),
.B(n_145),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_173),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_181),
.B1(n_186),
.B2(n_193),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_261),
.B1(n_262),
.B2(n_267),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_222),
.A2(n_179),
.B(n_194),
.C(n_181),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_260),
.A2(n_236),
.B(n_224),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_203),
.B1(n_197),
.B2(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_245),
.Y(n_265)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_194),
.B1(n_158),
.B2(n_182),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_194),
.B1(n_112),
.B2(n_158),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_242),
.B1(n_229),
.B2(n_244),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_280),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_271),
.B(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_174),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_216),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_226),
.B(n_171),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_219),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_279),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_252),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_162),
.B1(n_135),
.B2(n_167),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_281),
.A2(n_239),
.B1(n_234),
.B2(n_250),
.Y(n_311)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_221),
.B(n_240),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_215),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_307),
.B1(n_269),
.B2(n_260),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_266),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_291),
.B(n_309),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_294),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_231),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_308),
.C(n_257),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_236),
.B1(n_228),
.B2(n_229),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_302),
.A2(n_305),
.B1(n_315),
.B2(n_281),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_267),
.A2(n_236),
.B1(n_238),
.B2(n_226),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_232),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_256),
.B(n_272),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_311),
.A2(n_270),
.B1(n_282),
.B2(n_285),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_248),
.B1(n_249),
.B2(n_224),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_278),
.B(n_264),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_316),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_342),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_312),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_327),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_286),
.A2(n_284),
.B1(n_260),
.B2(n_262),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_286),
.A2(n_269),
.B1(n_278),
.B2(n_260),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_287),
.A2(n_277),
.B1(n_273),
.B2(n_283),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_275),
.Y(n_328)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_307),
.A2(n_283),
.B1(n_262),
.B2(n_256),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_336),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_307),
.A2(n_263),
.B1(n_274),
.B2(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_339),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_265),
.B1(n_279),
.B2(n_255),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_337),
.A2(n_321),
.B1(n_329),
.B2(n_326),
.Y(n_359)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_297),
.A2(n_298),
.B1(n_311),
.B2(n_295),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_345),
.B1(n_293),
.B2(n_306),
.Y(n_372)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_293),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_294),
.A2(n_247),
.B(n_250),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_233),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_346),
.C(n_304),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_302),
.A2(n_279),
.B1(n_241),
.B2(n_253),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_295),
.A2(n_232),
.B(n_233),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_322),
.A2(n_289),
.B1(n_299),
.B2(n_313),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_348),
.A2(n_364),
.B1(n_376),
.B2(n_227),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_308),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_351),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_343),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_365),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_299),
.Y(n_351)
);

OA22x2_ASAP7_75t_L g354 ( 
.A1(n_317),
.A2(n_315),
.B1(n_314),
.B2(n_310),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_374),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_357),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_343),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_359),
.A2(n_337),
.B1(n_324),
.B2(n_327),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_344),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_227),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_340),
.A2(n_291),
.B1(n_310),
.B2(n_301),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_328),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_366),
.Y(n_391)
);

XNOR2x2_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_296),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_128),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_312),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_375),
.C(n_333),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_300),
.B1(n_241),
.B2(n_255),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_300),
.B1(n_241),
.B2(n_255),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_247),
.C(n_239),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_324),
.A2(n_303),
.B1(n_253),
.B2(n_235),
.Y(n_376)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_378),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_379),
.A2(n_348),
.B1(n_359),
.B2(n_364),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_377),
.A2(n_324),
.B1(n_345),
.B2(n_342),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_393),
.B1(n_395),
.B2(n_362),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_386),
.Y(n_409)
);

AOI322xp5_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_319),
.A3(n_245),
.B1(n_341),
.B2(n_335),
.C1(n_332),
.C2(n_325),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_384),
.B(n_185),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_339),
.C(n_334),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_387),
.C(n_389),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_325),
.C(n_338),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_235),
.C(n_243),
.Y(n_389)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_392),
.B(n_150),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_361),
.A2(n_245),
.B1(n_204),
.B2(n_205),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_352),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_396),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_352),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_195),
.Y(n_397)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_368),
.A2(n_178),
.B(n_152),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_400),
.A2(n_403),
.B(n_370),
.Y(n_414)
);

INVx13_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_353),
.A2(n_177),
.B(n_212),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_209),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_388),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_210),
.Y(n_405)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_406),
.A2(n_425),
.B1(n_413),
.B2(n_395),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_401),
.A2(n_356),
.B1(n_354),
.B2(n_369),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_407),
.A2(n_411),
.B1(n_413),
.B2(n_417),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_419),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_410),
.A2(n_398),
.B1(n_399),
.B2(n_396),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_401),
.A2(n_356),
.B1(n_354),
.B2(n_369),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_380),
.A2(n_354),
.B1(n_371),
.B2(n_351),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_414),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_415),
.B(n_429),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_380),
.A2(n_370),
.B1(n_358),
.B2(n_362),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_375),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_358),
.C(n_206),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_422),
.Y(n_431)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_421),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_141),
.C(n_155),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_218),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_400),
.Y(n_443)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_428),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_427),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_434),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_408),
.C(n_419),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_385),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_436),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_438),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_440),
.A2(n_378),
.B1(n_184),
.B2(n_199),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_391),
.Y(n_441)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_442),
.A2(n_418),
.B1(n_402),
.B2(n_405),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_411),
.Y(n_452)
);

NAND2x1_ASAP7_75t_SL g444 ( 
.A(n_427),
.B(n_399),
.Y(n_444)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_392),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_447),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_448),
.Y(n_460)
);

FAx1_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_394),
.CI(n_382),
.CON(n_449),
.SN(n_449)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_402),
.B(n_391),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_404),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_393),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_456),
.Y(n_476)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_415),
.Y(n_456)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_432),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_461),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_424),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_422),
.C(n_414),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_463),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_398),
.C(n_403),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_429),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_464),
.B(n_451),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_465),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_468),
.A2(n_199),
.B1(n_162),
.B2(n_268),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_446),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_470),
.A2(n_451),
.B1(n_449),
.B2(n_378),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_437),
.C(n_456),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_471),
.B(n_473),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_467),
.A2(n_439),
.B1(n_430),
.B2(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_431),
.C(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_478),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_483),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_460),
.A2(n_449),
.B1(n_444),
.B2(n_446),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_477),
.B(n_482),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_462),
.C(n_461),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_112),
.C(n_167),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_485),
.Y(n_498)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_268),
.C(n_211),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_1),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_454),
.C(n_466),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_489),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_464),
.C(n_465),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_481),
.A2(n_196),
.B(n_111),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_490),
.A2(n_496),
.B(n_499),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_131),
.C(n_30),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_497),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_478),
.A2(n_131),
.B(n_30),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_473),
.C(n_476),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_479),
.A2(n_30),
.B(n_2),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_501),
.B(n_1),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_504),
.A2(n_506),
.B(n_6),
.Y(n_517)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_505),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_495),
.A2(n_483),
.B(n_487),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_492),
.Y(n_507)
);

AOI21xp33_ASAP7_75t_SL g515 ( 
.A1(n_507),
.A2(n_510),
.B(n_501),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_484),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_509),
.B(n_491),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_2),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_5),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_5),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_514),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_SL g519 ( 
.A1(n_515),
.A2(n_508),
.B(n_8),
.C(n_9),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_502),
.A2(n_12),
.B(n_7),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_7),
.C(n_8),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_503),
.B(n_510),
.Y(n_518)
);

AOI21x1_ASAP7_75t_L g522 ( 
.A1(n_518),
.A2(n_519),
.B(n_521),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_520),
.A2(n_512),
.B(n_9),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_8),
.C(n_10),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_522),
.B(n_11),
.Y(n_525)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_10),
.B(n_11),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_526),
.B(n_11),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_12),
.Y(n_528)
);


endmodule