module real_aes_795_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_0), .B(n_143), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_1), .A2(n_151), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_2), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_3), .B(n_143), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_4), .B(n_170), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_5), .B(n_170), .Y(n_473) );
INVx1_ASAP7_75t_L g139 ( .A(n_6), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_7), .B(n_170), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_8), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g543 ( .A(n_9), .B(n_168), .Y(n_543) );
AND2x2_ASAP7_75t_L g173 ( .A(n_10), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g184 ( .A(n_11), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g130 ( .A(n_12), .Y(n_130) );
AOI221x1_ASAP7_75t_L g448 ( .A1(n_13), .A2(n_25), .B1(n_143), .B2(n_151), .C(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_14), .B(n_170), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_16), .B(n_143), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_17), .A2(n_85), .B1(n_103), .B2(n_104), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_17), .Y(n_103) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_18), .A2(n_185), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_19), .B(n_128), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_20), .B(n_170), .Y(n_526) );
AO21x1_ASAP7_75t_L g468 ( .A1(n_21), .A2(n_143), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_22), .B(n_143), .Y(n_224) );
INVx1_ASAP7_75t_L g114 ( .A(n_23), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_24), .A2(n_89), .B1(n_134), .B2(n_143), .Y(n_133) );
NAND2x1_ASAP7_75t_L g460 ( .A(n_26), .B(n_170), .Y(n_460) );
NAND2x1_ASAP7_75t_L g501 ( .A(n_27), .B(n_168), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_28), .Y(n_752) );
OR2x2_ASAP7_75t_L g131 ( .A(n_29), .B(n_86), .Y(n_131) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_29), .A2(n_86), .B(n_130), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_30), .B(n_168), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_31), .B(n_170), .Y(n_542) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_32), .A2(n_174), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_33), .B(n_168), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_34), .A2(n_151), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_35), .B(n_170), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_36), .A2(n_151), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g141 ( .A(n_37), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g149 ( .A(n_37), .B(n_139), .Y(n_149) );
INVx1_ASAP7_75t_L g155 ( .A(n_37), .Y(n_155) );
OR2x6_ASAP7_75t_L g112 ( .A(n_38), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_39), .B(n_143), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_40), .B(n_143), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_41), .B(n_170), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_42), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_43), .B(n_168), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_44), .B(n_143), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_45), .A2(n_151), .B(n_166), .Y(n_165) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_46), .A2(n_101), .B1(n_729), .B2(n_740), .C1(n_753), .C2(n_757), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_46), .A2(n_60), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_46), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_47), .A2(n_151), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_48), .B(n_168), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_49), .A2(n_102), .B1(n_722), .B2(n_726), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_50), .B(n_168), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_51), .B(n_143), .Y(n_236) );
INVx1_ASAP7_75t_L g137 ( .A(n_52), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_52), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_53), .B(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g204 ( .A(n_54), .B(n_128), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_55), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_56), .B(n_170), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_57), .B(n_168), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_58), .A2(n_151), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_59), .B(n_143), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_60), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_61), .B(n_143), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_62), .A2(n_151), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g230 ( .A(n_63), .B(n_129), .Y(n_230) );
AO21x1_ASAP7_75t_L g470 ( .A1(n_64), .A2(n_151), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_65), .B(n_143), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_66), .B(n_168), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_67), .B(n_143), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_68), .B(n_168), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_69), .A2(n_93), .B1(n_151), .B2(n_153), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_70), .B(n_170), .Y(n_227) );
AND2x2_ASAP7_75t_L g484 ( .A(n_71), .B(n_129), .Y(n_484) );
INVx1_ASAP7_75t_L g142 ( .A(n_72), .Y(n_142) );
INVx1_ASAP7_75t_L g148 ( .A(n_72), .Y(n_148) );
AND2x2_ASAP7_75t_L g504 ( .A(n_73), .B(n_174), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_74), .B(n_168), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_75), .A2(n_151), .B(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_76), .A2(n_151), .B(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_77), .A2(n_151), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g221 ( .A(n_78), .B(n_129), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_79), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
AND2x2_ASAP7_75t_L g489 ( .A(n_81), .B(n_174), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_82), .B(n_143), .Y(n_528) );
AND2x2_ASAP7_75t_L g197 ( .A(n_83), .B(n_185), .Y(n_197) );
AND2x2_ASAP7_75t_L g469 ( .A(n_84), .B(n_211), .Y(n_469) );
INVx1_ASAP7_75t_L g104 ( .A(n_85), .Y(n_104) );
AND2x2_ASAP7_75t_L g463 ( .A(n_87), .B(n_174), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_88), .B(n_168), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_90), .B(n_170), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_91), .B(n_168), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_92), .A2(n_151), .B(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_94), .A2(n_151), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_95), .B(n_170), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_96), .B(n_170), .Y(n_494) );
BUFx2_ASAP7_75t_L g229 ( .A(n_97), .Y(n_229) );
BUFx2_ASAP7_75t_L g737 ( .A(n_98), .Y(n_737) );
BUFx2_ASAP7_75t_SL g761 ( .A(n_98), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_99), .A2(n_151), .B(n_541), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_105), .B(n_721), .Y(n_101) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_116), .B1(n_436), .B2(n_440), .Y(n_106) );
CKINVDCx11_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx6p67_ASAP7_75t_R g723 ( .A(n_108), .Y(n_723) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AND2x6_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x6_ASAP7_75t_SL g438 ( .A(n_111), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g728 ( .A(n_111), .B(n_112), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_111), .B(n_439), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_112), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_116), .A2(n_117), .B1(n_743), .B2(n_746), .Y(n_742) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_117), .A2(n_441), .B1(n_723), .B2(n_724), .Y(n_722) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_373), .Y(n_117) );
NAND3xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_289), .C(n_326), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_257), .C(n_272), .Y(n_119) );
OAI221xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_201), .B1(n_231), .B2(n_243), .C(n_244), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_123), .B(n_186), .Y(n_122) );
OAI22xp33_ASAP7_75t_SL g317 ( .A1(n_123), .A2(n_281), .B1(n_318), .B2(n_321), .Y(n_317) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_158), .Y(n_123) );
OAI21xp33_ASAP7_75t_SL g327 ( .A1(n_124), .A2(n_328), .B(n_334), .Y(n_327) );
OR2x2_ASAP7_75t_L g356 ( .A(n_124), .B(n_188), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_124), .B(n_276), .Y(n_357) );
INVx2_ASAP7_75t_L g388 ( .A(n_124), .Y(n_388) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_125), .B(n_248), .Y(n_369) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g243 ( .A(n_126), .B(n_161), .Y(n_243) );
BUFx3_ASAP7_75t_L g269 ( .A(n_126), .Y(n_269) );
AND2x2_ASAP7_75t_L g405 ( .A(n_126), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g428 ( .A(n_126), .B(n_189), .Y(n_428) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
AND2x4_ASAP7_75t_L g200 ( .A(n_127), .B(n_132), .Y(n_200) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_128), .A2(n_133), .B(n_150), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_128), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_128), .A2(n_192), .B(n_193), .Y(n_191) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_128), .A2(n_448), .B(n_452), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_128), .A2(n_491), .B(n_492), .Y(n_490) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_128), .A2(n_448), .B(n_452), .Y(n_591) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x4_ASAP7_75t_L g211 ( .A(n_130), .B(n_131), .Y(n_211) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g152 ( .A(n_137), .B(n_139), .Y(n_152) );
AND2x4_ASAP7_75t_L g170 ( .A(n_137), .B(n_147), .Y(n_170) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g151 ( .A(n_141), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
AND2x6_ASAP7_75t_L g168 ( .A(n_142), .B(n_145), .Y(n_168) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
AND2x4_ASAP7_75t_L g153 ( .A(n_152), .B(n_154), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_159), .B(n_189), .Y(n_348) );
INVx1_ASAP7_75t_L g385 ( .A(n_159), .Y(n_385) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_175), .Y(n_159) );
AND2x2_ASAP7_75t_L g199 ( .A(n_160), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g406 ( .A(n_160), .Y(n_406) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g249 ( .A(n_161), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_161), .B(n_175), .Y(n_250) );
AND2x2_ASAP7_75t_L g271 ( .A(n_161), .B(n_190), .Y(n_271) );
AND2x2_ASAP7_75t_L g353 ( .A(n_161), .B(n_176), .Y(n_353) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_173), .Y(n_161) );
INVx4_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_172), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_168), .B(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_171), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_171), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_171), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_171), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_171), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_171), .A2(n_239), .B(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_171), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_171), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_171), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_171), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_171), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_171), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_171), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_171), .A2(n_542), .B(n_543), .Y(n_541) );
INVx3_ASAP7_75t_L g214 ( .A(n_174), .Y(n_214) );
AND2x4_ASAP7_75t_SL g246 ( .A(n_175), .B(n_190), .Y(n_246) );
INVx1_ASAP7_75t_L g277 ( .A(n_175), .Y(n_277) );
INVx2_ASAP7_75t_L g285 ( .A(n_175), .Y(n_285) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_175), .Y(n_309) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_176), .Y(n_198) );
AOI21x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_184), .Y(n_176) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_177), .A2(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_183), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_185), .A2(n_224), .B(n_225), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_199), .Y(n_186) );
AND2x2_ASAP7_75t_L g424 ( .A(n_187), .B(n_287), .Y(n_424) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_189), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g335 ( .A(n_189), .B(n_250), .Y(n_335) );
AND2x2_ASAP7_75t_L g352 ( .A(n_189), .B(n_353), .Y(n_352) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x4_ASAP7_75t_L g276 ( .A(n_190), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g292 ( .A(n_190), .Y(n_292) );
AND2x2_ASAP7_75t_L g336 ( .A(n_190), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g343 ( .A(n_190), .B(n_344), .Y(n_343) );
NOR2x1_ASAP7_75t_L g358 ( .A(n_190), .B(n_249), .Y(n_358) );
BUFx2_ASAP7_75t_L g368 ( .A(n_190), .Y(n_368) );
AND2x2_ASAP7_75t_L g393 ( .A(n_190), .B(n_353), .Y(n_393) );
AND2x2_ASAP7_75t_L g414 ( .A(n_190), .B(n_415), .Y(n_414) );
OR2x6_ASAP7_75t_L g190 ( .A(n_191), .B(n_197), .Y(n_190) );
INVx1_ASAP7_75t_L g345 ( .A(n_198), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_199), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g375 ( .A(n_199), .B(n_246), .Y(n_375) );
INVx3_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
AND2x2_ASAP7_75t_L g415 ( .A(n_200), .B(n_337), .Y(n_415) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_202), .A2(n_245), .B1(n_250), .B2(n_251), .Y(n_244) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_212), .Y(n_202) );
INVx4_ASAP7_75t_L g242 ( .A(n_203), .Y(n_242) );
INVx2_ASAP7_75t_L g279 ( .A(n_203), .Y(n_279) );
NAND2x1_ASAP7_75t_L g305 ( .A(n_203), .B(n_222), .Y(n_305) );
OR2x2_ASAP7_75t_L g320 ( .A(n_203), .B(n_255), .Y(n_320) );
OR2x2_ASAP7_75t_SL g347 ( .A(n_203), .B(n_319), .Y(n_347) );
AND2x2_ASAP7_75t_L g360 ( .A(n_203), .B(n_234), .Y(n_360) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_203), .Y(n_381) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_211), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_211), .A2(n_236), .B(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_211), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g522 ( .A(n_211), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_211), .A2(n_539), .B(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g260 ( .A(n_212), .Y(n_260) );
AND2x2_ASAP7_75t_L g392 ( .A(n_212), .B(n_366), .Y(n_392) );
NOR2x1_ASAP7_75t_SL g212 ( .A(n_213), .B(n_222), .Y(n_212) );
AND2x2_ASAP7_75t_L g233 ( .A(n_213), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g409 ( .A(n_213), .B(n_332), .Y(n_409) );
AO21x1_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_213) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_256) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_214), .A2(n_457), .B(n_463), .Y(n_456) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_214), .A2(n_478), .B(n_484), .Y(n_477) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_214), .A2(n_478), .B(n_484), .Y(n_511) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_214), .A2(n_457), .B(n_463), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
OR2x2_ASAP7_75t_L g241 ( .A(n_222), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g252 ( .A(n_222), .B(n_242), .Y(n_252) );
AND2x2_ASAP7_75t_L g298 ( .A(n_222), .B(n_255), .Y(n_298) );
OR2x2_ASAP7_75t_L g319 ( .A(n_222), .B(n_234), .Y(n_319) );
INVx2_ASAP7_75t_SL g325 ( .A(n_222), .Y(n_325) );
AND2x2_ASAP7_75t_L g331 ( .A(n_222), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g341 ( .A(n_222), .B(n_324), .Y(n_341) );
BUFx2_ASAP7_75t_L g363 ( .A(n_222), .Y(n_363) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_230), .Y(n_222) );
INVx2_ASAP7_75t_L g410 ( .A(n_231), .Y(n_410) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_241), .Y(n_231) );
OR2x2_ASAP7_75t_L g435 ( .A(n_232), .B(n_279), .Y(n_435) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_233), .B(n_242), .Y(n_301) );
AND2x2_ASAP7_75t_L g372 ( .A(n_233), .B(n_252), .Y(n_372) );
INVx1_ASAP7_75t_L g254 ( .A(n_234), .Y(n_254) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
INVx1_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
INVx2_ASAP7_75t_L g332 ( .A(n_234), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g262 ( .A(n_242), .B(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g322 ( .A(n_242), .Y(n_322) );
INVx2_ASAP7_75t_SL g398 ( .A(n_243), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_245), .A2(n_300), .B1(n_302), .B2(n_306), .Y(n_299) );
AND2x2_ASAP7_75t_SL g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g426 ( .A(n_246), .B(n_282), .Y(n_426) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_248), .B(n_292), .Y(n_371) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g337 ( .A(n_249), .B(n_285), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_250), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g280 ( .A(n_251), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_251), .A2(n_395), .B1(n_399), .B2(n_401), .C(n_403), .Y(n_394) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g264 ( .A(n_252), .B(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_252), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_252), .B(n_295), .Y(n_350) );
INVx1_ASAP7_75t_SL g346 ( .A(n_253), .Y(n_346) );
AOI221xp5_ASAP7_75t_SL g374 ( .A1(n_253), .A2(n_264), .B1(n_375), .B2(n_376), .C(n_379), .Y(n_374) );
AOI322xp5_ASAP7_75t_L g407 ( .A1(n_253), .A2(n_325), .A3(n_352), .B1(n_408), .B2(n_410), .C1(n_411), .C2(n_414), .Y(n_407) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
BUFx2_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_255), .Y(n_266) );
INVx2_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
AND2x2_ASAP7_75t_L g365 ( .A(n_255), .B(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OA21x2_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_264), .B(n_267), .Y(n_257) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_258), .A2(n_428), .B(n_429), .C(n_433), .Y(n_427) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OR2x2_ASAP7_75t_L g316 ( .A(n_260), .B(n_278), .Y(n_316) );
OR2x2_ASAP7_75t_L g400 ( .A(n_260), .B(n_295), .Y(n_400) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g340 ( .A(n_262), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g418 ( .A(n_265), .Y(n_418) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OR2x2_ASAP7_75t_L g273 ( .A(n_269), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g308 ( .A(n_271), .B(n_309), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .A3(n_278), .B1(n_280), .B2(n_281), .C1(n_286), .C2(n_288), .Y(n_272) );
INVx1_ASAP7_75t_L g314 ( .A(n_273), .Y(n_314) );
OR2x2_ASAP7_75t_L g286 ( .A(n_275), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_275), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g297 ( .A(n_279), .B(n_298), .Y(n_297) );
OAI32xp33_ASAP7_75t_L g342 ( .A1(n_279), .A2(n_343), .A3(n_346), .B1(n_347), .B2(n_348), .Y(n_342) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g287 ( .A(n_282), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_282), .B(n_345), .Y(n_344) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_282), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g408 ( .A(n_282), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g329 ( .A(n_283), .Y(n_329) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_287), .B(n_353), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_310), .Y(n_289) );
OAI21xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .B(n_299), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_SL g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g359 ( .A(n_298), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_301), .A2(n_321), .B1(n_423), .B2(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_303), .A2(n_350), .B(n_351), .C(n_354), .Y(n_349) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx3_ASAP7_75t_L g431 ( .A(n_305), .Y(n_431) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g312 ( .A(n_309), .Y(n_312) );
AO21x1_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B(n_317), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g377 ( .A(n_312), .Y(n_377) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_318), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g333 ( .A(n_320), .Y(n_333) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g390 ( .A(n_323), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NOR3xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_349), .C(n_361), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
OAI21xp5_ASAP7_75t_SL g391 ( .A1(n_330), .A2(n_392), .B(n_393), .Y(n_391) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
O2A1O1Ixp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_336), .B(n_338), .C(n_342), .Y(n_334) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_344), .Y(n_434) );
INVx2_ASAP7_75t_L g419 ( .A(n_347), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_348), .A2(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g413 ( .A(n_353), .Y(n_413) );
OAI31xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .A3(n_358), .B(n_359), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g432 ( .A(n_360), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_367), .B(n_370), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
BUFx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g382 ( .A(n_365), .Y(n_382) );
AOI21xp33_ASAP7_75t_SL g429 ( .A1(n_367), .A2(n_430), .B(n_432), .Y(n_429) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_368), .B(n_388), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_368), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g378 ( .A(n_369), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND5xp2_ASAP7_75t_L g373 ( .A(n_374), .B(n_394), .C(n_407), .D(n_416), .E(n_427), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_386), .B2(n_389), .C(n_391), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_422), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_437), .Y(n_725) );
CKINVDCx11_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND4xp75_ASAP7_75t_L g441 ( .A(n_442), .B(n_631), .C(n_671), .D(n_700), .Y(n_441) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_593), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_550), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_485), .B(n_505), .Y(n_444) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_453), .Y(n_445) );
AND2x4_ASAP7_75t_L g549 ( .A(n_446), .B(n_510), .Y(n_549) );
INVx1_ASAP7_75t_SL g602 ( .A(n_446), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g637 ( .A1(n_446), .A2(n_638), .B(n_641), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_SL g641 ( .A1(n_446), .A2(n_642), .B(n_643), .C(n_644), .Y(n_641) );
NAND2x1_ASAP7_75t_L g682 ( .A(n_446), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_446), .B(n_643), .Y(n_704) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_447), .Y(n_581) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_464), .Y(n_453) );
AND2x2_ASAP7_75t_L g573 ( .A(n_454), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g654 ( .A(n_454), .B(n_510), .Y(n_654) );
INVx1_ASAP7_75t_L g714 ( .A(n_454), .Y(n_714) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g558 ( .A(n_455), .B(n_476), .Y(n_558) );
AND2x2_ASAP7_75t_L g683 ( .A(n_455), .B(n_477), .Y(n_683) );
AND2x2_ASAP7_75t_L g688 ( .A(n_455), .B(n_648), .Y(n_688) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp67_ASAP7_75t_L g564 ( .A(n_456), .Y(n_564) );
BUFx3_ASAP7_75t_L g597 ( .A(n_456), .Y(n_597) );
AND2x2_ASAP7_75t_L g643 ( .A(n_456), .B(n_477), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .Y(n_457) );
AND2x2_ASAP7_75t_L g628 ( .A(n_464), .B(n_507), .Y(n_628) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .Y(n_464) );
AND2x4_ASAP7_75t_L g510 ( .A(n_465), .B(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g620 ( .A(n_465), .B(n_604), .Y(n_620) );
AND2x2_ASAP7_75t_SL g663 ( .A(n_465), .B(n_591), .Y(n_663) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g599 ( .A(n_466), .Y(n_599) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g560 ( .A(n_467), .Y(n_560) );
OAI21x1_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_470), .B(n_474), .Y(n_467) );
INVx1_ASAP7_75t_L g475 ( .A(n_469), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_476), .B(n_560), .Y(n_563) );
AND2x2_ASAP7_75t_L g648 ( .A(n_476), .B(n_591), .Y(n_648) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g645 ( .A(n_477), .B(n_508), .Y(n_645) );
AND2x2_ASAP7_75t_L g665 ( .A(n_477), .B(n_591), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_483), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_485), .B(n_554), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_485), .A2(n_677), .B1(n_678), .B2(n_679), .C(n_681), .Y(n_676) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI332xp33_ASAP7_75t_L g710 ( .A1(n_486), .A2(n_570), .A3(n_577), .B1(n_636), .B2(n_711), .B3(n_712), .C1(n_713), .C2(n_715), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
AND2x2_ASAP7_75t_L g516 ( .A(n_487), .B(n_497), .Y(n_516) );
AND2x2_ASAP7_75t_L g533 ( .A(n_487), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g545 ( .A(n_487), .Y(n_545) );
AND2x2_ASAP7_75t_SL g605 ( .A(n_487), .B(n_546), .Y(n_605) );
INVx5_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2x1_ASAP7_75t_SL g567 ( .A(n_488), .B(n_534), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_488), .B(n_496), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_488), .B(n_497), .Y(n_578) );
BUFx2_ASAP7_75t_L g613 ( .A(n_488), .Y(n_613) );
AND2x2_ASAP7_75t_L g668 ( .A(n_488), .B(n_537), .Y(n_668) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OR2x2_ASAP7_75t_L g536 ( .A(n_496), .B(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g546 ( .A(n_496), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g586 ( .A(n_496), .Y(n_586) );
AND2x2_ASAP7_75t_L g656 ( .A(n_496), .B(n_555), .Y(n_656) );
AND2x2_ASAP7_75t_L g669 ( .A(n_496), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_496), .B(n_670), .Y(n_687) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_497), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
OAI32xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_512), .A3(n_517), .B1(n_531), .B2(n_548), .Y(n_505) );
INVx2_ASAP7_75t_L g614 ( .A(n_506), .Y(n_614) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g625 ( .A(n_507), .Y(n_625) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g559 ( .A(n_508), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g692 ( .A(n_508), .B(n_597), .Y(n_692) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g604 ( .A(n_511), .Y(n_604) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g592 ( .A(n_514), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_514), .B(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_SL g603 ( .A(n_515), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g680 ( .A(n_515), .Y(n_680) );
AND2x2_ASAP7_75t_L g698 ( .A(n_515), .B(n_560), .Y(n_698) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2xp67_ASAP7_75t_SL g642 ( .A(n_518), .B(n_571), .Y(n_642) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_519), .B(n_553), .Y(n_640) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g716 ( .A(n_520), .B(n_586), .Y(n_716) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g547 ( .A(n_521), .Y(n_547) );
INVx2_ASAP7_75t_L g588 ( .A(n_521), .Y(n_588) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_529), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_522), .B(n_530), .Y(n_529) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_522), .A2(n_523), .B(n_529), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_528), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_544), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_532), .B(n_590), .Y(n_675) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND3x2_ASAP7_75t_L g630 ( .A(n_533), .B(n_577), .C(n_586), .Y(n_630) );
AND2x2_ASAP7_75t_L g554 ( .A(n_534), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_534), .B(n_537), .Y(n_611) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g565 ( .A(n_536), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g555 ( .A(n_537), .Y(n_555) );
INVx1_ASAP7_75t_L g570 ( .A(n_537), .Y(n_570) );
BUFx3_ASAP7_75t_L g577 ( .A(n_537), .Y(n_577) );
AND2x2_ASAP7_75t_L g587 ( .A(n_537), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AND2x4_ASAP7_75t_L g596 ( .A(n_545), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_545), .B(n_555), .Y(n_639) );
AND2x2_ASAP7_75t_L g595 ( .A(n_546), .B(n_570), .Y(n_595) );
INVx2_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_556), .B(n_561), .C(n_582), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_551), .A2(n_678), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_554), .B(n_613), .Y(n_612) );
AOI211xp5_ASAP7_75t_SL g632 ( .A1(n_554), .A2(n_633), .B(n_637), .C(n_646), .Y(n_632) );
AND2x2_ASAP7_75t_L g618 ( .A(n_555), .B(n_578), .Y(n_618) );
OR2x2_ASAP7_75t_L g621 ( .A(n_555), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_558), .B(n_663), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_559), .B(n_604), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_559), .A2(n_585), .B1(n_665), .B2(n_668), .C(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g590 ( .A(n_560), .B(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g636 ( .A(n_560), .B(n_591), .Y(n_636) );
OAI221xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_565), .B1(n_568), .B2(n_572), .C(n_575), .Y(n_561) );
AND2x2_ASAP7_75t_L g707 ( .A(n_562), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g574 ( .A(n_563), .Y(n_574) );
INVx1_ASAP7_75t_L g660 ( .A(n_564), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_565), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g579 ( .A(n_567), .B(n_570), .Y(n_579) );
AND2x2_ASAP7_75t_L g655 ( .A(n_567), .B(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g580 ( .A(n_574), .B(n_581), .Y(n_580) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_579), .B(n_580), .Y(n_575) );
INVx1_ASAP7_75t_L g699 ( .A(n_576), .Y(n_699) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g678 ( .A(n_577), .B(n_605), .Y(n_678) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_578), .B(n_587), .Y(n_651) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_589), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_583), .A2(n_617), .B1(n_620), .B2(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g689 ( .A(n_583), .Y(n_689) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g609 ( .A(n_586), .Y(n_609) );
INVx1_ASAP7_75t_L g670 ( .A(n_588), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_590), .B(n_660), .Y(n_711) );
AND2x2_ASAP7_75t_L g679 ( .A(n_591), .B(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g672 ( .A1(n_592), .A2(n_673), .B(n_676), .C(n_684), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_615), .Y(n_593) );
AOI322xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .A3(n_598), .B1(n_600), .B2(n_605), .C1(n_606), .C2(n_614), .Y(n_594) );
CKINVDCx16_ASAP7_75t_R g712 ( .A(n_596), .Y(n_712) );
AND2x2_ASAP7_75t_L g662 ( .A(n_597), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g696 ( .A(n_597), .Y(n_696) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_SL g647 ( .A(n_599), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_599), .B(n_645), .Y(n_653) );
AND2x2_ASAP7_75t_L g677 ( .A(n_599), .B(n_643), .Y(n_677) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g649 ( .A(n_603), .Y(n_649) );
NAND2xp33_ASAP7_75t_SL g606 ( .A(n_607), .B(n_612), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI221xp5_ASAP7_75t_SL g652 ( .A1(n_608), .A2(n_653), .B1(n_654), .B2(n_655), .C(n_657), .Y(n_652) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g719 ( .A(n_611), .Y(n_719) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_619), .C(n_623), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g694 ( .A(n_618), .Y(n_694) );
INVx1_ASAP7_75t_L g626 ( .A(n_620), .Y(n_626) );
OR2x2_ASAP7_75t_L g713 ( .A(n_620), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g709 ( .A(n_621), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_629), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_625), .B(n_643), .Y(n_720) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_652), .Y(n_631) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_635), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g686 ( .A(n_639), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_649), .B(n_650), .Y(n_646) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AOI31xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .A3(n_664), .B(n_666), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_663), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B1(n_689), .B2(n_690), .C(n_693), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_697), .B2(n_699), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g697 ( .A(n_698), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_710), .C(n_717), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx4f_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_738), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_734), .B(n_737), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_SL g756 ( .A(n_735), .B(n_737), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_735), .A2(n_759), .B(n_762), .Y(n_758) );
INVx1_ASAP7_75t_SL g748 ( .A(n_738), .Y(n_748) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx3_ASAP7_75t_L g751 ( .A(n_739), .Y(n_751) );
BUFx2_ASAP7_75t_L g763 ( .A(n_739), .Y(n_763) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_747), .B(n_749), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_743), .Y(n_746) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_SL g749 ( .A(n_750), .B(n_752), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
CKINVDCx11_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
CKINVDCx8_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule