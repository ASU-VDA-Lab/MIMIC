module fake_jpeg_19646_n_285 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_93;
wire n_54;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_24),
.C(n_20),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_37),
.B1(n_29),
.B2(n_22),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_60),
.Y(n_69)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_19),
.B1(n_34),
.B2(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_27),
.B1(n_15),
.B2(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_66),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_63),
.A2(n_86),
.B(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_36),
.B1(n_37),
.B2(n_21),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_43),
.A3(n_41),
.B1(n_21),
.B2(n_22),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_74),
.A3(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_41),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_77),
.B1(n_89),
.B2(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_54),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_37),
.B1(n_22),
.B2(n_35),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_39),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_39),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_21),
.B(n_30),
.C(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_27),
.B1(n_35),
.B2(n_30),
.Y(n_86)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_26),
.B1(n_34),
.B2(n_39),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_27),
.B1(n_35),
.B2(n_25),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_42),
.B1(n_38),
.B2(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_48),
.A2(n_42),
.B(n_38),
.C(n_44),
.Y(n_96)
);

AND2x4_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_25),
.B1(n_23),
.B2(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_63),
.C(n_62),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_107),
.C(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_54),
.C(n_48),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_32),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_73),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_151),
.B(n_119),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_97),
.B1(n_66),
.B2(n_92),
.Y(n_129)
);

OAI22x1_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_151),
.B1(n_133),
.B2(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_141),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_104),
.B(n_123),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_138),
.B(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_81),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_72),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_71),
.B(n_69),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_84),
.C(n_82),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_145),
.C(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_69),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_124),
.B(n_74),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_115),
.B1(n_120),
.B2(n_104),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_148),
.B1(n_149),
.B2(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_77),
.C(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_65),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_115),
.B1(n_110),
.B2(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_110),
.A2(n_91),
.B1(n_83),
.B2(n_96),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_76),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_152),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_96),
.B1(n_97),
.B2(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_28),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_117),
.B1(n_114),
.B2(n_116),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_93),
.C(n_54),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_161),
.B(n_162),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2x1p5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_42),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_175),
.C(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_99),
.B1(n_78),
.B2(n_100),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_179),
.B1(n_181),
.B2(n_131),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_105),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_180),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_42),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_182),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_125),
.C(n_54),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_177),
.C(n_176),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_78),
.B1(n_85),
.B2(n_38),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_44),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_31),
.B1(n_33),
.B2(n_32),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_32),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_193),
.B(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_197),
.C(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_167),
.A2(n_145),
.B1(n_148),
.B2(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_188),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_151),
.B1(n_128),
.B2(n_150),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_196),
.Y(n_218)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_175),
.B1(n_183),
.B2(n_180),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_152),
.B(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_142),
.C(n_109),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_163),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_109),
.C(n_44),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_20),
.C(n_31),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_179),
.C(n_173),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_23),
.B(n_25),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_11),
.B1(n_16),
.B2(n_2),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_204),
.A2(n_155),
.B1(n_174),
.B2(n_166),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_207),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_214),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_156),
.B1(n_155),
.B2(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_159),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_220),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_87),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_172),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_170),
.C(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_223),
.C(n_20),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_159),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_224),
.B1(n_184),
.B2(n_20),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_170),
.C(n_20),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_87),
.B(n_1),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_233),
.B1(n_23),
.B2(n_33),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_193),
.C(n_201),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_229),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_194),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_201),
.B(n_203),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_230),
.A2(n_232),
.B(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_199),
.C(n_187),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.C(n_238),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_192),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_190),
.B1(n_205),
.B2(n_184),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_200),
.C(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_33),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_241),
.C(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_209),
.B1(n_224),
.B2(n_222),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_251),
.B1(n_255),
.B2(n_5),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_219),
.B(n_223),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_249),
.C(n_253),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_250),
.B1(n_3),
.B2(n_4),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_242),
.B1(n_233),
.B2(n_237),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_238),
.A2(n_6),
.B1(n_15),
.B2(n_2),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_8),
.C(n_15),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_6),
.B1(n_13),
.B2(n_3),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_234),
.C(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_259),
.Y(n_270)
);

FAx1_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_241),
.CI(n_228),
.CON(n_258),
.SN(n_258)
);

AOI31xp33_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_263),
.A3(n_248),
.B(n_250),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_235),
.C(n_10),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_262),
.B1(n_249),
.B2(n_12),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_254),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_264),
.A2(n_245),
.B(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_266),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_263),
.A2(n_252),
.B(n_253),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_269),
.B1(n_271),
.B2(n_258),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_260),
.A2(n_252),
.B(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_257),
.C(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_257),
.B(n_275),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_3),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_279),
.A3(n_4),
.B1(n_12),
.B2(n_13),
.C1(n_16),
.C2(n_1),
.Y(n_283)
);

OAI321xp33_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_0),
.A3(n_1),
.B1(n_12),
.B2(n_16),
.C(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_0),
.Y(n_285)
);


endmodule