module fake_aes_8396_n_711 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_711);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_711;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_26), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_57), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_4), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_70), .B(n_68), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_18), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_71), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_9), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_76), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_43), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_20), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_64), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_15), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_10), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_1), .Y(n_94) );
NOR2xp67_ASAP7_75t_L g95 ( .A(n_60), .B(n_59), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_25), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_78), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_69), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_47), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_51), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_10), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_61), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_49), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_52), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_75), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_33), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_65), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_4), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_35), .B(n_11), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_45), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_55), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_34), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_6), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_42), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_62), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_56), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_90), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
BUFx8_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
BUFx8_ASAP7_75t_L g132 ( .A(n_111), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_106), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_115), .A2(n_29), .B(n_74), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_99), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_115), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_111), .B(n_3), .Y(n_139) );
CKINVDCx6p67_ASAP7_75t_R g140 ( .A(n_97), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_87), .B(n_5), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_124), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_79), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_85), .B(n_6), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_92), .B(n_31), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_79), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_81), .Y(n_155) );
INVx5_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx4_ASAP7_75t_L g160 ( .A(n_103), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_100), .B(n_7), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_123), .A2(n_32), .B(n_72), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_108), .B(n_7), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_104), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_89), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_107), .B(n_8), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_81), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_89), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_93), .B(n_8), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_129), .A2(n_93), .B1(n_120), .B2(n_81), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_148), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_149), .B(n_114), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_129), .A2(n_81), .B1(n_105), .B2(n_80), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_154), .B(n_103), .Y(n_177) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_154), .B(n_126), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_147), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx6f_ASAP7_75t_SL g186 ( .A(n_152), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_131), .B(n_118), .Y(n_187) );
AND3x1_ASAP7_75t_L g188 ( .A(n_136), .B(n_113), .C(n_121), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_128), .B(n_126), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_128), .B(n_127), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_139), .B(n_101), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_139), .B(n_81), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_140), .B(n_125), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_155), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_166), .B(n_125), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_131), .A2(n_102), .B1(n_117), .B2(n_84), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_137), .B(n_110), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_148), .B(n_119), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_137), .B(n_119), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_143), .B(n_96), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_143), .B(n_112), .Y(n_206) );
BUFx4f_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_146), .B(n_109), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_156), .Y(n_211) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_171), .B(n_98), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_130), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_135), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_146), .B(n_86), .Y(n_216) );
INVx6_ASAP7_75t_L g217 ( .A(n_156), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_151), .B(n_95), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
AND2x6_ASAP7_75t_L g220 ( .A(n_165), .B(n_82), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_155), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_135), .Y(n_222) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_144), .B(n_9), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_151), .B(n_113), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_130), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_130), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_133), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_132), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_157), .A2(n_12), .B1(n_13), .B2(n_77), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_157), .B(n_13), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_158), .B(n_14), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_158), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_169), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_159), .B(n_67), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_196), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_233), .B(n_163), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_178), .A2(n_159), .B1(n_163), .B2(n_138), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_226), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_204), .B(n_132), .Y(n_243) );
AND2x6_ASAP7_75t_L g244 ( .A(n_189), .B(n_142), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_190), .B(n_132), .Y(n_245) );
AO22x1_ASAP7_75t_L g246 ( .A1(n_229), .A2(n_150), .B1(n_168), .B2(n_161), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_228), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_200), .B(n_164), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_177), .B(n_164), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_180), .B(n_156), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_202), .B(n_156), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_231), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_215), .B(n_141), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_227), .B(n_141), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_214), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_193), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_202), .B(n_156), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_224), .B(n_156), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
NOR2x1p5_ASAP7_75t_L g262 ( .A(n_229), .B(n_142), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_235), .B(n_138), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g265 ( .A(n_207), .B(n_134), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_187), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_207), .B(n_134), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_176), .B(n_133), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_178), .A2(n_169), .B(n_162), .C(n_22), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_181), .B(n_162), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_181), .B(n_184), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_184), .B(n_162), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_185), .B(n_162), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_185), .B(n_169), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_187), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_217), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_179), .B(n_169), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_226), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_179), .B(n_169), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_212), .B(n_17), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_192), .B(n_21), .Y(n_282) );
AND2x6_ASAP7_75t_SL g283 ( .A(n_174), .B(n_188), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_212), .A2(n_23), .B1(n_24), .B2(n_27), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_186), .A2(n_28), .B1(n_30), .B2(n_36), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_203), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_198), .B(n_38), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_193), .B(n_39), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_205), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_206), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_193), .B(n_44), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_225), .B(n_46), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_210), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_216), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_182), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_236), .B(n_174), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_174), .B(n_48), .Y(n_297) );
OAI22xp5_ASAP7_75t_SL g298 ( .A1(n_223), .A2(n_54), .B1(n_58), .B2(n_63), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_218), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_213), .B(n_66), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_223), .B(n_208), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_201), .B(n_191), .Y(n_302) );
NOR2xp33_ASAP7_75t_SL g303 ( .A(n_186), .B(n_193), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_193), .A2(n_195), .B1(n_220), .B2(n_208), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_195), .B(n_201), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_270), .A2(n_214), .B(n_222), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_257), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_272), .A2(n_214), .B(n_222), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_289), .B(n_195), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_275), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_237), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_264), .B(n_191), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_247), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_264), .B(n_191), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_273), .A2(n_214), .B(n_222), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_286), .A2(n_195), .B1(n_220), .B2(n_230), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_238), .B(n_194), .Y(n_319) );
OAI22x1_ASAP7_75t_L g320 ( .A1(n_241), .A2(n_195), .B1(n_232), .B2(n_230), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_305), .A2(n_172), .B1(n_175), .B2(n_222), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_244), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_258), .B(n_197), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_254), .B(n_220), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_304), .A2(n_172), .B1(n_175), .B2(n_194), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_245), .B(n_197), .Y(n_326) );
BUFx12f_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_242), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_295), .A2(n_232), .B(n_199), .C(n_209), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_258), .B(n_211), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_250), .A2(n_211), .B(n_199), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_290), .A2(n_217), .B1(n_220), .B2(n_234), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_294), .B(n_220), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_183), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_257), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_253), .A2(n_234), .B(n_209), .C(n_219), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_248), .B(n_183), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_239), .A2(n_219), .B1(n_221), .B2(n_301), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_262), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_303), .A2(n_221), .B1(n_293), .B2(n_301), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_252), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_271), .A2(n_274), .B(n_302), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_239), .A2(n_281), .B1(n_292), .B2(n_299), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_256), .B(n_246), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_244), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_300), .B(n_243), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_244), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_296), .B(n_268), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_257), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_300), .A2(n_297), .B1(n_298), .B2(n_268), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_249), .A2(n_263), .B(n_255), .C(n_267), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_255), .B(n_265), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_297), .B(n_244), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_265), .B(n_282), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_261), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_271), .A2(n_251), .B(n_259), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_266), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_351), .A2(n_276), .B1(n_284), .B2(n_285), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_327), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_344), .A2(n_284), .B1(n_288), .B2(n_291), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_287), .B(n_260), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_318), .A2(n_277), .B1(n_283), .B2(n_278), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_308), .A2(n_280), .B(n_257), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_324), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_307), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_343), .A2(n_269), .B1(n_346), .B2(n_309), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g368 ( .A1(n_326), .A2(n_320), .B(n_333), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_345), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_317), .A2(n_357), .B(n_342), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
NOR2xp33_ASAP7_75t_SL g373 ( .A(n_322), .B(n_347), .Y(n_373) );
CKINVDCx14_ASAP7_75t_R g374 ( .A(n_322), .Y(n_374) );
BUFx8_ASAP7_75t_L g375 ( .A(n_324), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_349), .A2(n_353), .B1(n_354), .B2(n_332), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_352), .A2(n_316), .B(n_314), .C(n_337), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_358), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_348), .B(n_307), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_334), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_SL g381 ( .A1(n_355), .A2(n_336), .B(n_329), .C(n_338), .Y(n_381) );
O2A1O1Ixp5_ASAP7_75t_L g382 ( .A1(n_321), .A2(n_354), .B(n_319), .C(n_325), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_331), .A2(n_340), .B(n_358), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_307), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_315), .Y(n_386) );
O2A1O1Ixp5_ASAP7_75t_L g387 ( .A1(n_323), .A2(n_356), .B(n_330), .C(n_312), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_310), .A2(n_311), .B(n_335), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_313), .B(n_328), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_335), .A2(n_350), .B(n_341), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_335), .A2(n_308), .B(n_306), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_371), .A2(n_350), .B(n_381), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_378), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_380), .B(n_350), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_374), .Y(n_395) );
BUFx8_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_359), .A2(n_376), .B1(n_363), .B2(n_365), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_389), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_386), .A2(n_384), .B1(n_373), .B2(n_369), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_377), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_375), .B(n_374), .Y(n_401) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_375), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_372), .B(n_379), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_369), .B(n_370), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_382), .A2(n_367), .B(n_361), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
AOI21x1_ASAP7_75t_L g407 ( .A1(n_391), .A2(n_383), .B(n_388), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_370), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_369), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_368), .A2(n_361), .B(n_383), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g413 ( .A1(n_379), .A2(n_385), .B1(n_366), .B2(n_387), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_362), .B1(n_390), .B2(n_388), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_381), .A2(n_391), .B(n_364), .Y(n_415) );
BUFx12f_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_364), .A2(n_178), .B1(n_264), .B2(n_380), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_375), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_378), .B(n_324), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_415), .A2(n_405), .B(n_411), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_393), .B(n_419), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_393), .B(n_419), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_398), .B(n_420), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_397), .B(n_400), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_416), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_392), .A2(n_407), .B(n_414), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_416), .Y(n_429) );
OAI21x1_ASAP7_75t_L g430 ( .A1(n_412), .A2(n_403), .B(n_417), .Y(n_430) );
OR2x6_ASAP7_75t_L g431 ( .A(n_413), .B(n_404), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_409), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_404), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_408), .B(n_418), .Y(n_435) );
AO21x2_ASAP7_75t_L g436 ( .A1(n_399), .A2(n_404), .B(n_420), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_420), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_410), .B(n_408), .C(n_406), .Y(n_438) );
OR2x6_ASAP7_75t_L g439 ( .A(n_418), .B(n_401), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_410), .B(n_409), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_395), .B(n_396), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_395), .B(n_396), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_380), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_418), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_416), .Y(n_447) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_415), .A2(n_405), .B(n_411), .Y(n_448) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_415), .A2(n_405), .B(n_411), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_393), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_398), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_415), .A2(n_405), .B(n_411), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_393), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_451), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_422), .B(n_423), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_427), .B(n_455), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_426), .A2(n_441), .B1(n_433), .B2(n_437), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_451), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_456), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_429), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_450), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_456), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_443), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_447), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_423), .B(n_432), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_432), .B(n_434), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_426), .B(n_432), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_434), .B(n_436), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_434), .B(n_436), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_430), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_436), .B(n_421), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_443), .A2(n_433), .A3(n_440), .B(n_441), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_436), .B(n_421), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_421), .B(n_425), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_452), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_435), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_428), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_430), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_421), .B(n_454), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_447), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_448), .B(n_454), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_424), .B(n_427), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_427), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_429), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_429), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_429), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_453), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_440), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_448), .B(n_454), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_457), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_458), .B(n_449), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_464), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_501), .B(n_443), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_458), .B(n_445), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_466), .B(n_446), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_479), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_461), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_483), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_461), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_490), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_499), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_469), .B(n_449), .Y(n_518) );
NOR2xp67_ASAP7_75t_L g519 ( .A(n_501), .B(n_443), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_469), .B(n_449), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_471), .B(n_455), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_490), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_462), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_468), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_472), .B(n_455), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_472), .B(n_455), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_473), .B(n_455), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_473), .B(n_455), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_468), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_462), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_480), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_480), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_478), .B(n_453), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_465), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_478), .B(n_453), .Y(n_536) );
INVx6_ASAP7_75t_L g537 ( .A(n_501), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_492), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_471), .B(n_431), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_466), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_470), .B(n_437), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_492), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_470), .B(n_431), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_476), .B(n_440), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_460), .B(n_446), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_502), .B(n_431), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_485), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_475), .B(n_431), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_475), .B(n_431), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_502), .B(n_439), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_477), .B(n_439), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_467), .B(n_439), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_477), .B(n_439), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_476), .B(n_438), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_467), .B(n_442), .Y(n_557) );
INVxp33_ASAP7_75t_L g558 ( .A(n_459), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_486), .B(n_439), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_506), .B(n_488), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_511), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_545), .A2(n_493), .B1(n_486), .B2(n_444), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_506), .B(n_488), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_556), .A2(n_444), .B(n_438), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_509), .B(n_497), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_514), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_543), .B(n_493), .Y(n_567) );
INVx3_ASAP7_75t_SL g568 ( .A(n_537), .Y(n_568) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_535), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_505), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_532), .B(n_494), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_539), .B(n_459), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_518), .B(n_504), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_518), .B(n_504), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_520), .B(n_525), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_549), .B(n_459), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_520), .B(n_491), .Y(n_577) );
NAND2x1_ASAP7_75t_SL g578 ( .A(n_519), .B(n_459), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_505), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_541), .B(n_491), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_531), .B(n_498), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_541), .B(n_498), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_516), .B(n_495), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_525), .B(n_487), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_522), .B(n_495), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_507), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_542), .B(n_497), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_526), .B(n_484), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_537), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_537), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_515), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_524), .B(n_496), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_526), .B(n_484), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_529), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_537), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_527), .B(n_484), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_523), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_487), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_530), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_542), .B(n_496), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_521), .B(n_463), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_528), .B(n_487), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_528), .B(n_481), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_557), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_533), .B(n_481), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_521), .B(n_463), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_540), .B(n_463), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_540), .B(n_463), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_533), .B(n_481), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_565), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_561), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_575), .B(n_536), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_586), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_560), .B(n_548), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_575), .B(n_560), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_596), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_563), .B(n_536), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_568), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_564), .A2(n_442), .B(n_553), .C(n_555), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_566), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_568), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_562), .A2(n_555), .B1(n_553), .B2(n_550), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_569), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_563), .B(n_550), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_573), .B(n_551), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_573), .B(n_510), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_574), .B(n_552), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_586), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_579), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_574), .B(n_551), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_562), .A2(n_508), .B(n_549), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_577), .B(n_512), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_607), .A2(n_546), .B(n_508), .C(n_559), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_590), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_577), .B(n_544), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_591), .A2(n_508), .B1(n_547), .B2(n_549), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_591), .B(n_499), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_596), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g644 ( .A1(n_589), .A2(n_517), .A3(n_552), .B(n_547), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_580), .B(n_558), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_584), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_588), .B(n_544), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_572), .B(n_554), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_621), .B(n_597), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
XNOR2x1_ASAP7_75t_L g652 ( .A(n_624), .B(n_581), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_642), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_638), .B(n_567), .C(n_571), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_614), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_636), .A2(n_576), .B(n_517), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_631), .B(n_587), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_630), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_619), .A2(n_578), .B(n_585), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_618), .B(n_606), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_633), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_639), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_622), .A2(n_576), .B1(n_602), .B2(n_610), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_642), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_641), .A2(n_576), .B(n_611), .C(n_609), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_618), .B(n_600), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_613), .B(n_595), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_643), .B(n_595), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_616), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_615), .B(n_588), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_623), .A2(n_612), .B1(n_608), .B2(n_594), .C1(n_599), .C2(n_601), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_637), .B(n_606), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_652), .A2(n_645), .B1(n_649), .B2(n_635), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_652), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_651), .A2(n_644), .B(n_593), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_658), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_659), .A2(n_645), .B(n_649), .C(n_625), .Y(n_677) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_650), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_665), .A2(n_617), .B1(n_631), .B2(n_629), .C(n_646), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_663), .A2(n_647), .A3(n_634), .B1(n_583), .B2(n_603), .C1(n_620), .C2(n_627), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_660), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_SL g682 ( .A1(n_654), .A2(n_503), .B(n_616), .C(n_632), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_650), .B(n_647), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_654), .A2(n_635), .B1(n_628), .B2(n_627), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_671), .A2(n_668), .B1(n_653), .B2(n_664), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_SL g686 ( .A1(n_656), .A2(n_503), .B(n_632), .C(n_604), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_680), .A2(n_655), .B1(n_661), .B2(n_662), .C(n_667), .Y(n_687) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_674), .A2(n_669), .B(n_672), .C(n_657), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_678), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_673), .A2(n_660), .B(n_670), .C(n_666), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g691 ( .A1(n_685), .A2(n_670), .B(n_628), .C(n_669), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_677), .A2(n_640), .B(n_620), .C(n_499), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_684), .B(n_640), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g694 ( .A1(n_679), .A2(n_615), .B(n_648), .C(n_634), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_687), .A2(n_688), .B1(n_691), .B2(n_690), .C(n_692), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_694), .B(n_678), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g697 ( .A1(n_689), .A2(n_675), .B(n_682), .C(n_686), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_693), .B(n_683), .C(n_676), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_691), .A2(n_681), .B(n_648), .C(n_582), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_695), .B(n_503), .C(n_534), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_696), .A2(n_538), .B1(n_513), .B2(n_474), .C(n_482), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_698), .A2(n_605), .B1(n_598), .B2(n_600), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_700), .Y(n_703) );
NAND4xp75_ASAP7_75t_L g704 ( .A(n_701), .B(n_697), .C(n_699), .D(n_605), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_704), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_703), .B(n_702), .Y(n_706) );
BUFx2_ASAP7_75t_L g707 ( .A(n_705), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_707), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_706), .B1(n_500), .B2(n_489), .C1(n_482), .C2(n_474), .Y(n_709) );
OR2x6_ASAP7_75t_L g710 ( .A(n_709), .B(n_489), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_710), .A2(n_598), .B1(n_608), .B2(n_612), .Y(n_711) );
endmodule