module fake_jpeg_31232_n_237 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_22),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_35),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_32),
.B1(n_24),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_66),
.B1(n_30),
.B2(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_68),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_24),
.B1(n_35),
.B2(n_29),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_73),
.B1(n_75),
.B2(n_29),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_36),
.B1(n_33),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_25),
.B1(n_39),
.B2(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_40),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_18),
.B1(n_27),
.B2(n_28),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_35),
.B1(n_29),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_44),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_20),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_88),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_20),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_87),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_50),
.B1(n_51),
.B2(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_98),
.B1(n_104),
.B2(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_102),
.B1(n_107),
.B2(n_109),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_23),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_17),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_17),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_38),
.B1(n_45),
.B2(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_106),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_38),
.B1(n_45),
.B2(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_42),
.B1(n_48),
.B2(n_47),
.Y(n_105)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_53),
.A2(n_48),
.B1(n_47),
.B2(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_42),
.B1(n_49),
.B2(n_43),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_0),
.B(n_1),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_1),
.B(n_2),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_49),
.B1(n_47),
.B2(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_65),
.B1(n_47),
.B2(n_5),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_1),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_2),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_79),
.B1(n_99),
.B2(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_79),
.B1(n_82),
.B2(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_97),
.B(n_6),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_150),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_90),
.B(n_96),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_139),
.C(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_107),
.B1(n_109),
.B2(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_126),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_102),
.B1(n_84),
.B2(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_85),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_106),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_106),
.B1(n_78),
.B2(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_143),
.B1(n_120),
.B2(n_111),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_117),
.A3(n_126),
.B1(n_113),
.B2(n_131),
.C1(n_112),
.C2(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_2),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_120),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_106),
.B(n_117),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_150),
.B(n_111),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_119),
.B1(n_130),
.B2(n_100),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_119),
.B1(n_116),
.B2(n_151),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_134),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_148),
.C(n_149),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_184),
.C(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_139),
.B(n_144),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_185),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_183),
.B1(n_160),
.B2(n_161),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_180),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_145),
.B1(n_116),
.B2(n_119),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_110),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_130),
.B(n_124),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_124),
.B(n_103),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_193),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_160),
.C(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_197),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_176),
.B1(n_159),
.B2(n_177),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_168),
.C(n_158),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_199),
.C(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_153),
.C(n_158),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_168),
.C(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_205),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_169),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_124),
.B(n_65),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_182),
.B(n_185),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_7),
.B(n_8),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_7),
.C(n_8),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_169),
.B1(n_78),
.B2(n_9),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_169),
.B1(n_198),
.B2(n_188),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_124),
.CI(n_8),
.CON(n_214),
.SN(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_216),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_7),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_204),
.B1(n_200),
.B2(n_209),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_212),
.B1(n_215),
.B2(n_218),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_203),
.C(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_207),
.C(n_9),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_219),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_229),
.B(n_214),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_222),
.B(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_232),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_214),
.C(n_225),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_227),
.C(n_10),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_235),
.A2(n_234),
.B1(n_10),
.B2(n_12),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_9),
.Y(n_237)
);


endmodule