module fake_jpeg_4352_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_17),
.B1(n_32),
.B2(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_7),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_32),
.CON(n_49),
.SN(n_49)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_49),
.B1(n_70),
.B2(n_21),
.Y(n_74)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_24),
.B1(n_25),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_22),
.B1(n_30),
.B2(n_19),
.Y(n_91)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_24),
.B1(n_25),
.B2(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_43),
.B1(n_22),
.B2(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_59),
.Y(n_84)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_26),
.B(n_34),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_34),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_8),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_16),
.B1(n_29),
.B2(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_29),
.B1(n_44),
.B2(n_38),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_65),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_52),
.B1(n_50),
.B2(n_65),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_19),
.B1(n_30),
.B2(n_22),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_31),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_49),
.B1(n_61),
.B2(n_71),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_19),
.B1(n_31),
.B2(n_23),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_105),
.B1(n_120),
.B2(n_84),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_113),
.B(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_107),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_111),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_62),
.C(n_47),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_117),
.CI(n_55),
.CON(n_142),
.SN(n_142)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_69),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_57),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_116),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_48),
.B(n_37),
.C(n_23),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_37),
.B(n_31),
.C(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_55),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_121),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_46),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_27),
.C(n_67),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_131),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_31),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_125),
.A2(n_126),
.B(n_134),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_81),
.B(n_95),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_95),
.B1(n_87),
.B2(n_76),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_129),
.A2(n_104),
.B1(n_133),
.B2(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_78),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_66),
.B1(n_56),
.B2(n_80),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_143),
.B1(n_83),
.B2(n_99),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_86),
.B(n_78),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_86),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_0),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_107),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_87),
.B1(n_80),
.B2(n_56),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_27),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_100),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_141),
.Y(n_195)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_168),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_158),
.B(n_133),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_157),
.B(n_159),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_98),
.Y(n_162)
);

OAI22x1_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_133),
.B1(n_149),
.B2(n_148),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_96),
.B(n_116),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_175),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_96),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_67),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_128),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_187),
.B(n_177),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_138),
.C(n_137),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_146),
.B1(n_149),
.B2(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_125),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_126),
.C(n_125),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_142),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_193),
.C(n_176),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_151),
.C(n_141),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_176),
.C(n_153),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_142),
.C(n_148),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_136),
.B1(n_134),
.B2(n_139),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_211),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_156),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_220),
.B1(n_200),
.B2(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_141),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_226),
.C(n_229),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_221),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_187),
.B(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_166),
.B1(n_159),
.B2(n_139),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_157),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_153),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_172),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_171),
.C(n_152),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_182),
.C(n_179),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_202),
.B1(n_183),
.B2(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_237),
.C(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_180),
.C(n_195),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_218),
.Y(n_253)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_200),
.C(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_196),
.C(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_236),
.C(n_243),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_248),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_160),
.B1(n_167),
.B2(n_152),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_144),
.B1(n_135),
.B2(n_73),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_220),
.A2(n_73),
.B1(n_144),
.B2(n_169),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_248),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_254),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_205),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_216),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_258),
.Y(n_279)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_269),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_211),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_230),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_264),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_265),
.B(n_268),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_214),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_229),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_210),
.C(n_207),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_225),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_272),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_213),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_228),
.B(n_234),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_212),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_278),
.B(n_281),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_233),
.B1(n_246),
.B2(n_247),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_276),
.B1(n_256),
.B2(n_258),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_246),
.B1(n_250),
.B2(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_266),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_286),
.B(n_8),
.Y(n_302)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_245),
.C(n_231),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_15),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_251),
.A3(n_239),
.B1(n_144),
.B2(n_114),
.C1(n_90),
.C2(n_169),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_15),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_301),
.B1(n_8),
.B2(n_9),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_254),
.C(n_255),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_299),
.C(n_279),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_169),
.B1(n_114),
.B2(n_3),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_114),
.C(n_2),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.C(n_1),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_1),
.C(n_3),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_7),
.B1(n_12),
.B2(n_10),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_297),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_300),
.B(n_3),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_302),
.B(n_9),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_15),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_12),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_308),
.C(n_310),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_274),
.B(n_284),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g320 ( 
.A(n_307),
.B(n_4),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_284),
.C(n_4),
.Y(n_308)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_3),
.C(n_4),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_6),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_290),
.C(n_291),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_320),
.B(n_6),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_5),
.B1(n_6),
.B2(n_313),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_304),
.B(n_306),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_325),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_327),
.Y(n_329)
);

NAND4xp25_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_5),
.C(n_6),
.D(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_318),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_315),
.B(n_326),
.C(n_329),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_328),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule