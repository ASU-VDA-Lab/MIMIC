module fake_ibex_869_n_4078 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_4078);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4078;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_3870;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_787;
wire n_2860;
wire n_2448;
wire n_4002;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1841;
wire n_1070;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_784;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_3199;
wire n_1616;
wire n_2723;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3733;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_2424;
wire n_1237;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3797;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3584;
wire n_998;
wire n_1395;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_4047;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_803;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_3948;
wire n_3719;
wire n_1599;
wire n_1539;
wire n_1400;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_817;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2352;
wire n_2263;
wire n_2212;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3908;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_4048;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_785;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_804;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3349;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_786;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3576;
wire n_3109;
wire n_1961;
wire n_3491;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_946;
wire n_1547;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_3380;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3742;
wire n_3791;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_3296;
wire n_1911;
wire n_2293;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_1488;
wire n_849;
wire n_3225;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3067;
wire n_1074;
wire n_3596;
wire n_3557;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3823;
wire n_3369;
wire n_3606;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_2148;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2961;
wire n_2996;
wire n_2704;
wire n_2770;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_3247;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2673;
wire n_2430;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_866;

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_760),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_232),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_464),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_600),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_268),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_132),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_604),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_299),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_661),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_396),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_180),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_698),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_33),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_151),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_475),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_614),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_87),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_753),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_83),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_727),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_615),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_417),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_159),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_260),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_85),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_222),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_368),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_643),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_24),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_631),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_256),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_576),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_127),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_175),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_19),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_768),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_590),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_491),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_650),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_726),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_296),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_12),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_732),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_520),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_99),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_438),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_710),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_200),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_212),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_411),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_68),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_98),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_367),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_372),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_82),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_4),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_540),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_328),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_200),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_367),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_71),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_475),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_720),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_515),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_577),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_524),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_648),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_463),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_661),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_425),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_769),
.Y(n_851)
);

BUFx10_ASAP7_75t_L g852 ( 
.A(n_89),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_364),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_739),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_170),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_458),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_247),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_331),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_530),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_210),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_559),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_406),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_66),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_40),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_359),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_730),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_549),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_469),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_389),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_552),
.Y(n_871)
);

CKINVDCx14_ASAP7_75t_R g872 ( 
.A(n_262),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_553),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_733),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_618),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_147),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_46),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_25),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_39),
.Y(n_879)
);

BUFx10_ASAP7_75t_L g880 ( 
.A(n_0),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_393),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_327),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_114),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_450),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_298),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_754),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_627),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_538),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_183),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_147),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_94),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_580),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_571),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_189),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_77),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_764),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_669),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_135),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_394),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_468),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_195),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_254),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_606),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_498),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_161),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_115),
.Y(n_907)
);

BUFx10_ASAP7_75t_L g908 ( 
.A(n_780),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_746),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_680),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_13),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_225),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_388),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_748),
.Y(n_914)
);

CKINVDCx14_ASAP7_75t_R g915 ( 
.A(n_388),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_744),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_352),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_414),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_699),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_70),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_587),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_579),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_415),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_208),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_233),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_755),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_171),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_474),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_248),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_728),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_664),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_563),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_767),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_344),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_567),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_319),
.Y(n_936)
);

BUFx10_ASAP7_75t_L g937 ( 
.A(n_696),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_744),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_614),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_539),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_772),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_137),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_526),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_720),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_741),
.Y(n_945)
);

CKINVDCx16_ASAP7_75t_R g946 ( 
.A(n_625),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_219),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_588),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_771),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_257),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_252),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_765),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_499),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_235),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_516),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_770),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_612),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_747),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_604),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_370),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_773),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_579),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_751),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_390),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_369),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_621),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_493),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_386),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_721),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_420),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_132),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_778),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_364),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_27),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_755),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_728),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_502),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_509),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_672),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_245),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_6),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_246),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_626),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_766),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_76),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_464),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_500),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_23),
.Y(n_988)
);

CKINVDCx16_ASAP7_75t_R g989 ( 
.A(n_756),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_773),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_749),
.Y(n_991)
);

BUFx2_ASAP7_75t_SL g992 ( 
.A(n_61),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_623),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_432),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_525),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_451),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_2),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_32),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_669),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_389),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_644),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_591),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_750),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_736),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_649),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_398),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_570),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_201),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_306),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_286),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_256),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_329),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_225),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_623),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_555),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_376),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_745),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_586),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_52),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_44),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_467),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_124),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_234),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_264),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_496),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_761),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_190),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_633),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_571),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_272),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_411),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_199),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_559),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_16),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_528),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_205),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_206),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_266),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_370),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_221),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_609),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_391),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_692),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_729),
.Y(n_1044)
);

BUFx8_ASAP7_75t_SL g1045 ( 
.A(n_470),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_469),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_519),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_470),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_105),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_201),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_430),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_196),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_624),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_738),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_108),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_43),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_688),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_327),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_751),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_306),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_42),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_187),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_439),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_381),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_55),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_443),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_519),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_591),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_292),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_253),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_630),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_418),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_7),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_350),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_435),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_397),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_588),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_192),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_21),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_740),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_176),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_496),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_245),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_679),
.Y(n_1084)
);

BUFx5_ASAP7_75t_L g1085 ( 
.A(n_566),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_610),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_125),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_2),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_515),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_699),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_580),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_615),
.Y(n_1092)
);

BUFx10_ASAP7_75t_L g1093 ( 
.A(n_618),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_466),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_743),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_718),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_698),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_40),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_657),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_288),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_59),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_58),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_65),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_53),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_269),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_705),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_366),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_543),
.Y(n_1108)
);

CKINVDCx16_ASAP7_75t_R g1109 ( 
.A(n_742),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_427),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_562),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_221),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_573),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_761),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_148),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_353),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_296),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_479),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_680),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_93),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_759),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_127),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_492),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_297),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_448),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_723),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_468),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_631),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_772),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_68),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_302),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_730),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_446),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_458),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_535),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_520),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_766),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_673),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_208),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_767),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_274),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_706),
.Y(n_1142)
);

CKINVDCx16_ASAP7_75t_R g1143 ( 
.A(n_454),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_175),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_589),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_382),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_427),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_750),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_384),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_351),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_691),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_111),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_692),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_115),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_242),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_205),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_66),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_305),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_172),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_533),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_131),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_589),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_352),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_737),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_196),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_611),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_335),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_612),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_34),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_445),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_565),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_268),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_662),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_597),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_209),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_251),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_758),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_605),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_299),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_442),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_609),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_206),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_57),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_545),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_676),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_303),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_734),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_467),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_735),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_567),
.Y(n_1190)
);

BUFx8_ASAP7_75t_SL g1191 ( 
.A(n_399),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_474),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_705),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_514),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_34),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_415),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_360),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_461),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_392),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_49),
.Y(n_1200)
);

CKINVDCx16_ASAP7_75t_R g1201 ( 
.A(n_616),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_709),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_660),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_616),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_562),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_732),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_139),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_321),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_610),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_139),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_180),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_298),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_305),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_754),
.Y(n_1214)
);

BUFx2_ASAP7_75t_SL g1215 ( 
.A(n_251),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_595),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_779),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_518),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_267),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_712),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_431),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_726),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_4),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_551),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_154),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_683),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_483),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_272),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_161),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_41),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_619),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_356),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_763),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_136),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_79),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_412),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_636),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_155),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_122),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_779),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_731),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_35),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_711),
.Y(n_1243)
);

BUFx10_ASAP7_75t_L g1244 ( 
.A(n_80),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_252),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_517),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_706),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_752),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_596),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_398),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_267),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_136),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_86),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_482),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_677),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_72),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_769),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_749),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_799),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1085),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_877),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_939),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_920),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_815),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_998),
.B(n_0),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_SL g1266 ( 
.A(n_880),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_815),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_831),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1223),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_939),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1235),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_831),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1085),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1256),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_872),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_915),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_939),
.Y(n_1277)
);

CKINVDCx16_ASAP7_75t_R g1278 ( 
.A(n_880),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_835),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1098),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1085),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_946),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_989),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1049),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_835),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1098),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_836),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1017),
.B(n_1043),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1077),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_911),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_836),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1017),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_863),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_811),
.B(n_0),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_894),
.B(n_1),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1043),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_863),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1193),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1193),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1258),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_984),
.B(n_1),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_864),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_864),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1258),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1183),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1182),
.B(n_1),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_793),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1109),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_822),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1183),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_880),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1133),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1045),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1202),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1191),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_841),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1143),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_988),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1034),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1231),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1144),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1061),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_895),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1079),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1088),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1201),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1252),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1090),
.B(n_3),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1102),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_942),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1130),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1157),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1169),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_818),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1195),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_832),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_911),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_792),
.B(n_2),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1200),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_838),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1244),
.Y(n_1341)
);

INVxp67_ASAP7_75t_SL g1342 ( 
.A(n_809),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_881),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1244),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_905),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1178),
.B(n_3),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_913),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_809),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1203),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1244),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_878),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1065),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_974),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_878),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_879),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_981),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_879),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_999),
.B(n_3),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_936),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1020),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1085),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_972),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1020),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_985),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1000),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1001),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_997),
.B(n_1019),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1073),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1056),
.Y(n_1369)
);

BUFx2_ASAP7_75t_SL g1370 ( 
.A(n_1085),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1073),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1129),
.B(n_1173),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_796),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1035),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_992),
.Y(n_1375)
);

XNOR2xp5_ASAP7_75t_L g1376 ( 
.A(n_1042),
.B(n_4),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_796),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_786),
.Y(n_1378)
);

CKINVDCx16_ASAP7_75t_R g1379 ( 
.A(n_786),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_819),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_819),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_830),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1259),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1266),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1278),
.B(n_1085),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1280),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1311),
.B(n_830),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1311),
.B(n_855),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1286),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1271),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1337),
.B(n_1085),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_SL g1392 ( 
.A(n_1266),
.B(n_1101),
.Y(n_1392)
);

NAND2x1_ASAP7_75t_L g1393 ( 
.A(n_1341),
.B(n_851),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1292),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1330),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1341),
.B(n_1344),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1381),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1296),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1298),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1271),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1381),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1299),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1350),
.B(n_855),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_L g1404 ( 
.A(n_1261),
.B(n_1103),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1264),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1267),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1367),
.B(n_1104),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1263),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1300),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1304),
.B(n_1230),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1342),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1269),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1348),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1262),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1274),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1268),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1340),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1352),
.B(n_1349),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1270),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1277),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1288),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1272),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1279),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1373),
.B(n_1085),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1377),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1285),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1382),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1307),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1260),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1309),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1316),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1273),
.A2(n_1361),
.B(n_1281),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1318),
.B(n_1242),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1287),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1293),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1319),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1322),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1324),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1325),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1329),
.B(n_965),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1331),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1330),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1297),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1302),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1303),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1332),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1340),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1333),
.B(n_965),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1335),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1351),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1305),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1281),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1310),
.Y(n_1454)
);

CKINVDCx16_ASAP7_75t_R g1455 ( 
.A(n_1379),
.Y(n_1455)
);

XNOR2xp5_ASAP7_75t_L g1456 ( 
.A(n_1317),
.B(n_1051),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1361),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1330),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1339),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1369),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1334),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1378),
.B(n_882),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1330),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1323),
.Y(n_1464)
);

AND2x6_ASAP7_75t_L g1465 ( 
.A(n_1294),
.B(n_1257),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1370),
.B(n_980),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1291),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1275),
.B(n_781),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1354),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1355),
.B(n_980),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1357),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1356),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1360),
.B(n_994),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1353),
.B(n_781),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1363),
.A2(n_862),
.B(n_851),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1368),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1371),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1375),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1314),
.B(n_783),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1320),
.A2(n_783),
.B1(n_789),
.B2(n_784),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1364),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1372),
.B(n_994),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1265),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1328),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1338),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1338),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1376),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1276),
.B(n_884),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1336),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1294),
.B(n_784),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1346),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1358),
.B(n_1009),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1295),
.B(n_1009),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1295),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1301),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1301),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1306),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1306),
.B(n_789),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1313),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1315),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1282),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1343),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1345),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1283),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1347),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_R g1506 ( 
.A(n_1284),
.B(n_790),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1289),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1308),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1359),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1312),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1321),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1326),
.B(n_1012),
.Y(n_1512)
);

NAND2xp33_ASAP7_75t_R g1513 ( 
.A(n_1327),
.B(n_794),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1362),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1365),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1366),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1374),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1266),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1266),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1290),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1280),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1311),
.B(n_794),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1278),
.B(n_1255),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1266),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1266),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1266),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1381),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1280),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1290),
.B(n_1012),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1266),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1266),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1280),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1280),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1266),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1280),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1280),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1280),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1278),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1290),
.B(n_1026),
.Y(n_1539)
);

BUFx10_ASAP7_75t_L g1540 ( 
.A(n_1266),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_SL g1541 ( 
.A(n_1266),
.B(n_1026),
.Y(n_1541)
);

CKINVDCx8_ASAP7_75t_R g1542 ( 
.A(n_1278),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1290),
.B(n_1066),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1259),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1266),
.Y(n_1545)
);

BUFx8_ASAP7_75t_L g1546 ( 
.A(n_1266),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1271),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1280),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1266),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1278),
.B(n_795),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1266),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1266),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1266),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1280),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1311),
.B(n_1066),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1278),
.B(n_795),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1280),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1280),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1290),
.B(n_1219),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1266),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1330),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1290),
.B(n_1219),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1311),
.B(n_1257),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1280),
.Y(n_1564)
);

CKINVDCx6p67_ASAP7_75t_R g1565 ( 
.A(n_1266),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1266),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1266),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1369),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1290),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1280),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1271),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1290),
.B(n_862),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1261),
.B(n_786),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1280),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1266),
.Y(n_1575)
);

XOR2xp5_ASAP7_75t_L g1576 ( 
.A(n_1271),
.B(n_1092),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1266),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1483),
.B(n_797),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1386),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1478),
.B(n_886),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1397),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1494),
.A2(n_785),
.B1(n_787),
.B2(n_782),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1485),
.A2(n_806),
.B(n_791),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1434),
.B(n_797),
.Y(n_1584)
);

NAND2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_857),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1527),
.Y(n_1586)
);

AND2x2_ASAP7_75t_SL g1587 ( 
.A(n_1455),
.B(n_1541),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1383),
.B(n_1215),
.Y(n_1588)
);

BUFx4f_ASAP7_75t_L g1589 ( 
.A(n_1565),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1540),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1446),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1495),
.A2(n_808),
.B1(n_820),
.B2(n_814),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1389),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1396),
.B(n_788),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1540),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1527),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1418),
.B(n_1568),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1541),
.B(n_942),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1544),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1446),
.B(n_885),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1475),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1546),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1546),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1484),
.B(n_812),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1542),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1393),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1491),
.B(n_942),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1491),
.B(n_942),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1486),
.B(n_889),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1475),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1496),
.A2(n_825),
.B1(n_837),
.B2(n_824),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1407),
.B(n_890),
.Y(n_1613)
);

AND2x6_ASAP7_75t_L g1614 ( 
.A(n_1496),
.B(n_893),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1520),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1556),
.B(n_812),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1521),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1528),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1433),
.Y(n_1619)
);

AND2x2_ASAP7_75t_SL g1620 ( 
.A(n_1435),
.B(n_893),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1464),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1396),
.B(n_839),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1532),
.Y(n_1623)
);

BUFx4f_ASAP7_75t_L g1624 ( 
.A(n_1491),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1404),
.B(n_853),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1522),
.B(n_891),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1496),
.B(n_942),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1434),
.B(n_798),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1451),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1424),
.B(n_800),
.C(n_798),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1451),
.Y(n_1631)
);

AO21x1_ASAP7_75t_L g1632 ( 
.A1(n_1391),
.A2(n_1539),
.B(n_1529),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_SL g1633 ( 
.A(n_1512),
.Y(n_1633)
);

CKINVDCx11_ASAP7_75t_R g1634 ( 
.A(n_1408),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1479),
.B(n_1480),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1411),
.B(n_800),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1533),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1460),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1535),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1536),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1476),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1412),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1429),
.B(n_801),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1497),
.A2(n_859),
.B1(n_861),
.B2(n_856),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1424),
.B(n_802),
.C(n_801),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1573),
.B(n_812),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1537),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1413),
.B(n_892),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1497),
.B(n_954),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1436),
.B(n_816),
.Y(n_1650)
);

INVx6_ASAP7_75t_L g1651 ( 
.A(n_1387),
.Y(n_1651)
);

AND2x6_ASAP7_75t_L g1652 ( 
.A(n_1497),
.B(n_900),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1548),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1554),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1444),
.B(n_1467),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1557),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1474),
.B(n_816),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1415),
.Y(n_1658)
);

INVx4_ASAP7_75t_L g1659 ( 
.A(n_1384),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1501),
.B(n_1507),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1555),
.Y(n_1661)
);

AND2x6_ASAP7_75t_L g1662 ( 
.A(n_1387),
.B(n_900),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1431),
.B(n_954),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1462),
.B(n_896),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1508),
.B(n_802),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1555),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1388),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1388),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1432),
.B(n_803),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1569),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1401),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1466),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1472),
.Y(n_1674)
);

NAND3x1_ASAP7_75t_L g1675 ( 
.A(n_1514),
.B(n_1126),
.C(n_1113),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1518),
.Y(n_1676)
);

AND2x2_ASAP7_75t_SL g1677 ( 
.A(n_1512),
.B(n_910),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1558),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1439),
.B(n_803),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1564),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1490),
.B(n_897),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1563),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1498),
.B(n_1385),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1510),
.B(n_804),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1506),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1570),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1466),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1469),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1574),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1405),
.B(n_852),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1440),
.B(n_954),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1563),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1403),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1471),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1442),
.B(n_804),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1394),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1410),
.B(n_898),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1403),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1406),
.B(n_852),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1398),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1492),
.B(n_867),
.Y(n_1701)
);

CKINVDCx16_ASAP7_75t_R g1702 ( 
.A(n_1468),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1416),
.B(n_852),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1481),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1422),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1423),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1477),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1425),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1519),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1426),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1489),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1447),
.B(n_805),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1493),
.B(n_899),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1399),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1493),
.B(n_1523),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1402),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1450),
.B(n_954),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1459),
.B(n_1414),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1409),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1492),
.B(n_954),
.Y(n_1720)
);

NAND2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1550),
.B(n_888),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1419),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1420),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1441),
.B(n_805),
.Y(n_1724)
);

AND2x4_ASAP7_75t_SL g1725 ( 
.A(n_1516),
.B(n_1504),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1499),
.B(n_1500),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1441),
.B(n_807),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1449),
.B(n_807),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1449),
.B(n_810),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1502),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1465),
.A2(n_813),
.B1(n_817),
.B2(n_810),
.Y(n_1731)
);

CKINVDCx6p67_ASAP7_75t_R g1732 ( 
.A(n_1516),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1427),
.Y(n_1733)
);

INVx8_ASAP7_75t_L g1734 ( 
.A(n_1524),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1465),
.B(n_813),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1421),
.B(n_901),
.Y(n_1736)
);

INVx4_ASAP7_75t_L g1737 ( 
.A(n_1525),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1572),
.A2(n_1141),
.B1(n_1160),
.B2(n_1128),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1482),
.B(n_902),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1392),
.B(n_1032),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1465),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1428),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1445),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1452),
.Y(n_1744)
);

INVx4_ASAP7_75t_SL g1745 ( 
.A(n_1516),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1572),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1454),
.B(n_908),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1529),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1539),
.B(n_821),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1543),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1543),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1559),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1559),
.A2(n_823),
.B1(n_826),
.B2(n_821),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1562),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1562),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1470),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1470),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1473),
.B(n_823),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1473),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1391),
.Y(n_1760)
);

AND2x6_ASAP7_75t_L g1761 ( 
.A(n_1482),
.B(n_910),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1511),
.B(n_978),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1430),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1526),
.B(n_903),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1390),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1530),
.A2(n_1192),
.B1(n_1245),
.B2(n_1166),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1453),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1531),
.B(n_1534),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1545),
.B(n_904),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1395),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1457),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1549),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1551),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1552),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_SL g1775 ( 
.A(n_1553),
.B(n_1567),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1395),
.Y(n_1776)
);

AND2x6_ASAP7_75t_L g1777 ( 
.A(n_1488),
.B(n_978),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1560),
.B(n_1032),
.Y(n_1778)
);

OR2x6_ASAP7_75t_L g1779 ( 
.A(n_1487),
.B(n_979),
.Y(n_1779)
);

OR2x6_ASAP7_75t_L g1780 ( 
.A(n_1513),
.B(n_979),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1566),
.A2(n_875),
.B1(n_883),
.B2(n_873),
.Y(n_1781)
);

INVx4_ASAP7_75t_L g1782 ( 
.A(n_1575),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1505),
.B(n_907),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1395),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1443),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1443),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1509),
.B(n_912),
.Y(n_1787)
);

OR2x6_ASAP7_75t_L g1788 ( 
.A(n_1517),
.B(n_993),
.Y(n_1788)
);

AND2x6_ASAP7_75t_L g1789 ( 
.A(n_1458),
.B(n_993),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1576),
.B(n_826),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1458),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1461),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1400),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1463),
.B(n_827),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1463),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1456),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1561),
.B(n_827),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1561),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1547),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1571),
.B(n_914),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1503),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1417),
.B(n_916),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1448),
.B(n_917),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1515),
.A2(n_906),
.B1(n_923),
.B2(n_887),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1483),
.B(n_828),
.Y(n_1805)
);

AND2x6_ASAP7_75t_L g1806 ( 
.A(n_1483),
.B(n_995),
.Y(n_1806)
);

INVx4_ASAP7_75t_L g1807 ( 
.A(n_1540),
.Y(n_1807)
);

OR2x6_ASAP7_75t_L g1808 ( 
.A(n_1538),
.B(n_995),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1478),
.B(n_919),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1386),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1546),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1478),
.B(n_921),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1386),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1483),
.B(n_925),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1397),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1386),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1475),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1475),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1483),
.B(n_828),
.Y(n_1819)
);

AND3x1_ASAP7_75t_L g1820 ( 
.A(n_1488),
.B(n_928),
.C(n_926),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1386),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1397),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1556),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1483),
.B(n_829),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1478),
.B(n_922),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1386),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1418),
.B(n_908),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1418),
.B(n_908),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1483),
.B(n_829),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1483),
.A2(n_933),
.B1(n_938),
.B2(n_929),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1386),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1397),
.Y(n_1832)
);

AO21x2_ASAP7_75t_L g1833 ( 
.A1(n_1433),
.A2(n_943),
.B(n_940),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1483),
.B(n_833),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1386),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1541),
.B(n_1032),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1418),
.B(n_909),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1478),
.B(n_924),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1541),
.B(n_1032),
.Y(n_1839)
);

CKINVDCx16_ASAP7_75t_R g1840 ( 
.A(n_1556),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1386),
.Y(n_1841)
);

CKINVDCx16_ASAP7_75t_R g1842 ( 
.A(n_1556),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1591),
.A2(n_1655),
.B1(n_1597),
.B2(n_1646),
.Y(n_1843)
);

AND2x6_ASAP7_75t_SL g1844 ( 
.A(n_1788),
.B(n_945),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1738),
.B(n_1251),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1635),
.A2(n_952),
.B1(n_959),
.B2(n_947),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1579),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1593),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1634),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1738),
.B(n_1255),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1756),
.B(n_833),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1591),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1757),
.B(n_834),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1715),
.A2(n_840),
.B1(n_842),
.B2(n_834),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1814),
.A2(n_1806),
.B1(n_1630),
.B2(n_1645),
.Y(n_1855)
);

NOR2xp67_ASAP7_75t_L g1856 ( 
.A(n_1590),
.B(n_5),
.Y(n_1856)
);

NAND2x1_ASAP7_75t_L g1857 ( 
.A(n_1714),
.B(n_1032),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1759),
.B(n_1251),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1814),
.A2(n_842),
.B1(n_843),
.B2(n_840),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1806),
.A2(n_844),
.B1(n_845),
.B2(n_843),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1600),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1806),
.A2(n_971),
.B1(n_975),
.B2(n_962),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1590),
.B(n_976),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1617),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1683),
.A2(n_1750),
.B(n_1751),
.C(n_1748),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1746),
.B(n_844),
.Y(n_1866)
);

O2A1O1Ixp5_ASAP7_75t_L g1867 ( 
.A1(n_1632),
.A2(n_1095),
.B(n_1111),
.C(n_1087),
.Y(n_1867)
);

OAI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1599),
.A2(n_1248),
.B1(n_846),
.B2(n_847),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1618),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1808),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1578),
.B(n_1805),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1578),
.B(n_845),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1718),
.A2(n_1004),
.B1(n_1005),
.B2(n_991),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1638),
.B(n_846),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1805),
.B(n_847),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1766),
.B(n_848),
.Y(n_1876)
);

BUFx3_ASAP7_75t_L g1877 ( 
.A(n_1732),
.Y(n_1877)
);

NOR3xp33_ASAP7_75t_L g1878 ( 
.A(n_1766),
.B(n_1243),
.C(n_951),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1808),
.Y(n_1879)
);

BUFx12f_ASAP7_75t_L g1880 ( 
.A(n_1602),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1672),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1718),
.A2(n_1023),
.B1(n_1036),
.B2(n_1006),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1819),
.B(n_848),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1808),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1819),
.B(n_849),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1687),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1824),
.B(n_850),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1824),
.B(n_850),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1623),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1827),
.B(n_854),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1687),
.B(n_1624),
.Y(n_1891)
);

A2O1A1Ixp33_ASAP7_75t_L g1892 ( 
.A1(n_1752),
.A2(n_1044),
.B(n_1046),
.C(n_1037),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1829),
.B(n_858),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1741),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1629),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1637),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1828),
.B(n_1837),
.Y(n_1897)
);

NAND2xp33_ASAP7_75t_L g1898 ( 
.A(n_1741),
.B(n_858),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1639),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1661),
.B(n_1666),
.Y(n_1900)
);

OR2x6_ASAP7_75t_L g1901 ( 
.A(n_1734),
.B(n_1087),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1640),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1834),
.B(n_860),
.Y(n_1903)
);

NAND2x1p5_ASAP7_75t_L g1904 ( 
.A(n_1661),
.B(n_1095),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1834),
.B(n_860),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1587),
.A2(n_1120),
.B1(n_1142),
.B2(n_868),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1724),
.B(n_865),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1650),
.B(n_865),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1724),
.B(n_866),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1630),
.A2(n_1057),
.B1(n_1059),
.B2(n_1054),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1629),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1631),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1727),
.B(n_866),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1727),
.B(n_868),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1647),
.Y(n_1915)
);

INVxp33_ASAP7_75t_SL g1916 ( 
.A(n_1705),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1758),
.B(n_869),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1631),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1731),
.A2(n_871),
.B1(n_874),
.B2(n_870),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1584),
.A2(n_1081),
.B1(n_1089),
.B2(n_1071),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1661),
.B(n_870),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1653),
.Y(n_1922)
);

OAI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1840),
.A2(n_874),
.B1(n_876),
.B2(n_871),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1584),
.B(n_876),
.Y(n_1924)
);

NAND3xp33_ASAP7_75t_L g1925 ( 
.A(n_1783),
.B(n_1118),
.C(n_1117),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1628),
.B(n_1749),
.Y(n_1926)
);

BUFx12f_ASAP7_75t_L g1927 ( 
.A(n_1603),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1654),
.Y(n_1928)
);

INVx8_ASAP7_75t_L g1929 ( 
.A(n_1734),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1714),
.B(n_1119),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1716),
.B(n_1120),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1716),
.B(n_1122),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1719),
.B(n_1122),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1719),
.B(n_1123),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1620),
.B(n_1123),
.Y(n_1935)
);

BUFx8_ASAP7_75t_L g1936 ( 
.A(n_1633),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1754),
.B(n_1131),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1628),
.B(n_1131),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1656),
.B(n_1134),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1592),
.A2(n_1099),
.B1(n_1100),
.B2(n_1091),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1631),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1678),
.B(n_1134),
.Y(n_1942)
);

AND2x6_ASAP7_75t_SL g1943 ( 
.A(n_1788),
.B(n_1106),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1680),
.B(n_1136),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1657),
.B(n_1136),
.Y(n_1945)
);

NAND2x1p5_ASAP7_75t_L g1946 ( 
.A(n_1666),
.B(n_1111),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1686),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1689),
.B(n_1137),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1820),
.A2(n_1753),
.B1(n_1594),
.B2(n_1713),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1696),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1700),
.B(n_1137),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1760),
.A2(n_1121),
.B(n_1108),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1645),
.A2(n_1125),
.B1(n_1127),
.B2(n_1124),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1820),
.A2(n_1140),
.B1(n_1142),
.B2(n_1138),
.Y(n_1954)
);

NAND3xp33_ASAP7_75t_SL g1955 ( 
.A(n_1711),
.B(n_1140),
.C(n_1138),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1810),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1813),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1585),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1666),
.B(n_1145),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1641),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1790),
.B(n_1793),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1651),
.B(n_1145),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1589),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1614),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1749),
.B(n_1643),
.Y(n_1965)
);

A2O1A1Ixp33_ASAP7_75t_L g1966 ( 
.A1(n_1816),
.A2(n_1151),
.B(n_1152),
.C(n_1132),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1601),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1811),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1610),
.A2(n_1755),
.B1(n_1669),
.B2(n_1679),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_SL g1970 ( 
.A(n_1605),
.Y(n_1970)
);

A2O1A1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1821),
.A2(n_1165),
.B(n_1168),
.C(n_1159),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1643),
.A2(n_1174),
.B1(n_1177),
.B2(n_1170),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1669),
.B(n_1146),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1651),
.B(n_1146),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1679),
.B(n_1147),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1826),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1831),
.Y(n_1977)
);

BUFx3_ASAP7_75t_L g1978 ( 
.A(n_1792),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1695),
.B(n_1147),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1695),
.B(n_1149),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1673),
.A2(n_1712),
.B(n_1735),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1712),
.B(n_1149),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1835),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1665),
.B(n_1150),
.Y(n_1984)
);

O2A1O1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1636),
.A2(n_1180),
.B(n_1184),
.C(n_1179),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1684),
.B(n_1150),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1728),
.B(n_1153),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1677),
.B(n_1153),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1601),
.Y(n_1989)
);

A2O1A1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1841),
.A2(n_1204),
.B(n_1208),
.C(n_1187),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1601),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1729),
.B(n_1154),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1753),
.B(n_1154),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1613),
.B(n_1155),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1761),
.A2(n_1662),
.B1(n_1693),
.B2(n_1692),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1642),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1594),
.A2(n_1681),
.B1(n_1662),
.B2(n_1625),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1761),
.A2(n_1216),
.B1(n_1225),
.B2(n_1209),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1706),
.B(n_1733),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1611),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1722),
.B(n_1155),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1604),
.B(n_1156),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1611),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1588),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1723),
.B(n_1688),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1694),
.B(n_1158),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1707),
.B(n_1158),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1743),
.B(n_1161),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1744),
.B(n_1162),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1708),
.B(n_1162),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1662),
.A2(n_1167),
.B1(n_1171),
.B2(n_1163),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1710),
.B(n_1163),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1742),
.B(n_1167),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1621),
.B(n_1171),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1616),
.B(n_1172),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1693),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1830),
.B(n_1172),
.Y(n_2017)
);

INVx4_ASAP7_75t_L g2018 ( 
.A(n_1595),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1595),
.B(n_1175),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_1800),
.B(n_1803),
.C(n_1802),
.Y(n_2020)
);

BUFx3_ASAP7_75t_L g2021 ( 
.A(n_1807),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1583),
.B(n_1175),
.Y(n_2022)
);

INVx8_ASAP7_75t_L g2023 ( 
.A(n_1734),
.Y(n_2023)
);

OR2x6_ASAP7_75t_L g2024 ( 
.A(n_1588),
.B(n_1189),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1817),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1625),
.B(n_1176),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1690),
.B(n_1181),
.Y(n_2027)
);

NAND2x1p5_ASAP7_75t_L g2028 ( 
.A(n_1615),
.B(n_1189),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1583),
.B(n_1181),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1699),
.B(n_1185),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1703),
.B(n_1185),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1619),
.A2(n_1232),
.B(n_1226),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1747),
.B(n_1186),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1761),
.B(n_1186),
.Y(n_2034)
);

AOI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1619),
.A2(n_1234),
.B(n_1247),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1817),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1761),
.B(n_1190),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1662),
.B(n_1194),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1818),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1818),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1725),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1745),
.B(n_1249),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1582),
.B(n_1194),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1726),
.B(n_1196),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1612),
.B(n_1196),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1668),
.B(n_1197),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1644),
.B(n_1197),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1622),
.B(n_927),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1622),
.B(n_930),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1667),
.A2(n_1253),
.B1(n_1254),
.B2(n_1250),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1674),
.B(n_909),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1692),
.Y(n_2052)
);

A2O1A1Ixp33_ASAP7_75t_SL g2053 ( 
.A1(n_1664),
.A2(n_1213),
.B(n_1221),
.C(n_1207),
.Y(n_2053)
);

BUFx5_ASAP7_75t_L g2054 ( 
.A(n_1789),
.Y(n_2054)
);

INVx2_ASAP7_75t_SL g2055 ( 
.A(n_1704),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1762),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1762),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1698),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1682),
.B(n_932),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1619),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1648),
.B(n_934),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1701),
.B(n_935),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1660),
.B(n_941),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_1762),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1701),
.B(n_1614),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_1780),
.Y(n_2066)
);

OAI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1763),
.A2(n_1213),
.B(n_1207),
.Y(n_2067)
);

AND2x6_ASAP7_75t_SL g2068 ( 
.A(n_1779),
.B(n_1780),
.Y(n_2068)
);

OR2x6_ASAP7_75t_SL g2069 ( 
.A(n_1658),
.B(n_944),
.Y(n_2069)
);

NAND2x1_ASAP7_75t_L g2070 ( 
.A(n_1614),
.B(n_1058),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1833),
.A2(n_1221),
.B(n_949),
.Y(n_2071)
);

NOR2xp67_ASAP7_75t_L g2072 ( 
.A(n_1607),
.B(n_5),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1626),
.B(n_948),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1720),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1581),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1606),
.B(n_950),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1606),
.B(n_953),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1840),
.Y(n_2078)
);

AND2x4_ASAP7_75t_L g2079 ( 
.A(n_1745),
.B(n_918),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1614),
.B(n_955),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1739),
.B(n_956),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1823),
.B(n_909),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1607),
.B(n_957),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1721),
.B(n_960),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1586),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1659),
.B(n_958),
.Y(n_2086)
);

OR2x6_ASAP7_75t_L g2087 ( 
.A(n_1779),
.B(n_1659),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1697),
.B(n_961),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1676),
.B(n_963),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1596),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1670),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1676),
.B(n_964),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1580),
.B(n_1825),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1671),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1809),
.B(n_966),
.Y(n_2095)
);

INVx5_ASAP7_75t_L g2096 ( 
.A(n_1652),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1709),
.B(n_967),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_1777),
.A2(n_969),
.B1(n_970),
.B2(n_968),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1812),
.B(n_973),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_1793),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_1685),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1709),
.B(n_977),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1815),
.Y(n_2103)
);

AND2x6_ASAP7_75t_SL g2104 ( 
.A(n_1801),
.B(n_1799),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1842),
.B(n_931),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1737),
.B(n_982),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1737),
.B(n_983),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1842),
.B(n_931),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1633),
.B(n_986),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1652),
.A2(n_937),
.B1(n_990),
.B2(n_931),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1822),
.Y(n_2111)
);

INVx4_ASAP7_75t_L g2112 ( 
.A(n_1782),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1782),
.B(n_987),
.Y(n_2113)
);

OAI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_1702),
.A2(n_1224),
.B1(n_1227),
.B2(n_1222),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_SL g2115 ( 
.A(n_1652),
.B(n_937),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1794),
.B(n_996),
.Y(n_2116)
);

INVx3_ASAP7_75t_L g2117 ( 
.A(n_1832),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_1772),
.B(n_1018),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1767),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1838),
.B(n_1002),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1804),
.B(n_937),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_1787),
.B(n_1773),
.Y(n_2122)
);

NAND2xp33_ASAP7_75t_SL g2123 ( 
.A(n_1768),
.B(n_1238),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_1774),
.B(n_1003),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1797),
.B(n_1007),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1652),
.B(n_1008),
.Y(n_2126)
);

AOI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_1777),
.A2(n_1736),
.B1(n_1781),
.B2(n_1769),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1771),
.B(n_1010),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1775),
.B(n_1011),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_1764),
.B(n_1013),
.Y(n_2130)
);

BUFx3_ASAP7_75t_L g2131 ( 
.A(n_1765),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1608),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1775),
.B(n_1014),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1730),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1777),
.B(n_1015),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_1675),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1777),
.B(n_1016),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1609),
.Y(n_2138)
);

OR2x6_ASAP7_75t_L g2139 ( 
.A(n_1796),
.B(n_1058),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1740),
.B(n_1021),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_1778),
.A2(n_1093),
.B1(n_1164),
.B2(n_990),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1847),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1848),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_1929),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1864),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1871),
.B(n_1627),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_2060),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1869),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1889),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_2060),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1896),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1871),
.B(n_1649),
.Y(n_2152)
);

NOR3xp33_ASAP7_75t_SL g2153 ( 
.A(n_1849),
.B(n_1024),
.C(n_1022),
.Y(n_2153)
);

INVx4_ASAP7_75t_L g2154 ( 
.A(n_1929),
.Y(n_2154)
);

A2O1A1Ixp33_ASAP7_75t_L g2155 ( 
.A1(n_1865),
.A2(n_1836),
.B(n_1839),
.C(n_1598),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1899),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1916),
.B(n_1025),
.Y(n_2157)
);

AOI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_1868),
.A2(n_1027),
.B1(n_1029),
.B2(n_1028),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1902),
.Y(n_2159)
);

NOR3xp33_ASAP7_75t_SL g2160 ( 
.A(n_1996),
.B(n_1031),
.C(n_1030),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1915),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1852),
.B(n_990),
.Y(n_2162)
);

BUFx10_ASAP7_75t_L g2163 ( 
.A(n_1970),
.Y(n_2163)
);

NOR3xp33_ASAP7_75t_SL g2164 ( 
.A(n_1955),
.B(n_1038),
.C(n_1033),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_1900),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_2086),
.B(n_1039),
.Y(n_2166)
);

INVx4_ASAP7_75t_L g2167 ( 
.A(n_1929),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1926),
.B(n_1040),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_2060),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1922),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1928),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1947),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_2018),
.B(n_1795),
.Y(n_2173)
);

INVx2_ASAP7_75t_SL g2174 ( 
.A(n_2023),
.Y(n_2174)
);

NOR3xp33_ASAP7_75t_SL g2175 ( 
.A(n_2123),
.B(n_1047),
.C(n_1041),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_2018),
.B(n_1795),
.Y(n_2176)
);

O2A1O1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_1892),
.A2(n_1139),
.B(n_1188),
.C(n_1148),
.Y(n_2177)
);

BUFx2_ASAP7_75t_SL g2178 ( 
.A(n_2021),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1950),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1956),
.Y(n_2180)
);

NOR3xp33_ASAP7_75t_SL g2181 ( 
.A(n_2122),
.B(n_1050),
.C(n_1048),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1965),
.B(n_1052),
.Y(n_2182)
);

A2O1A1Ixp33_ASAP7_75t_L g2183 ( 
.A1(n_1981),
.A2(n_1691),
.B(n_1717),
.C(n_1663),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_2086),
.B(n_1053),
.Y(n_2184)
);

INVx3_ASAP7_75t_L g2185 ( 
.A(n_1900),
.Y(n_2185)
);

NAND2xp33_ASAP7_75t_SL g2186 ( 
.A(n_2112),
.B(n_1055),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1957),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1976),
.B(n_1060),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1977),
.Y(n_2189)
);

AND2x6_ASAP7_75t_L g2190 ( 
.A(n_1964),
.B(n_1058),
.Y(n_2190)
);

INVxp67_ASAP7_75t_L g2191 ( 
.A(n_2100),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1880),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1983),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_2112),
.B(n_1789),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1969),
.B(n_1062),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1897),
.B(n_1961),
.Y(n_2196)
);

BUFx3_ASAP7_75t_L g2197 ( 
.A(n_2023),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1949),
.B(n_1063),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2005),
.Y(n_2199)
);

CKINVDCx8_ASAP7_75t_R g2200 ( 
.A(n_2023),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_1936),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1872),
.B(n_1064),
.Y(n_2202)
);

AO22x1_ASAP7_75t_L g2203 ( 
.A1(n_1936),
.A2(n_1789),
.B1(n_1069),
.B2(n_1072),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1872),
.B(n_1068),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2119),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1937),
.Y(n_2206)
);

CKINVDCx16_ASAP7_75t_R g2207 ( 
.A(n_2069),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_L g2208 ( 
.A(n_1879),
.B(n_1074),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1875),
.B(n_1075),
.Y(n_2209)
);

INVx2_ASAP7_75t_SL g2210 ( 
.A(n_1877),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_2096),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_1870),
.B(n_1789),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1861),
.B(n_1076),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1937),
.Y(n_2214)
);

BUFx4f_ASAP7_75t_L g2215 ( 
.A(n_1927),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1875),
.B(n_1078),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1883),
.B(n_1080),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1930),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_L g2219 ( 
.A(n_1884),
.B(n_1082),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1930),
.Y(n_2220)
);

INVx8_ASAP7_75t_L g2221 ( 
.A(n_1901),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1901),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_1958),
.B(n_5),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_2004),
.B(n_6),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2096),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1883),
.B(n_1083),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_2096),
.Y(n_2227)
);

BUFx2_ASAP7_75t_L g2228 ( 
.A(n_2087),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_2087),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2087),
.B(n_6),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1931),
.Y(n_2231)
);

BUFx2_ASAP7_75t_L g2232 ( 
.A(n_1901),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_1845),
.B(n_1210),
.Y(n_2233)
);

INVx4_ASAP7_75t_L g2234 ( 
.A(n_2068),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1999),
.A2(n_1086),
.B1(n_1094),
.B2(n_1084),
.Y(n_2235)
);

OR2x4_ASAP7_75t_L g2236 ( 
.A(n_1876),
.B(n_1058),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_2139),
.Y(n_2237)
);

BUFx4f_ASAP7_75t_L g2238 ( 
.A(n_2024),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2056),
.B(n_7),
.Y(n_2239)
);

NAND3xp33_ASAP7_75t_SL g2240 ( 
.A(n_2127),
.B(n_1220),
.C(n_1105),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1843),
.B(n_1096),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1885),
.B(n_1107),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1885),
.B(n_1110),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1866),
.B(n_1112),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1866),
.B(n_1114),
.Y(n_2245)
);

CKINVDCx16_ASAP7_75t_R g2246 ( 
.A(n_2024),
.Y(n_2246)
);

AOI22x1_ASAP7_75t_L g2247 ( 
.A1(n_2071),
.A2(n_1791),
.B1(n_1798),
.B2(n_1784),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_2024),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1931),
.Y(n_2249)
);

INVx4_ASAP7_75t_L g2250 ( 
.A(n_1844),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1932),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_R g2252 ( 
.A(n_2078),
.B(n_1115),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1932),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_1850),
.B(n_1116),
.Y(n_2254)
);

BUFx4f_ASAP7_75t_L g2255 ( 
.A(n_2139),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1935),
.B(n_1093),
.Y(n_2256)
);

AOI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_1878),
.A2(n_1164),
.B1(n_1093),
.B2(n_1198),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1988),
.B(n_1164),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1933),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1970),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1851),
.B(n_1199),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1933),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2091),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1934),
.Y(n_2264)
);

NOR3xp33_ASAP7_75t_SL g2265 ( 
.A(n_2114),
.B(n_1923),
.C(n_2129),
.Y(n_2265)
);

AOI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_2020),
.A2(n_1206),
.B1(n_1211),
.B2(n_1205),
.Y(n_2266)
);

BUFx12f_ASAP7_75t_L g2267 ( 
.A(n_2055),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_1860),
.B(n_1212),
.Y(n_2268)
);

NAND2x1_ASAP7_75t_L g2269 ( 
.A(n_1895),
.B(n_1784),
.Y(n_2269)
);

BUFx8_ASAP7_75t_L g2270 ( 
.A(n_1968),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2115),
.B(n_1214),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_2096),
.Y(n_2272)
);

INVx3_ASAP7_75t_L g2273 ( 
.A(n_1960),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2121),
.A2(n_1218),
.B1(n_1228),
.B2(n_1217),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1984),
.B(n_1986),
.Y(n_2275)
);

NOR3xp33_ASAP7_75t_SL g2276 ( 
.A(n_2133),
.B(n_1233),
.C(n_1229),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1851),
.B(n_1236),
.Y(n_2277)
);

INVx3_ASAP7_75t_L g2278 ( 
.A(n_1960),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_1895),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1853),
.B(n_1237),
.Y(n_2280)
);

NAND2x1p5_ASAP7_75t_L g2281 ( 
.A(n_1964),
.B(n_1067),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_2115),
.B(n_2011),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_1967),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1934),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2139),
.Y(n_2285)
);

BUFx12f_ASAP7_75t_L g2286 ( 
.A(n_1943),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2094),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_1862),
.A2(n_1070),
.B1(n_1097),
.B2(n_1067),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1853),
.B(n_1858),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2057),
.B(n_1239),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1858),
.B(n_1240),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_1904),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_1978),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1846),
.B(n_1241),
.Y(n_2294)
);

INVx5_ASAP7_75t_L g2295 ( 
.A(n_2064),
.Y(n_2295)
);

BUFx12f_ASAP7_75t_L g2296 ( 
.A(n_2104),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2006),
.Y(n_2297)
);

INVx1_ASAP7_75t_SL g2298 ( 
.A(n_2131),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2016),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2006),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1920),
.B(n_1952),
.Y(n_2301)
);

INVxp67_ASAP7_75t_SL g2302 ( 
.A(n_1904),
.Y(n_2302)
);

AND2x2_ASAP7_75t_SL g2303 ( 
.A(n_2079),
.B(n_1067),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2052),
.Y(n_2304)
);

NOR3xp33_ASAP7_75t_SL g2305 ( 
.A(n_1920),
.B(n_1246),
.C(n_7),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2063),
.B(n_8),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2013),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2013),
.Y(n_2308)
);

INVx1_ASAP7_75t_SL g2309 ( 
.A(n_2065),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2007),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2010),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_R g2312 ( 
.A(n_1963),
.B(n_8),
.Y(n_2312)
);

AOI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_1945),
.A2(n_1070),
.B1(n_1097),
.B2(n_1067),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2012),
.Y(n_2314)
);

NAND3xp33_ASAP7_75t_SL g2315 ( 
.A(n_1997),
.B(n_1786),
.C(n_1776),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_2134),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2103),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_1989),
.Y(n_2318)
);

INVx4_ASAP7_75t_L g2319 ( 
.A(n_2079),
.Y(n_2319)
);

INVx4_ASAP7_75t_L g2320 ( 
.A(n_2054),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1906),
.B(n_1770),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1972),
.B(n_8),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1939),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2111),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_2028),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_2008),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1939),
.B(n_9),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_2009),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1942),
.B(n_9),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_SL g2330 ( 
.A(n_1925),
.B(n_9),
.C(n_10),
.Y(n_2330)
);

BUFx2_ASAP7_75t_L g2331 ( 
.A(n_2014),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1942),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1944),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_R g2334 ( 
.A(n_2136),
.B(n_10),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1944),
.B(n_10),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1948),
.Y(n_2336)
);

BUFx5_ASAP7_75t_L g2337 ( 
.A(n_2138),
.Y(n_2337)
);

INVx4_ASAP7_75t_L g2338 ( 
.A(n_2054),
.Y(n_2338)
);

INVx4_ASAP7_75t_L g2339 ( 
.A(n_2054),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_1991),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2015),
.B(n_11),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_L g2342 ( 
.A1(n_1890),
.A2(n_1097),
.B1(n_1135),
.B2(n_1070),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1948),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_1908),
.A2(n_1097),
.B1(n_1135),
.B2(n_1070),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2066),
.B(n_11),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2044),
.B(n_2098),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2101),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2118),
.B(n_1770),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2083),
.B(n_2089),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1951),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1951),
.B(n_11),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_1993),
.B(n_12),
.Y(n_2352)
);

NOR3xp33_ASAP7_75t_SL g2353 ( 
.A(n_1966),
.B(n_13),
.C(n_14),
.Y(n_2353)
);

OR2x2_ASAP7_75t_L g2354 ( 
.A(n_1859),
.B(n_13),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_1938),
.B(n_1910),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_R g2356 ( 
.A(n_2041),
.B(n_14),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2058),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2001),
.Y(n_2358)
);

BUFx2_ASAP7_75t_L g2359 ( 
.A(n_2028),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2002),
.B(n_14),
.Y(n_2360)
);

INVx1_ASAP7_75t_SL g2361 ( 
.A(n_2065),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1881),
.Y(n_2362)
);

BUFx4f_ASAP7_75t_L g2363 ( 
.A(n_1863),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1886),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2042),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_1946),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1953),
.B(n_1855),
.Y(n_2367)
);

INVx2_ASAP7_75t_SL g2368 ( 
.A(n_1863),
.Y(n_2368)
);

BUFx3_ASAP7_75t_L g2369 ( 
.A(n_2042),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2075),
.Y(n_2370)
);

NOR3xp33_ASAP7_75t_SL g2371 ( 
.A(n_1971),
.B(n_15),
.C(n_16),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2118),
.B(n_1785),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2093),
.B(n_15),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2085),
.Y(n_2374)
);

OR2x6_ASAP7_75t_L g2375 ( 
.A(n_1856),
.B(n_1135),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_1946),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2090),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2092),
.B(n_2097),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2117),
.Y(n_2379)
);

CKINVDCx6p67_ASAP7_75t_R g2380 ( 
.A(n_2105),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_2108),
.Y(n_2381)
);

NOR3xp33_ASAP7_75t_SL g2382 ( 
.A(n_1990),
.B(n_15),
.C(n_16),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2067),
.B(n_17),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1887),
.Y(n_2384)
);

CKINVDCx14_ASAP7_75t_R g2385 ( 
.A(n_2051),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2067),
.B(n_17),
.Y(n_2386)
);

CKINVDCx20_ASAP7_75t_R g2387 ( 
.A(n_1954),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1888),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_1854),
.B(n_17),
.Y(n_2389)
);

CKINVDCx20_ASAP7_75t_R g2390 ( 
.A(n_1919),
.Y(n_2390)
);

BUFx5_ASAP7_75t_L g2391 ( 
.A(n_2074),
.Y(n_2391)
);

BUFx3_ASAP7_75t_L g2392 ( 
.A(n_2082),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2027),
.B(n_18),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1893),
.B(n_1903),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1905),
.Y(n_2395)
);

BUFx3_ASAP7_75t_L g2396 ( 
.A(n_2109),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1973),
.Y(n_2397)
);

AND2x6_ASAP7_75t_SL g2398 ( 
.A(n_2084),
.B(n_18),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2000),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_1857),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1911),
.Y(n_2401)
);

NOR3xp33_ASAP7_75t_SL g2402 ( 
.A(n_1940),
.B(n_19),
.C(n_20),
.Y(n_2402)
);

INVxp67_ASAP7_75t_L g2403 ( 
.A(n_2038),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1975),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_1924),
.B(n_19),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_1979),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1907),
.B(n_20),
.Y(n_2407)
);

AND2x6_ASAP7_75t_L g2408 ( 
.A(n_1912),
.B(n_1918),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_2072),
.B(n_1874),
.Y(n_2409)
);

INVx5_ASAP7_75t_L g2410 ( 
.A(n_1941),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_R g2411 ( 
.A(n_1898),
.B(n_20),
.Y(n_2411)
);

OR2x2_ASAP7_75t_SL g2412 ( 
.A(n_2022),
.B(n_21),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2034),
.B(n_22),
.Y(n_2413)
);

BUFx2_ASAP7_75t_L g2414 ( 
.A(n_2034),
.Y(n_2414)
);

INVx5_ASAP7_75t_L g2415 ( 
.A(n_2003),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1980),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_1909),
.B(n_22),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1867),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_L g2419 ( 
.A(n_2130),
.B(n_2110),
.C(n_2053),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1982),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1913),
.B(n_23),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2030),
.B(n_23),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2102),
.B(n_24),
.Y(n_2423)
);

INVx4_ASAP7_75t_L g2424 ( 
.A(n_2054),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2025),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1914),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_2037),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_1917),
.B(n_24),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_R g2429 ( 
.A(n_2037),
.B(n_25),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2036),
.Y(n_2430)
);

BUFx4f_ASAP7_75t_L g2431 ( 
.A(n_2132),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_R g2432 ( 
.A(n_2048),
.B(n_26),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_R g2433 ( 
.A(n_2048),
.B(n_26),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_SL g2434 ( 
.A1(n_1873),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2434)
);

AND2x2_ASAP7_75t_SL g2435 ( 
.A(n_1995),
.B(n_27),
.Y(n_2435)
);

INVx2_ASAP7_75t_SL g2436 ( 
.A(n_1921),
.Y(n_2436)
);

A2O1A1Ixp33_ASAP7_75t_L g2437 ( 
.A1(n_1985),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_2437)
);

AOI22xp33_ASAP7_75t_L g2438 ( 
.A1(n_2031),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2438)
);

NAND2xp33_ASAP7_75t_SL g2439 ( 
.A(n_2135),
.B(n_29),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2049),
.Y(n_2440)
);

AOI22xp5_ASAP7_75t_SL g2441 ( 
.A1(n_2033),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2441)
);

INVx1_ASAP7_75t_SL g2442 ( 
.A(n_2080),
.Y(n_2442)
);

INVx2_ASAP7_75t_SL g2443 ( 
.A(n_1959),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1873),
.Y(n_2444)
);

HB1xp67_ASAP7_75t_L g2445 ( 
.A(n_2049),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2022),
.B(n_31),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_1882),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2026),
.B(n_31),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_1882),
.Y(n_2449)
);

INVx5_ASAP7_75t_L g2450 ( 
.A(n_2039),
.Y(n_2450)
);

INVx5_ASAP7_75t_L g2451 ( 
.A(n_2040),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2135),
.B(n_33),
.Y(n_2452)
);

BUFx3_ASAP7_75t_L g2453 ( 
.A(n_2070),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2017),
.B(n_32),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2029),
.B(n_33),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1987),
.Y(n_2456)
);

XNOR2x1_ASAP7_75t_L g2457 ( 
.A(n_1940),
.B(n_35),
.Y(n_2457)
);

INVx1_ASAP7_75t_SL g2458 ( 
.A(n_2080),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2029),
.B(n_34),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_1992),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2126),
.Y(n_2461)
);

CKINVDCx20_ASAP7_75t_R g2462 ( 
.A(n_2019),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2050),
.B(n_35),
.Y(n_2463)
);

NOR3xp33_ASAP7_75t_SL g2464 ( 
.A(n_2106),
.B(n_36),
.C(n_37),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2062),
.B(n_37),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2017),
.B(n_2043),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2045),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2062),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2045),
.Y(n_2469)
);

INVx4_ASAP7_75t_L g2470 ( 
.A(n_1891),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2046),
.B(n_36),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2061),
.B(n_1994),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_1962),
.B(n_1974),
.Y(n_2473)
);

NOR3xp33_ASAP7_75t_SL g2474 ( 
.A(n_2107),
.B(n_2113),
.C(n_2073),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2061),
.B(n_36),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_1998),
.B(n_37),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2124),
.Y(n_2477)
);

OR2x6_ASAP7_75t_L g2478 ( 
.A(n_2076),
.B(n_38),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2128),
.B(n_38),
.Y(n_2479)
);

AND2x4_ASAP7_75t_L g2480 ( 
.A(n_2077),
.B(n_2116),
.Y(n_2480)
);

HB1xp67_ASAP7_75t_L g2481 ( 
.A(n_2047),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2047),
.Y(n_2482)
);

INVx4_ASAP7_75t_L g2483 ( 
.A(n_1894),
.Y(n_2483)
);

HB1xp67_ASAP7_75t_L g2484 ( 
.A(n_2137),
.Y(n_2484)
);

AND2x4_ASAP7_75t_L g2485 ( 
.A(n_2125),
.B(n_38),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2088),
.B(n_2081),
.Y(n_2486)
);

AOI211xp5_ASAP7_75t_L g2487 ( 
.A1(n_2095),
.A2(n_2120),
.B(n_2099),
.C(n_2059),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2032),
.B(n_2035),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2140),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_2141),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_1900),
.Y(n_2491)
);

AOI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_1871),
.A2(n_39),
.B(n_40),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_1849),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2018),
.B(n_39),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_1916),
.B(n_41),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_1900),
.Y(n_2496)
);

BUFx2_ASAP7_75t_L g2497 ( 
.A(n_1852),
.Y(n_2497)
);

O2A1O1Ixp5_ASAP7_75t_L g2498 ( 
.A1(n_1867),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_1847),
.Y(n_2499)
);

INVx3_ASAP7_75t_SL g2500 ( 
.A(n_1929),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_1847),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_1871),
.B(n_42),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2060),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_1847),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_1847),
.Y(n_2505)
);

AND2x6_ASAP7_75t_L g2506 ( 
.A(n_1964),
.B(n_43),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_1847),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1847),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2060),
.Y(n_2509)
);

BUFx6f_ASAP7_75t_L g2510 ( 
.A(n_2060),
.Y(n_2510)
);

NOR3xp33_ASAP7_75t_SL g2511 ( 
.A(n_1849),
.B(n_44),
.C(n_45),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_R g2512 ( 
.A(n_1929),
.B(n_44),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_1871),
.B(n_45),
.Y(n_2513)
);

BUFx12f_ASAP7_75t_L g2514 ( 
.A(n_1849),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_1847),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_1878),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2516)
);

CKINVDCx16_ASAP7_75t_R g2517 ( 
.A(n_2069),
.Y(n_2517)
);

HB1xp67_ASAP7_75t_L g2518 ( 
.A(n_1852),
.Y(n_2518)
);

AOI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_1871),
.A2(n_46),
.B(n_47),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_1871),
.B(n_47),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_1900),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_1847),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_1871),
.B(n_48),
.Y(n_2523)
);

INVx4_ASAP7_75t_L g2524 ( 
.A(n_1929),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_1847),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_1852),
.B(n_49),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_1852),
.B(n_49),
.Y(n_2527)
);

INVx5_ASAP7_75t_L g2528 ( 
.A(n_1929),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1847),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_1929),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2060),
.Y(n_2531)
);

INVxp67_ASAP7_75t_SL g2532 ( 
.A(n_1852),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1847),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1847),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_1847),
.Y(n_2535)
);

AND2x4_ASAP7_75t_L g2536 ( 
.A(n_2018),
.B(n_48),
.Y(n_2536)
);

INVx4_ASAP7_75t_L g2537 ( 
.A(n_1929),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_1852),
.B(n_51),
.Y(n_2538)
);

AOI22x1_ASAP7_75t_L g2539 ( 
.A1(n_2071),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2539)
);

AOI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_1916),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_2018),
.B(n_50),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_1916),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_1871),
.B(n_53),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_1847),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2060),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_1871),
.B(n_54),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_1847),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_1852),
.B(n_54),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_1847),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_R g2550 ( 
.A(n_1929),
.B(n_55),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_1847),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_1847),
.Y(n_2552)
);

AOI22xp33_ASAP7_75t_L g2553 ( 
.A1(n_1878),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_1929),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_1916),
.B(n_56),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_1929),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_1852),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_1852),
.B(n_57),
.Y(n_2558)
);

BUFx2_ASAP7_75t_L g2559 ( 
.A(n_1852),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_1852),
.B(n_56),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_1852),
.B(n_58),
.Y(n_2561)
);

BUFx3_ASAP7_75t_L g2562 ( 
.A(n_1929),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_1871),
.B(n_59),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_1878),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_1900),
.Y(n_2565)
);

BUFx10_ASAP7_75t_L g2566 ( 
.A(n_1970),
.Y(n_2566)
);

INVx5_ASAP7_75t_L g2567 ( 
.A(n_1929),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_1871),
.B(n_60),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_1847),
.Y(n_2569)
);

BUFx3_ASAP7_75t_L g2570 ( 
.A(n_1929),
.Y(n_2570)
);

OAI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_1865),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_R g2572 ( 
.A(n_1929),
.B(n_62),
.Y(n_2572)
);

BUFx2_ASAP7_75t_L g2573 ( 
.A(n_1852),
.Y(n_2573)
);

AOI22xp33_ASAP7_75t_L g2574 ( 
.A1(n_1878),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2574)
);

NAND3xp33_ASAP7_75t_SL g2575 ( 
.A(n_2127),
.B(n_63),
.C(n_64),
.Y(n_2575)
);

OR2x6_ASAP7_75t_L g2576 ( 
.A(n_1929),
.B(n_63),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_1852),
.B(n_64),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_1847),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_R g2579 ( 
.A(n_1929),
.B(n_65),
.Y(n_2579)
);

AO21x2_ASAP7_75t_L g2580 ( 
.A1(n_2071),
.A2(n_65),
.B(n_66),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_1849),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_1847),
.Y(n_2582)
);

BUFx10_ASAP7_75t_L g2583 ( 
.A(n_1970),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2488),
.A2(n_67),
.B(n_68),
.Y(n_2584)
);

OAI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2498),
.A2(n_67),
.B(n_69),
.Y(n_2585)
);

AOI221xp5_ASAP7_75t_L g2586 ( 
.A1(n_2196),
.A2(n_70),
.B1(n_67),
.B2(n_69),
.C(n_71),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2199),
.B(n_69),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2532),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2532),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2145),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2528),
.Y(n_2591)
);

OAI21x1_ASAP7_75t_L g2592 ( 
.A1(n_2247),
.A2(n_70),
.B(n_71),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2457),
.B(n_72),
.Y(n_2593)
);

BUFx6f_ASAP7_75t_L g2594 ( 
.A(n_2528),
.Y(n_2594)
);

OAI21x1_ASAP7_75t_L g2595 ( 
.A1(n_2281),
.A2(n_72),
.B(n_73),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2289),
.B(n_73),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2488),
.A2(n_73),
.B(n_74),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2289),
.B(n_74),
.Y(n_2598)
);

BUFx2_ASAP7_75t_L g2599 ( 
.A(n_2576),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2528),
.Y(n_2600)
);

OAI21x1_ASAP7_75t_L g2601 ( 
.A1(n_2281),
.A2(n_74),
.B(n_75),
.Y(n_2601)
);

OAI21x1_ASAP7_75t_L g2602 ( 
.A1(n_2418),
.A2(n_75),
.B(n_76),
.Y(n_2602)
);

AO31x2_ASAP7_75t_L g2603 ( 
.A1(n_2155),
.A2(n_79),
.A3(n_77),
.B(n_78),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2206),
.B(n_78),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2214),
.B(n_79),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2444),
.B(n_80),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2472),
.A2(n_81),
.B(n_82),
.Y(n_2607)
);

AND2x6_ASAP7_75t_L g2608 ( 
.A(n_2230),
.B(n_83),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_SL g2609 ( 
.A(n_2255),
.B(n_85),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2557),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2447),
.B(n_84),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2151),
.Y(n_2612)
);

AOI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2472),
.A2(n_84),
.B(n_86),
.Y(n_2613)
);

AOI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2486),
.A2(n_84),
.B(n_87),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2486),
.A2(n_88),
.B(n_89),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2528),
.B(n_88),
.Y(n_2616)
);

OAI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2498),
.A2(n_90),
.B(n_91),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_2567),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2449),
.B(n_90),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2323),
.B(n_91),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2255),
.B(n_92),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2557),
.B(n_92),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2156),
.Y(n_2623)
);

OAI21x1_ASAP7_75t_SL g2624 ( 
.A1(n_2320),
.A2(n_93),
.B(n_94),
.Y(n_2624)
);

OAI21xp33_ASAP7_75t_L g2625 ( 
.A1(n_2355),
.A2(n_95),
.B(n_96),
.Y(n_2625)
);

NAND2xp33_ASAP7_75t_L g2626 ( 
.A(n_2567),
.B(n_776),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2332),
.B(n_2333),
.Y(n_2627)
);

OAI21x1_ASAP7_75t_L g2628 ( 
.A1(n_2211),
.A2(n_2272),
.B(n_2225),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2514),
.Y(n_2629)
);

OAI21xp5_ASAP7_75t_L g2630 ( 
.A1(n_2146),
.A2(n_95),
.B(n_96),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2146),
.A2(n_97),
.B(n_98),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2211),
.A2(n_97),
.B(n_99),
.Y(n_2632)
);

NAND2x1p5_ASAP7_75t_L g2633 ( 
.A(n_2567),
.B(n_100),
.Y(n_2633)
);

OAI21x1_ASAP7_75t_L g2634 ( 
.A1(n_2225),
.A2(n_100),
.B(n_101),
.Y(n_2634)
);

INVx4_ASAP7_75t_L g2635 ( 
.A(n_2567),
.Y(n_2635)
);

NAND3xp33_ASAP7_75t_L g2636 ( 
.A(n_2402),
.B(n_101),
.C(n_102),
.Y(n_2636)
);

AOI211x1_ASAP7_75t_L g2637 ( 
.A1(n_2526),
.A2(n_2538),
.B(n_2558),
.C(n_2527),
.Y(n_2637)
);

AO22x2_ASAP7_75t_L g2638 ( 
.A1(n_2240),
.A2(n_2236),
.B1(n_2575),
.B2(n_2230),
.Y(n_2638)
);

AOI21xp33_ASAP7_75t_L g2639 ( 
.A1(n_2419),
.A2(n_2386),
.B(n_2383),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2336),
.B(n_102),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2343),
.B(n_103),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2350),
.B(n_103),
.Y(n_2642)
);

CKINVDCx20_ASAP7_75t_R g2643 ( 
.A(n_2500),
.Y(n_2643)
);

OAI21x1_ASAP7_75t_L g2644 ( 
.A1(n_2272),
.A2(n_104),
.B(n_105),
.Y(n_2644)
);

OAI21x1_ASAP7_75t_L g2645 ( 
.A1(n_2165),
.A2(n_104),
.B(n_106),
.Y(n_2645)
);

AOI211x1_ASAP7_75t_L g2646 ( 
.A1(n_2465),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2646)
);

AOI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2152),
.A2(n_107),
.B(n_109),
.Y(n_2647)
);

AO31x2_ASAP7_75t_L g2648 ( 
.A1(n_2571),
.A2(n_111),
.A3(n_109),
.B(n_110),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2518),
.B(n_110),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2159),
.Y(n_2650)
);

O2A1O1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2177),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_2651)
);

OA21x2_ASAP7_75t_L g2652 ( 
.A1(n_2539),
.A2(n_112),
.B(n_113),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2154),
.Y(n_2653)
);

OA21x2_ASAP7_75t_L g2654 ( 
.A1(n_2446),
.A2(n_116),
.B(n_117),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2297),
.B(n_2300),
.Y(n_2655)
);

BUFx12f_ASAP7_75t_L g2656 ( 
.A(n_2192),
.Y(n_2656)
);

OAI21x1_ASAP7_75t_L g2657 ( 
.A1(n_2165),
.A2(n_116),
.B(n_117),
.Y(n_2657)
);

CKINVDCx6p67_ASAP7_75t_R g2658 ( 
.A(n_2207),
.Y(n_2658)
);

NAND3xp33_ASAP7_75t_SL g2659 ( 
.A(n_2512),
.B(n_118),
.C(n_119),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2468),
.B(n_118),
.Y(n_2660)
);

OAI21x1_ASAP7_75t_L g2661 ( 
.A1(n_2185),
.A2(n_119),
.B(n_120),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2307),
.B(n_120),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2147),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2390),
.B(n_121),
.Y(n_2664)
);

BUFx3_ASAP7_75t_L g2665 ( 
.A(n_2270),
.Y(n_2665)
);

OAI21x1_ASAP7_75t_L g2666 ( 
.A1(n_2185),
.A2(n_121),
.B(n_122),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2154),
.B(n_123),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_2147),
.Y(n_2668)
);

NAND3x1_ASAP7_75t_L g2669 ( 
.A(n_2495),
.B(n_123),
.C(n_124),
.Y(n_2669)
);

OR2x2_ASAP7_75t_L g2670 ( 
.A(n_2254),
.B(n_125),
.Y(n_2670)
);

OAI21x1_ASAP7_75t_L g2671 ( 
.A1(n_2491),
.A2(n_126),
.B(n_128),
.Y(n_2671)
);

OAI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2152),
.A2(n_126),
.B(n_128),
.Y(n_2672)
);

OAI21xp5_ASAP7_75t_L g2673 ( 
.A1(n_2394),
.A2(n_129),
.B(n_130),
.Y(n_2673)
);

A2O1A1Ixp33_ASAP7_75t_L g2674 ( 
.A1(n_2487),
.A2(n_134),
.B(n_129),
.C(n_133),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2171),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2308),
.B(n_133),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2147),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_SL g2678 ( 
.A(n_2238),
.B(n_134),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2518),
.B(n_135),
.Y(n_2679)
);

OAI21x1_ASAP7_75t_SL g2680 ( 
.A1(n_2320),
.A2(n_2339),
.B(n_2338),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2440),
.B(n_2445),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2238),
.B(n_2246),
.Y(n_2682)
);

INVx2_ASAP7_75t_SL g2683 ( 
.A(n_2197),
.Y(n_2683)
);

O2A1O1Ixp5_ASAP7_75t_L g2684 ( 
.A1(n_2282),
.A2(n_140),
.B(n_137),
.C(n_138),
.Y(n_2684)
);

AOI21xp33_ASAP7_75t_L g2685 ( 
.A1(n_2383),
.A2(n_138),
.B(n_140),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2440),
.B(n_141),
.Y(n_2686)
);

OAI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2491),
.A2(n_141),
.B(n_142),
.Y(n_2687)
);

AOI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2355),
.A2(n_2301),
.B(n_2373),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2445),
.B(n_2426),
.Y(n_2689)
);

OAI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2394),
.A2(n_142),
.B(n_143),
.Y(n_2690)
);

INVx3_ASAP7_75t_L g2691 ( 
.A(n_2167),
.Y(n_2691)
);

NOR2xp67_ASAP7_75t_L g2692 ( 
.A(n_2167),
.B(n_143),
.Y(n_2692)
);

AO21x1_ASAP7_75t_L g2693 ( 
.A1(n_2571),
.A2(n_144),
.B(n_145),
.Y(n_2693)
);

AOI21x1_ASAP7_75t_L g2694 ( 
.A1(n_2375),
.A2(n_146),
.B(n_148),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2524),
.B(n_146),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2275),
.B(n_149),
.Y(n_2696)
);

OAI21x1_ASAP7_75t_L g2697 ( 
.A1(n_2496),
.A2(n_149),
.B(n_150),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2497),
.B(n_150),
.Y(n_2698)
);

OAI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_2576),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2180),
.Y(n_2700)
);

AOI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2373),
.A2(n_152),
.B(n_153),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2303),
.B(n_154),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2384),
.B(n_156),
.Y(n_2703)
);

OAI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2502),
.A2(n_157),
.B(n_158),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2236),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_2705)
);

OAI21x1_ASAP7_75t_L g2706 ( 
.A1(n_2496),
.A2(n_160),
.B(n_162),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2435),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2388),
.B(n_163),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2193),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2395),
.B(n_164),
.Y(n_2710)
);

AO31x2_ASAP7_75t_L g2711 ( 
.A1(n_2386),
.A2(n_167),
.A3(n_165),
.B(n_166),
.Y(n_2711)
);

OAI22xp5_ASAP7_75t_L g2712 ( 
.A1(n_2412),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_2712)
);

OAI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_2502),
.A2(n_168),
.B(n_169),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2409),
.A2(n_169),
.B(n_170),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2397),
.B(n_172),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2501),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2404),
.B(n_173),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2406),
.B(n_174),
.Y(n_2718)
);

BUFx2_ASAP7_75t_L g2719 ( 
.A(n_2576),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2466),
.A2(n_177),
.B(n_178),
.Y(n_2720)
);

OAI21x1_ASAP7_75t_L g2721 ( 
.A1(n_2521),
.A2(n_178),
.B(n_179),
.Y(n_2721)
);

OA21x2_ASAP7_75t_L g2722 ( 
.A1(n_2446),
.A2(n_179),
.B(n_181),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2416),
.B(n_181),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2420),
.B(n_182),
.Y(n_2724)
);

OAI21x1_ASAP7_75t_L g2725 ( 
.A1(n_2565),
.A2(n_182),
.B(n_183),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2513),
.A2(n_184),
.B(n_185),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2218),
.B(n_184),
.Y(n_2727)
);

OAI21x1_ASAP7_75t_L g2728 ( 
.A1(n_2565),
.A2(n_185),
.B(n_186),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2220),
.B(n_186),
.Y(n_2729)
);

AOI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2466),
.A2(n_187),
.B(n_188),
.Y(n_2730)
);

OAI21x1_ASAP7_75t_L g2731 ( 
.A1(n_2315),
.A2(n_188),
.B(n_189),
.Y(n_2731)
);

INVx2_ASAP7_75t_SL g2732 ( 
.A(n_2556),
.Y(n_2732)
);

AOI21xp33_ASAP7_75t_L g2733 ( 
.A1(n_2177),
.A2(n_190),
.B(n_191),
.Y(n_2733)
);

AOI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2183),
.A2(n_191),
.B(n_192),
.Y(n_2734)
);

OAI21x1_ASAP7_75t_L g2735 ( 
.A1(n_2315),
.A2(n_193),
.B(n_194),
.Y(n_2735)
);

OAI21x1_ASAP7_75t_L g2736 ( 
.A1(n_2292),
.A2(n_2366),
.B(n_2269),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_SL g2737 ( 
.A1(n_2434),
.A2(n_193),
.B(n_194),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2231),
.B(n_195),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2249),
.B(n_197),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2569),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2251),
.B(n_197),
.Y(n_2741)
);

BUFx10_ASAP7_75t_L g2742 ( 
.A(n_2201),
.Y(n_2742)
);

NAND2x1p5_ASAP7_75t_L g2743 ( 
.A(n_2524),
.B(n_198),
.Y(n_2743)
);

OA21x2_ASAP7_75t_L g2744 ( 
.A1(n_2455),
.A2(n_198),
.B(n_199),
.Y(n_2744)
);

INVx4_ASAP7_75t_L g2745 ( 
.A(n_2537),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2363),
.B(n_202),
.Y(n_2746)
);

OAI21xp33_ASAP7_75t_L g2747 ( 
.A1(n_2341),
.A2(n_202),
.B(n_203),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2559),
.B(n_2573),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2253),
.B(n_2259),
.Y(n_2749)
);

BUFx6f_ASAP7_75t_L g2750 ( 
.A(n_2150),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2262),
.B(n_2264),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2284),
.B(n_203),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2456),
.B(n_204),
.Y(n_2753)
);

AO31x2_ASAP7_75t_L g2754 ( 
.A1(n_2455),
.A2(n_209),
.A3(n_204),
.B(n_207),
.Y(n_2754)
);

AOI221x1_ASAP7_75t_L g2755 ( 
.A1(n_2575),
.A2(n_211),
.B1(n_207),
.B2(n_210),
.C(n_212),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2578),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2363),
.B(n_211),
.Y(n_2757)
);

AND2x6_ASAP7_75t_L g2758 ( 
.A(n_2494),
.B(n_213),
.Y(n_2758)
);

OAI21x1_ASAP7_75t_L g2759 ( 
.A1(n_2292),
.A2(n_213),
.B(n_214),
.Y(n_2759)
);

OAI21x1_ASAP7_75t_L g2760 ( 
.A1(n_2366),
.A2(n_214),
.B(n_215),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2513),
.A2(n_215),
.B(n_216),
.Y(n_2761)
);

A2O1A1Ixp33_ASAP7_75t_L g2762 ( 
.A1(n_2439),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2142),
.Y(n_2763)
);

AOI21x1_ASAP7_75t_L g2764 ( 
.A1(n_2375),
.A2(n_217),
.B(n_218),
.Y(n_2764)
);

OR2x2_ASAP7_75t_L g2765 ( 
.A(n_2233),
.B(n_219),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2537),
.Y(n_2766)
);

OAI21x1_ASAP7_75t_L g2767 ( 
.A1(n_2459),
.A2(n_220),
.B(n_222),
.Y(n_2767)
);

AOI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2520),
.A2(n_220),
.B(n_223),
.Y(n_2768)
);

NOR2xp33_ASAP7_75t_L g2769 ( 
.A(n_2387),
.B(n_223),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2520),
.A2(n_224),
.B(n_226),
.Y(n_2770)
);

OAI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2523),
.A2(n_224),
.B(n_226),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2150),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2467),
.B(n_227),
.Y(n_2773)
);

OAI21x1_ASAP7_75t_L g2774 ( 
.A1(n_2459),
.A2(n_227),
.B(n_228),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2346),
.B(n_228),
.Y(n_2775)
);

AOI221x1_ASAP7_75t_L g2776 ( 
.A1(n_2240),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.C(n_232),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2460),
.B(n_231),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2358),
.B(n_233),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2191),
.B(n_2432),
.Y(n_2779)
);

OAI21x1_ASAP7_75t_L g2780 ( 
.A1(n_2401),
.A2(n_234),
.B(n_235),
.Y(n_2780)
);

O2A1O1Ixp5_ASAP7_75t_L g2781 ( 
.A1(n_2321),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2143),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_2215),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_SL g2784 ( 
.A(n_2222),
.B(n_238),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2310),
.B(n_239),
.Y(n_2785)
);

AO31x2_ASAP7_75t_L g2786 ( 
.A1(n_2288),
.A2(n_241),
.A3(n_239),
.B(n_240),
.Y(n_2786)
);

A2O1A1Ixp33_ASAP7_75t_L g2787 ( 
.A1(n_2523),
.A2(n_243),
.B(n_240),
.C(n_242),
.Y(n_2787)
);

CKINVDCx11_ASAP7_75t_R g2788 ( 
.A(n_2200),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2543),
.A2(n_243),
.B(n_244),
.Y(n_2789)
);

AND3x4_ASAP7_75t_L g2790 ( 
.A(n_2511),
.B(n_2153),
.C(n_2160),
.Y(n_2790)
);

NAND3x1_ASAP7_75t_L g2791 ( 
.A(n_2555),
.B(n_247),
.C(n_248),
.Y(n_2791)
);

O2A1O1Ixp33_ASAP7_75t_L g2792 ( 
.A1(n_2437),
.A2(n_253),
.B(n_249),
.C(n_250),
.Y(n_2792)
);

OAI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2543),
.A2(n_249),
.B(n_250),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2270),
.Y(n_2794)
);

AOI21xp5_ASAP7_75t_L g2795 ( 
.A1(n_2546),
.A2(n_254),
.B(n_255),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_SL g2796 ( 
.A(n_2298),
.B(n_255),
.Y(n_2796)
);

INVx4_ASAP7_75t_SL g2797 ( 
.A(n_2506),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2311),
.B(n_258),
.Y(n_2798)
);

OAI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2546),
.A2(n_259),
.B(n_260),
.Y(n_2799)
);

OA22x2_ASAP7_75t_L g2800 ( 
.A1(n_2222),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_2800)
);

AO31x2_ASAP7_75t_L g2801 ( 
.A1(n_2288),
.A2(n_265),
.A3(n_261),
.B(n_263),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2191),
.B(n_263),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2433),
.B(n_265),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2563),
.A2(n_266),
.B(n_269),
.Y(n_2804)
);

AO31x2_ASAP7_75t_L g2805 ( 
.A1(n_2492),
.A2(n_273),
.A3(n_270),
.B(n_271),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2314),
.B(n_270),
.Y(n_2806)
);

OAI21x1_ASAP7_75t_L g2807 ( 
.A1(n_2273),
.A2(n_271),
.B(n_273),
.Y(n_2807)
);

AOI22xp5_ASAP7_75t_SL g2808 ( 
.A1(n_2517),
.A2(n_2506),
.B1(n_2234),
.B2(n_2250),
.Y(n_2808)
);

AOI221xp5_ASAP7_75t_SL g2809 ( 
.A1(n_2492),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_2809)
);

BUFx2_ASAP7_75t_L g2810 ( 
.A(n_2550),
.Y(n_2810)
);

AO22x2_ASAP7_75t_L g2811 ( 
.A1(n_2494),
.A2(n_2541),
.B1(n_2536),
.B2(n_2248),
.Y(n_2811)
);

A2O1A1Ixp33_ASAP7_75t_L g2812 ( 
.A1(n_2563),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2568),
.A2(n_2402),
.B1(n_2434),
.B2(n_2481),
.Y(n_2813)
);

OAI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2568),
.A2(n_278),
.B(n_279),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2469),
.B(n_278),
.Y(n_2815)
);

CKINVDCx20_ASAP7_75t_R g2816 ( 
.A(n_2572),
.Y(n_2816)
);

A2O1A1Ixp33_ASAP7_75t_L g2817 ( 
.A1(n_2519),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2817)
);

BUFx6f_ASAP7_75t_L g2818 ( 
.A(n_2150),
.Y(n_2818)
);

OAI21x1_ASAP7_75t_L g2819 ( 
.A1(n_2273),
.A2(n_280),
.B(n_281),
.Y(n_2819)
);

OAI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2519),
.A2(n_282),
.B(n_283),
.Y(n_2820)
);

HB1xp67_ASAP7_75t_L g2821 ( 
.A(n_2298),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2482),
.B(n_282),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2148),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_SL g2824 ( 
.A1(n_2375),
.A2(n_283),
.B(n_284),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2149),
.B(n_284),
.Y(n_2825)
);

OAI22x1_ASAP7_75t_L g2826 ( 
.A1(n_2250),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_2826)
);

AO31x2_ASAP7_75t_L g2827 ( 
.A1(n_2327),
.A2(n_288),
.A3(n_285),
.B(n_287),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_2579),
.B(n_289),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2405),
.A2(n_289),
.B(n_290),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2161),
.B(n_290),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2170),
.B(n_2172),
.Y(n_2831)
);

INVx3_ASAP7_75t_L g2832 ( 
.A(n_2173),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2562),
.B(n_291),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2179),
.B(n_291),
.Y(n_2834)
);

AOI221xp5_ASAP7_75t_L g2835 ( 
.A1(n_2257),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.C(n_295),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2187),
.B(n_293),
.Y(n_2836)
);

OAI21x1_ASAP7_75t_L g2837 ( 
.A1(n_2278),
.A2(n_294),
.B(n_295),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2256),
.B(n_297),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2189),
.B(n_2499),
.Y(n_2839)
);

OAI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2367),
.A2(n_300),
.B(n_301),
.Y(n_2840)
);

OAI21x1_ASAP7_75t_L g2841 ( 
.A1(n_2278),
.A2(n_300),
.B(n_301),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2504),
.B(n_2505),
.Y(n_2842)
);

OAI21x1_ASAP7_75t_L g2843 ( 
.A1(n_2302),
.A2(n_304),
.B(n_307),
.Y(n_2843)
);

INVx2_ASAP7_75t_SL g2844 ( 
.A(n_2570),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2507),
.B(n_307),
.Y(n_2845)
);

AOI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2405),
.A2(n_308),
.B(n_309),
.Y(n_2846)
);

OR2x2_ASAP7_75t_L g2847 ( 
.A(n_2347),
.B(n_310),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2258),
.B(n_311),
.Y(n_2848)
);

A2O1A1Ixp33_ASAP7_75t_L g2849 ( 
.A1(n_2329),
.A2(n_2335),
.B(n_2351),
.C(n_2407),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2508),
.B(n_311),
.Y(n_2850)
);

OAI21x1_ASAP7_75t_L g2851 ( 
.A1(n_2302),
.A2(n_312),
.B(n_313),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2515),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_SL g2853 ( 
.A1(n_2169),
.A2(n_312),
.B(n_313),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2522),
.B(n_314),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2407),
.A2(n_315),
.B(n_316),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2525),
.B(n_316),
.Y(n_2856)
);

HB1xp67_ASAP7_75t_L g2857 ( 
.A(n_2536),
.Y(n_2857)
);

AO22x2_ASAP7_75t_L g2858 ( 
.A1(n_2541),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2326),
.B(n_317),
.Y(n_2859)
);

AOI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2417),
.A2(n_318),
.B(n_320),
.Y(n_2860)
);

OAI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2367),
.A2(n_322),
.B(n_323),
.Y(n_2861)
);

INVx1_ASAP7_75t_SL g2862 ( 
.A(n_2178),
.Y(n_2862)
);

NAND3xp33_ASAP7_75t_SL g2863 ( 
.A(n_2312),
.B(n_322),
.C(n_323),
.Y(n_2863)
);

OAI21x1_ASAP7_75t_L g2864 ( 
.A1(n_2362),
.A2(n_324),
.B(n_325),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2529),
.B(n_326),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2533),
.B(n_329),
.Y(n_2866)
);

CKINVDCx11_ASAP7_75t_R g2867 ( 
.A(n_2163),
.Y(n_2867)
);

OAI21xp33_ASAP7_75t_L g2868 ( 
.A1(n_2305),
.A2(n_330),
.B(n_331),
.Y(n_2868)
);

AOI21xp5_ASAP7_75t_SL g2869 ( 
.A1(n_2169),
.A2(n_330),
.B(n_332),
.Y(n_2869)
);

O2A1O1Ixp33_ASAP7_75t_SL g2870 ( 
.A1(n_2271),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_2870)
);

OAI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2364),
.A2(n_333),
.B(n_334),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2328),
.B(n_335),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2166),
.B(n_336),
.Y(n_2873)
);

AO31x2_ASAP7_75t_L g2874 ( 
.A1(n_2335),
.A2(n_338),
.A3(n_336),
.B(n_337),
.Y(n_2874)
);

OAI21xp33_ASAP7_75t_L g2875 ( 
.A1(n_2305),
.A2(n_2438),
.B(n_2371),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2534),
.B(n_2535),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_2215),
.Y(n_2877)
);

AO21x1_ASAP7_75t_L g2878 ( 
.A1(n_2452),
.A2(n_337),
.B(n_338),
.Y(n_2878)
);

AO21x2_ASAP7_75t_L g2879 ( 
.A1(n_2580),
.A2(n_339),
.B(n_340),
.Y(n_2879)
);

BUFx5_ASAP7_75t_L g2880 ( 
.A(n_2190),
.Y(n_2880)
);

INVx3_ASAP7_75t_L g2881 ( 
.A(n_2173),
.Y(n_2881)
);

O2A1O1Ixp5_ASAP7_75t_L g2882 ( 
.A1(n_2348),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_2882)
);

INVx6_ASAP7_75t_L g2883 ( 
.A(n_2163),
.Y(n_2883)
);

AO31x2_ASAP7_75t_L g2884 ( 
.A1(n_2351),
.A2(n_345),
.A3(n_343),
.B(n_344),
.Y(n_2884)
);

OR2x2_ASAP7_75t_L g2885 ( 
.A(n_2331),
.B(n_345),
.Y(n_2885)
);

OAI21xp5_ASAP7_75t_L g2886 ( 
.A1(n_2417),
.A2(n_346),
.B(n_347),
.Y(n_2886)
);

OAI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2421),
.A2(n_348),
.B(n_349),
.Y(n_2887)
);

INVx2_ASAP7_75t_SL g2888 ( 
.A(n_2221),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2544),
.B(n_348),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2429),
.B(n_349),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2547),
.B(n_350),
.Y(n_2891)
);

NAND3x1_ASAP7_75t_L g2892 ( 
.A(n_2540),
.B(n_351),
.C(n_353),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2549),
.Y(n_2893)
);

OAI21x1_ASAP7_75t_L g2894 ( 
.A1(n_2372),
.A2(n_354),
.B(n_355),
.Y(n_2894)
);

A2O1A1Ixp33_ASAP7_75t_L g2895 ( 
.A1(n_2428),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_2895)
);

OAI21x1_ASAP7_75t_L g2896 ( 
.A1(n_2379),
.A2(n_357),
.B(n_358),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2551),
.B(n_357),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2552),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2582),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2473),
.B(n_2481),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2221),
.Y(n_2901)
);

INVx2_ASAP7_75t_SL g2902 ( 
.A(n_2221),
.Y(n_2902)
);

BUFx2_ASAP7_75t_L g2903 ( 
.A(n_2316),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2356),
.B(n_361),
.Y(n_2904)
);

O2A1O1Ixp5_ASAP7_75t_L g2905 ( 
.A1(n_2413),
.A2(n_365),
.B(n_362),
.C(n_363),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2389),
.B(n_371),
.Y(n_2906)
);

OAI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2475),
.A2(n_371),
.B(n_372),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2184),
.B(n_373),
.Y(n_2908)
);

AND3x4_ASAP7_75t_L g2909 ( 
.A(n_2511),
.B(n_373),
.C(n_374),
.Y(n_2909)
);

AO31x2_ASAP7_75t_L g2910 ( 
.A1(n_2338),
.A2(n_376),
.A3(n_374),
.B(n_375),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2360),
.B(n_375),
.Y(n_2911)
);

OAI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2454),
.A2(n_2476),
.B(n_2403),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2168),
.B(n_2182),
.Y(n_2913)
);

HB1xp67_ASAP7_75t_L g2914 ( 
.A(n_2223),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_2392),
.B(n_377),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2168),
.B(n_378),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2182),
.B(n_379),
.Y(n_2917)
);

OAI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2476),
.A2(n_380),
.B(n_381),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2144),
.B(n_382),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2198),
.B(n_383),
.Y(n_2920)
);

AOI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2542),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_2921)
);

OAI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2237),
.A2(n_2322),
.B1(n_2371),
.B2(n_2353),
.Y(n_2922)
);

INVx1_ASAP7_75t_SL g2923 ( 
.A(n_2359),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2198),
.B(n_385),
.Y(n_2924)
);

OAI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2403),
.A2(n_387),
.B(n_390),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2205),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2370),
.Y(n_2927)
);

OA21x2_ASAP7_75t_L g2928 ( 
.A1(n_2344),
.A2(n_393),
.B(n_394),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2393),
.B(n_395),
.Y(n_2929)
);

AOI21x1_ASAP7_75t_L g2930 ( 
.A1(n_2427),
.A2(n_400),
.B(n_401),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2374),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2489),
.B(n_2377),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2322),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2933)
);

OAI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2352),
.A2(n_402),
.B(n_403),
.Y(n_2934)
);

OAI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2463),
.A2(n_404),
.B(n_405),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2263),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2422),
.B(n_405),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2306),
.B(n_2354),
.Y(n_2938)
);

OAI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2463),
.A2(n_406),
.B(n_407),
.Y(n_2939)
);

INVx1_ASAP7_75t_SL g2940 ( 
.A(n_2285),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2248),
.B(n_407),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2244),
.B(n_2245),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2287),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2244),
.B(n_408),
.Y(n_2944)
);

INVx3_ASAP7_75t_L g2945 ( 
.A(n_2176),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2195),
.A2(n_408),
.B(n_409),
.Y(n_2946)
);

AO21x2_ASAP7_75t_L g2947 ( 
.A1(n_2313),
.A2(n_409),
.B(n_410),
.Y(n_2947)
);

INVx3_ASAP7_75t_L g2948 ( 
.A(n_2176),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2245),
.B(n_410),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2503),
.A2(n_2510),
.B(n_2509),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2239),
.Y(n_2951)
);

OAI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2195),
.A2(n_412),
.B(n_413),
.Y(n_2952)
);

OR2x2_ASAP7_75t_L g2953 ( 
.A(n_2380),
.B(n_413),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2317),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2324),
.Y(n_2955)
);

OA21x2_ASAP7_75t_L g2956 ( 
.A1(n_2342),
.A2(n_416),
.B(n_417),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2509),
.A2(n_416),
.B(n_418),
.Y(n_2957)
);

AO22x2_ASAP7_75t_L g2958 ( 
.A1(n_2239),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_SL g2959 ( 
.A1(n_2334),
.A2(n_2441),
.B1(n_2232),
.B2(n_2223),
.Y(n_2959)
);

AO31x2_ASAP7_75t_L g2960 ( 
.A1(n_2339),
.A2(n_422),
.A3(n_419),
.B(n_421),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2548),
.Y(n_2961)
);

CKINVDCx20_ASAP7_75t_R g2962 ( 
.A(n_2643),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2842),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2688),
.B(n_2427),
.Y(n_2964)
);

INVx6_ASAP7_75t_L g2965 ( 
.A(n_2745),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_SL g2966 ( 
.A1(n_2705),
.A2(n_2325),
.B(n_2234),
.Y(n_2966)
);

OA21x2_ASAP7_75t_L g2967 ( 
.A1(n_2639),
.A2(n_2330),
.B(n_2464),
.Y(n_2967)
);

NOR2x1_ASAP7_75t_SL g2968 ( 
.A(n_2635),
.B(n_2478),
.Y(n_2968)
);

OAI21x1_ASAP7_75t_L g2969 ( 
.A1(n_2950),
.A2(n_2304),
.B(n_2299),
.Y(n_2969)
);

AO21x2_ASAP7_75t_L g2970 ( 
.A1(n_2639),
.A2(n_2330),
.B(n_2353),
.Y(n_2970)
);

AND2x4_ASAP7_75t_L g2971 ( 
.A(n_2797),
.B(n_2228),
.Y(n_2971)
);

OR2x2_ASAP7_75t_L g2972 ( 
.A(n_2900),
.B(n_2224),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2842),
.Y(n_2973)
);

OAI21x1_ASAP7_75t_L g2974 ( 
.A1(n_2680),
.A2(n_2592),
.B(n_2628),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2593),
.B(n_2560),
.Y(n_2975)
);

OR2x2_ASAP7_75t_L g2976 ( 
.A(n_2681),
.B(n_2689),
.Y(n_2976)
);

AOI221x1_ASAP7_75t_SL g2977 ( 
.A1(n_2664),
.A2(n_2224),
.B1(n_2398),
.B2(n_2423),
.C(n_2345),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2763),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2779),
.B(n_2561),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2797),
.B(n_2229),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2635),
.Y(n_2981)
);

AND2x4_ASAP7_75t_SL g2982 ( 
.A(n_2745),
.B(n_2566),
.Y(n_2982)
);

OAI21x1_ASAP7_75t_L g2983 ( 
.A1(n_2731),
.A2(n_2531),
.B(n_2510),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2590),
.Y(n_2984)
);

NAND2x1p5_ASAP7_75t_L g2985 ( 
.A(n_2594),
.B(n_2174),
.Y(n_2985)
);

OAI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2849),
.A2(n_2813),
.B(n_2913),
.Y(n_2986)
);

HB1xp67_ASAP7_75t_L g2987 ( 
.A(n_2610),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2591),
.B(n_2227),
.Y(n_2988)
);

HB1xp67_ASAP7_75t_L g2989 ( 
.A(n_2821),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2782),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2594),
.Y(n_2991)
);

INVx1_ASAP7_75t_SL g2992 ( 
.A(n_2923),
.Y(n_2992)
);

BUFx4_ASAP7_75t_R g2993 ( 
.A(n_2665),
.Y(n_2993)
);

NOR2xp33_ASAP7_75t_L g2994 ( 
.A(n_2599),
.B(n_2381),
.Y(n_2994)
);

BUFx2_ASAP7_75t_SL g2995 ( 
.A(n_2794),
.Y(n_2995)
);

BUFx3_ASAP7_75t_L g2996 ( 
.A(n_2788),
.Y(n_2996)
);

INVxp67_ASAP7_75t_SL g2997 ( 
.A(n_2626),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2893),
.Y(n_2998)
);

OAI21x1_ASAP7_75t_L g2999 ( 
.A1(n_2735),
.A2(n_2545),
.B(n_2531),
.Y(n_2999)
);

AOI21x1_ASAP7_75t_L g3000 ( 
.A1(n_2638),
.A2(n_2203),
.B(n_2461),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2623),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2898),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2602),
.A2(n_2545),
.B(n_2531),
.Y(n_3003)
);

OA21x2_ASAP7_75t_L g3004 ( 
.A1(n_2617),
.A2(n_2464),
.B(n_2458),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2617),
.A2(n_2382),
.B(n_2411),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2927),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2931),
.Y(n_3007)
);

AO31x2_ASAP7_75t_L g3008 ( 
.A1(n_2813),
.A2(n_2424),
.A3(n_2414),
.B(n_2448),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2650),
.Y(n_3009)
);

HB1xp67_ASAP7_75t_L g3010 ( 
.A(n_2588),
.Y(n_3010)
);

BUFx2_ASAP7_75t_L g3011 ( 
.A(n_2594),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2912),
.B(n_2309),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2719),
.B(n_2385),
.Y(n_3013)
);

AOI22xp33_ASAP7_75t_SL g3014 ( 
.A1(n_2811),
.A2(n_2506),
.B1(n_2345),
.B2(n_2319),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2938),
.B(n_2477),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2932),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2875),
.A2(n_2478),
.B1(n_2423),
.B2(n_2490),
.Y(n_3017)
);

OAI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2737),
.A2(n_2478),
.B1(n_2319),
.B2(n_2286),
.Y(n_3018)
);

OAI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2737),
.A2(n_2296),
.B1(n_2368),
.B2(n_2442),
.Y(n_3019)
);

OAI21x1_ASAP7_75t_SL g3020 ( 
.A1(n_2705),
.A2(n_2553),
.B(n_2516),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2875),
.A2(n_2490),
.B1(n_2485),
.B2(n_2479),
.Y(n_3021)
);

NAND2xp33_ASAP7_75t_L g3022 ( 
.A(n_2608),
.B(n_2506),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2608),
.A2(n_2490),
.B1(n_2485),
.B2(n_2479),
.Y(n_3023)
);

OAI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2585),
.A2(n_2471),
.B(n_2382),
.Y(n_3024)
);

OAI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2784),
.A2(n_2442),
.B1(n_2458),
.B2(n_2295),
.Y(n_3025)
);

O2A1O1Ixp33_ASAP7_75t_SL g3026 ( 
.A1(n_2707),
.A2(n_2484),
.B(n_2188),
.C(n_2268),
.Y(n_3026)
);

OA21x2_ASAP7_75t_L g3027 ( 
.A1(n_2585),
.A2(n_2361),
.B(n_2309),
.Y(n_3027)
);

OAI22xp5_ASAP7_75t_SL g3028 ( 
.A1(n_2959),
.A2(n_2462),
.B1(n_2574),
.B2(n_2564),
.Y(n_3028)
);

OAI21x1_ASAP7_75t_SL g3029 ( 
.A1(n_2925),
.A2(n_2470),
.B(n_2483),
.Y(n_3029)
);

BUFx8_ASAP7_75t_L g3030 ( 
.A(n_2656),
.Y(n_3030)
);

O2A1O1Ixp33_ASAP7_75t_L g3031 ( 
.A1(n_2712),
.A2(n_2202),
.B(n_2209),
.C(n_2204),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2811),
.B(n_2577),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_SL g3033 ( 
.A1(n_2707),
.A2(n_2190),
.B1(n_2241),
.B2(n_2252),
.Y(n_3033)
);

OAI221xp5_ASAP7_75t_L g3034 ( 
.A1(n_2868),
.A2(n_2265),
.B1(n_2181),
.B2(n_2266),
.C(n_2261),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2675),
.Y(n_3035)
);

OAI21x1_ASAP7_75t_L g3036 ( 
.A1(n_2595),
.A2(n_2601),
.B(n_2780),
.Y(n_3036)
);

BUFx2_ASAP7_75t_SL g3037 ( 
.A(n_2816),
.Y(n_3037)
);

BUFx10_ASAP7_75t_L g3038 ( 
.A(n_2783),
.Y(n_3038)
);

AO21x2_ASAP7_75t_L g3039 ( 
.A1(n_2625),
.A2(n_2188),
.B(n_2261),
.Y(n_3039)
);

OAI21x1_ASAP7_75t_L g3040 ( 
.A1(n_2864),
.A2(n_2337),
.B(n_2357),
.Y(n_3040)
);

OAI21x1_ASAP7_75t_L g3041 ( 
.A1(n_2871),
.A2(n_2337),
.B(n_2391),
.Y(n_3041)
);

NOR2xp33_ASAP7_75t_L g3042 ( 
.A(n_2810),
.B(n_2157),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2756),
.Y(n_3043)
);

BUFx3_ASAP7_75t_L g3044 ( 
.A(n_2903),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2926),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2823),
.Y(n_3046)
);

NOR2x1_ASAP7_75t_R g3047 ( 
.A(n_2867),
.B(n_2493),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2932),
.Y(n_3048)
);

AO21x2_ASAP7_75t_L g3049 ( 
.A1(n_2625),
.A2(n_2280),
.B(n_2277),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2831),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2839),
.Y(n_3051)
);

NAND3xp33_ASAP7_75t_L g3052 ( 
.A(n_2755),
.B(n_2265),
.C(n_2181),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2876),
.Y(n_3053)
);

BUFx6f_ASAP7_75t_L g3054 ( 
.A(n_2600),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2852),
.Y(n_3055)
);

NAND2x1p5_ASAP7_75t_L g3056 ( 
.A(n_2600),
.B(n_2530),
.Y(n_3056)
);

AND2x4_ASAP7_75t_L g3057 ( 
.A(n_2591),
.B(n_2227),
.Y(n_3057)
);

AO21x2_ASAP7_75t_L g3058 ( 
.A1(n_2840),
.A2(n_2280),
.B(n_2277),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2899),
.Y(n_3059)
);

BUFx8_ASAP7_75t_L g3060 ( 
.A(n_2608),
.Y(n_3060)
);

AO21x2_ASAP7_75t_L g3061 ( 
.A1(n_2840),
.A2(n_2291),
.B(n_2204),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2638),
.A2(n_2318),
.B(n_2283),
.Y(n_3062)
);

O2A1O1Ixp33_ASAP7_75t_SL g3063 ( 
.A1(n_2762),
.A2(n_2202),
.B(n_2216),
.C(n_2209),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2636),
.A2(n_2361),
.B1(n_2291),
.B2(n_2276),
.Y(n_3064)
);

OAI21x1_ASAP7_75t_L g3065 ( 
.A1(n_2736),
.A2(n_2337),
.B(n_2391),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2612),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_2790),
.B(n_2396),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2857),
.B(n_2349),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2912),
.B(n_2391),
.Y(n_3069)
);

OAI22xp5_ASAP7_75t_SL g3070 ( 
.A1(n_2909),
.A2(n_2581),
.B1(n_2554),
.B2(n_2295),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2922),
.A2(n_2318),
.B(n_2283),
.Y(n_3071)
);

OAI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2942),
.A2(n_2217),
.B(n_2216),
.Y(n_3072)
);

AOI22xp33_ASAP7_75t_L g3073 ( 
.A1(n_2608),
.A2(n_2480),
.B1(n_2443),
.B2(n_2436),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2700),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2709),
.Y(n_3075)
);

OAI21x1_ASAP7_75t_SL g3076 ( 
.A1(n_2925),
.A2(n_2470),
.B(n_2483),
.Y(n_3076)
);

OR2x2_ASAP7_75t_L g3077 ( 
.A(n_2923),
.B(n_2365),
.Y(n_3077)
);

AO21x2_ASAP7_75t_L g3078 ( 
.A1(n_2861),
.A2(n_2226),
.B(n_2217),
.Y(n_3078)
);

INVx4_ASAP7_75t_L g3079 ( 
.A(n_2618),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2716),
.Y(n_3080)
);

OAI21x1_ASAP7_75t_SL g3081 ( 
.A1(n_2712),
.A2(n_2907),
.B(n_2673),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2748),
.B(n_2162),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2740),
.Y(n_3083)
);

OAI21x1_ASAP7_75t_L g3084 ( 
.A1(n_2767),
.A2(n_2190),
.B(n_2290),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2589),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2936),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_SL g3087 ( 
.A(n_2784),
.B(n_2276),
.Y(n_3087)
);

OAI21x1_ASAP7_75t_L g3088 ( 
.A1(n_2774),
.A2(n_2213),
.B(n_2283),
.Y(n_3088)
);

HB1xp67_ASAP7_75t_L g3089 ( 
.A(n_2914),
.Y(n_3089)
);

NAND2x1p5_ASAP7_75t_L g3090 ( 
.A(n_2618),
.B(n_2194),
.Y(n_3090)
);

OAI21x1_ASAP7_75t_L g3091 ( 
.A1(n_2896),
.A2(n_2340),
.B(n_2318),
.Y(n_3091)
);

OAI21x1_ASAP7_75t_SL g3092 ( 
.A1(n_2907),
.A2(n_2242),
.B(n_2226),
.Y(n_3092)
);

O2A1O1Ixp33_ASAP7_75t_L g3093 ( 
.A1(n_2733),
.A2(n_2242),
.B(n_2243),
.C(n_2294),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2627),
.B(n_2415),
.Y(n_3094)
);

A2O1A1Ixp33_ASAP7_75t_L g3095 ( 
.A1(n_2868),
.A2(n_2186),
.B(n_2164),
.C(n_2175),
.Y(n_3095)
);

OAI21xp33_ASAP7_75t_SL g3096 ( 
.A1(n_2820),
.A2(n_2243),
.B(n_2294),
.Y(n_3096)
);

OAI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2921),
.A2(n_2295),
.B1(n_2369),
.B2(n_2235),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2845),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2627),
.Y(n_3099)
);

OAI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2921),
.A2(n_2295),
.B1(n_2158),
.B2(n_2376),
.Y(n_3100)
);

OAI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2607),
.A2(n_2474),
.B(n_2164),
.Y(n_3101)
);

AO21x2_ASAP7_75t_L g3102 ( 
.A1(n_2861),
.A2(n_2474),
.B(n_2212),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_2940),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2655),
.B(n_2415),
.Y(n_3104)
);

AOI21xp33_ASAP7_75t_SL g3105 ( 
.A1(n_2877),
.A2(n_2260),
.B(n_2210),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2859),
.B(n_2175),
.Y(n_3106)
);

AO21x2_ASAP7_75t_L g3107 ( 
.A1(n_2820),
.A2(n_2212),
.B(n_2194),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2758),
.A2(n_2480),
.B1(n_2378),
.B2(n_2349),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_2872),
.B(n_2160),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2943),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2618),
.B(n_2653),
.Y(n_3111)
);

OAI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2636),
.A2(n_2274),
.B1(n_2450),
.B2(n_2415),
.Y(n_3112)
);

OAI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2584),
.A2(n_2378),
.B(n_2431),
.Y(n_3113)
);

OR2x2_ASAP7_75t_L g3114 ( 
.A(n_2765),
.B(n_2293),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2922),
.A2(n_2425),
.B(n_2399),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2954),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_2653),
.Y(n_3117)
);

CKINVDCx5p33_ASAP7_75t_R g3118 ( 
.A(n_2629),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2955),
.Y(n_3119)
);

OAI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_2597),
.A2(n_2431),
.B(n_2408),
.Y(n_3120)
);

NAND2xp33_ASAP7_75t_R g3121 ( 
.A(n_2616),
.B(n_2153),
.Y(n_3121)
);

OAI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2614),
.A2(n_2408),
.B(n_2415),
.Y(n_3122)
);

AND2x6_ASAP7_75t_L g3123 ( 
.A(n_2616),
.B(n_2227),
.Y(n_3123)
);

OAI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2613),
.A2(n_2408),
.B(n_2450),
.Y(n_3124)
);

OAI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2720),
.A2(n_2408),
.B(n_2450),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2587),
.Y(n_3126)
);

OR2x2_ASAP7_75t_L g3127 ( 
.A(n_2670),
.B(n_2208),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2749),
.Y(n_3128)
);

A2O1A1Ixp33_ASAP7_75t_L g3129 ( 
.A1(n_2651),
.A2(n_2219),
.B(n_2400),
.C(n_2453),
.Y(n_3129)
);

BUFx24_ASAP7_75t_SL g3130 ( 
.A(n_2808),
.Y(n_3130)
);

CKINVDCx16_ASAP7_75t_R g3131 ( 
.A(n_2808),
.Y(n_3131)
);

BUFx8_ASAP7_75t_L g3132 ( 
.A(n_2667),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2802),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_2649),
.B(n_2267),
.Y(n_3134)
);

CKINVDCx11_ASAP7_75t_R g3135 ( 
.A(n_2742),
.Y(n_3135)
);

OAI21x1_ASAP7_75t_L g3136 ( 
.A1(n_2894),
.A2(n_2430),
.B(n_2451),
.Y(n_3136)
);

BUFx10_ASAP7_75t_L g3137 ( 
.A(n_2667),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2679),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2751),
.Y(n_3139)
);

AO21x2_ASAP7_75t_L g3140 ( 
.A1(n_2630),
.A2(n_2451),
.B(n_2410),
.Y(n_3140)
);

OAI21x1_ASAP7_75t_L g3141 ( 
.A1(n_2632),
.A2(n_2451),
.B(n_2279),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2682),
.B(n_2566),
.Y(n_3142)
);

INVx1_ASAP7_75t_SL g3143 ( 
.A(n_2940),
.Y(n_3143)
);

O2A1O1Ixp33_ASAP7_75t_L g3144 ( 
.A1(n_2733),
.A2(n_2583),
.B(n_425),
.C(n_423),
.Y(n_3144)
);

OAI21x1_ASAP7_75t_L g3145 ( 
.A1(n_2634),
.A2(n_2279),
.B(n_2410),
.Y(n_3145)
);

OAI21x1_ASAP7_75t_L g3146 ( 
.A1(n_2644),
.A2(n_2279),
.B(n_2410),
.Y(n_3146)
);

O2A1O1Ixp33_ASAP7_75t_L g3147 ( 
.A1(n_2674),
.A2(n_2583),
.B(n_428),
.C(n_424),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2606),
.B(n_424),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2827),
.Y(n_3149)
);

AND2x4_ASAP7_75t_L g3150 ( 
.A(n_2691),
.B(n_426),
.Y(n_3150)
);

A2O1A1Ixp33_ASAP7_75t_L g3151 ( 
.A1(n_2747),
.A2(n_429),
.B(n_426),
.C(n_428),
.Y(n_3151)
);

CKINVDCx20_ASAP7_75t_R g3152 ( 
.A(n_2658),
.Y(n_3152)
);

INVx3_ASAP7_75t_L g3153 ( 
.A(n_2691),
.Y(n_3153)
);

OA21x2_ASAP7_75t_L g3154 ( 
.A1(n_2809),
.A2(n_429),
.B(n_430),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2758),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2611),
.B(n_433),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2862),
.B(n_434),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2827),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2803),
.B(n_434),
.Y(n_3159)
);

O2A1O1Ixp5_ASAP7_75t_SL g3160 ( 
.A1(n_2796),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_3160)
);

OR2x6_ASAP7_75t_L g3161 ( 
.A(n_2633),
.B(n_436),
.Y(n_3161)
);

OAI21x1_ASAP7_75t_L g3162 ( 
.A1(n_2807),
.A2(n_437),
.B(n_438),
.Y(n_3162)
);

HB1xp67_ASAP7_75t_L g3163 ( 
.A(n_2663),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2654),
.Y(n_3164)
);

OR2x2_ASAP7_75t_L g3165 ( 
.A(n_2847),
.B(n_439),
.Y(n_3165)
);

AO31x2_ASAP7_75t_L g3166 ( 
.A1(n_2693),
.A2(n_442),
.A3(n_440),
.B(n_441),
.Y(n_3166)
);

AO21x1_ASAP7_75t_L g3167 ( 
.A1(n_2633),
.A2(n_440),
.B(n_441),
.Y(n_3167)
);

AOI22xp33_ASAP7_75t_L g3168 ( 
.A1(n_2758),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2596),
.B(n_2598),
.Y(n_3169)
);

AOI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_2758),
.A2(n_447),
.B1(n_444),
.B2(n_446),
.Y(n_3170)
);

AO21x2_ASAP7_75t_L g3171 ( 
.A1(n_2630),
.A2(n_780),
.B(n_447),
.Y(n_3171)
);

NAND2x1p5_ASAP7_75t_L g3172 ( 
.A(n_2862),
.B(n_448),
.Y(n_3172)
);

NAND3xp33_ASAP7_75t_L g3173 ( 
.A(n_2776),
.B(n_449),
.C(n_450),
.Y(n_3173)
);

OAI21x1_ASAP7_75t_L g3174 ( 
.A1(n_2819),
.A2(n_449),
.B(n_451),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2874),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_2766),
.Y(n_3176)
);

OAI21x1_ASAP7_75t_L g3177 ( 
.A1(n_2837),
.A2(n_452),
.B(n_453),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_2766),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2654),
.Y(n_3179)
);

A2O1A1Ixp33_ASAP7_75t_L g3180 ( 
.A1(n_2747),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2722),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2874),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2722),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2874),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2884),
.Y(n_3185)
);

OAI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2730),
.A2(n_455),
.B(n_456),
.Y(n_3186)
);

AO21x2_ASAP7_75t_L g3187 ( 
.A1(n_2672),
.A2(n_2952),
.B(n_2946),
.Y(n_3187)
);

BUFx2_ASAP7_75t_L g3188 ( 
.A(n_2888),
.Y(n_3188)
);

O2A1O1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_2699),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_SL g3190 ( 
.A1(n_2858),
.A2(n_460),
.B1(n_457),
.B2(n_459),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2619),
.B(n_459),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2744),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2884),
.Y(n_3193)
);

OAI21x1_ASAP7_75t_L g3194 ( 
.A1(n_2841),
.A2(n_460),
.B(n_461),
.Y(n_3194)
);

CKINVDCx5p33_ASAP7_75t_R g3195 ( 
.A(n_2742),
.Y(n_3195)
);

OAI21x1_ASAP7_75t_L g3196 ( 
.A1(n_2734),
.A2(n_462),
.B(n_463),
.Y(n_3196)
);

INVx3_ASAP7_75t_L g3197 ( 
.A(n_2695),
.Y(n_3197)
);

INVx3_ASAP7_75t_L g3198 ( 
.A(n_2832),
.Y(n_3198)
);

CKINVDCx20_ASAP7_75t_R g3199 ( 
.A(n_2883),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2858),
.A2(n_466),
.B1(n_462),
.B2(n_465),
.Y(n_3200)
);

AOI21x1_ASAP7_75t_L g3201 ( 
.A1(n_2930),
.A2(n_465),
.B(n_471),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2951),
.B(n_471),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2884),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2825),
.Y(n_3204)
);

OAI21x1_ASAP7_75t_L g3205 ( 
.A1(n_2843),
.A2(n_472),
.B(n_473),
.Y(n_3205)
);

BUFx8_ASAP7_75t_L g3206 ( 
.A(n_2833),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2773),
.B(n_472),
.Y(n_3207)
);

OA21x2_ASAP7_75t_L g3208 ( 
.A1(n_2851),
.A2(n_476),
.B(n_477),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2830),
.Y(n_3209)
);

AND2x4_ASAP7_75t_L g3210 ( 
.A(n_2832),
.B(n_477),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2834),
.Y(n_3211)
);

AND2x4_ASAP7_75t_L g3212 ( 
.A(n_2881),
.B(n_478),
.Y(n_3212)
);

OAI21x1_ASAP7_75t_L g3213 ( 
.A1(n_2759),
.A2(n_2760),
.B(n_2657),
.Y(n_3213)
);

AOI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_2652),
.A2(n_2773),
.B(n_2690),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2836),
.Y(n_3215)
);

OAI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_2946),
.A2(n_478),
.B(n_479),
.Y(n_3216)
);

OR2x2_ASAP7_75t_L g3217 ( 
.A(n_2885),
.B(n_480),
.Y(n_3217)
);

NAND2x1p5_ASAP7_75t_L g3218 ( 
.A(n_2901),
.B(n_480),
.Y(n_3218)
);

OAI21x1_ASAP7_75t_L g3219 ( 
.A1(n_2645),
.A2(n_481),
.B(n_483),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2850),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_2775),
.A2(n_485),
.B1(n_481),
.B2(n_484),
.Y(n_3221)
);

NAND2x1p5_ASAP7_75t_L g3222 ( 
.A(n_2902),
.B(n_484),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2744),
.Y(n_3223)
);

CKINVDCx20_ASAP7_75t_R g3224 ( 
.A(n_2883),
.Y(n_3224)
);

BUFx2_ASAP7_75t_SL g3225 ( 
.A(n_2833),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2854),
.Y(n_3226)
);

NAND2x1p5_ASAP7_75t_L g3227 ( 
.A(n_2683),
.B(n_485),
.Y(n_3227)
);

OAI21x1_ASAP7_75t_L g3228 ( 
.A1(n_2661),
.A2(n_486),
.B(n_487),
.Y(n_3228)
);

O2A1O1Ixp33_ASAP7_75t_SL g3229 ( 
.A1(n_2702),
.A2(n_488),
.B(n_486),
.C(n_487),
.Y(n_3229)
);

OAI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2952),
.A2(n_488),
.B(n_489),
.Y(n_3230)
);

BUFx4f_ASAP7_75t_L g3231 ( 
.A(n_2743),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_2958),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_3232)
);

INVx3_ASAP7_75t_L g3233 ( 
.A(n_2881),
.Y(n_3233)
);

OAI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2690),
.A2(n_490),
.B(n_492),
.Y(n_3234)
);

AO21x2_ASAP7_75t_L g3235 ( 
.A1(n_2672),
.A2(n_778),
.B(n_493),
.Y(n_3235)
);

CKINVDCx5p33_ASAP7_75t_R g3236 ( 
.A(n_2732),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_2652),
.A2(n_494),
.B(n_495),
.Y(n_3237)
);

OAI21x1_ASAP7_75t_L g3238 ( 
.A1(n_2666),
.A2(n_494),
.B(n_495),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2856),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2865),
.Y(n_3240)
);

OAI21x1_ASAP7_75t_L g3241 ( 
.A1(n_2671),
.A2(n_497),
.B(n_498),
.Y(n_3241)
);

OA21x2_ASAP7_75t_L g3242 ( 
.A1(n_2684),
.A2(n_497),
.B(n_499),
.Y(n_3242)
);

AOI221x1_ASAP7_75t_L g3243 ( 
.A1(n_2958),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.C(n_503),
.Y(n_3243)
);

CKINVDCx5p33_ASAP7_75t_R g3244 ( 
.A(n_2844),
.Y(n_3244)
);

INVx3_ASAP7_75t_L g3245 ( 
.A(n_2945),
.Y(n_3245)
);

AND2x4_ASAP7_75t_L g3246 ( 
.A(n_2945),
.B(n_501),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2687),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2866),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2889),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_2911),
.B(n_503),
.Y(n_3250)
);

OAI21x1_ASAP7_75t_L g3251 ( 
.A1(n_2697),
.A2(n_504),
.B(n_505),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2891),
.Y(n_3252)
);

OAI21x1_ASAP7_75t_L g3253 ( 
.A1(n_2706),
.A2(n_504),
.B(n_505),
.Y(n_3253)
);

NOR2xp33_ASAP7_75t_L g3254 ( 
.A(n_2904),
.B(n_506),
.Y(n_3254)
);

OA21x2_ASAP7_75t_L g3255 ( 
.A1(n_2781),
.A2(n_506),
.B(n_507),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_2916),
.A2(n_507),
.B(n_508),
.Y(n_3256)
);

OAI21x1_ASAP7_75t_L g3257 ( 
.A1(n_2721),
.A2(n_508),
.B(n_509),
.Y(n_3257)
);

INVx1_ASAP7_75t_SL g3258 ( 
.A(n_2948),
.Y(n_3258)
);

AOI221x1_ASAP7_75t_L g3259 ( 
.A1(n_2826),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.C(n_513),
.Y(n_3259)
);

OAI21x1_ASAP7_75t_L g3260 ( 
.A1(n_2725),
.A2(n_510),
.B(n_511),
.Y(n_3260)
);

OAI21x1_ASAP7_75t_L g3261 ( 
.A1(n_2728),
.A2(n_512),
.B(n_513),
.Y(n_3261)
);

BUFx3_ASAP7_75t_L g3262 ( 
.A(n_2948),
.Y(n_3262)
);

CKINVDCx20_ASAP7_75t_R g3263 ( 
.A(n_2953),
.Y(n_3263)
);

INVxp67_ASAP7_75t_L g3264 ( 
.A(n_2919),
.Y(n_3264)
);

NAND2x1p5_ASAP7_75t_L g3265 ( 
.A(n_2919),
.B(n_514),
.Y(n_3265)
);

AOI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_2659),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_2743),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_2863),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3045),
.Y(n_3269)
);

BUFx3_ASAP7_75t_L g3270 ( 
.A(n_3135),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2984),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_2987),
.B(n_2961),
.Y(n_3272)
);

BUFx2_ASAP7_75t_L g3273 ( 
.A(n_3132),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3028),
.A2(n_2800),
.B1(n_2586),
.B2(n_2769),
.Y(n_3274)
);

AOI221xp5_ASAP7_75t_L g3275 ( 
.A1(n_3018),
.A2(n_2933),
.B1(n_2908),
.B2(n_2873),
.C(n_2696),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2975),
.B(n_2622),
.Y(n_3276)
);

BUFx2_ASAP7_75t_L g3277 ( 
.A(n_3132),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3082),
.B(n_2698),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2978),
.Y(n_3279)
);

AOI22xp33_ASAP7_75t_SL g3280 ( 
.A1(n_3060),
.A2(n_2757),
.B1(n_2624),
.B2(n_2933),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_3028),
.A2(n_2835),
.B1(n_2890),
.B2(n_2828),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_2979),
.B(n_2838),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2990),
.Y(n_3283)
);

AOI21xp33_ASAP7_75t_L g3284 ( 
.A1(n_3031),
.A2(n_3093),
.B(n_3096),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3250),
.B(n_2848),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_3159),
.B(n_2915),
.Y(n_3286)
);

OAI211xp5_ASAP7_75t_SL g3287 ( 
.A1(n_3127),
.A2(n_2660),
.B(n_2906),
.C(n_2678),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3128),
.B(n_2934),
.Y(n_3288)
);

AOI222xp33_ASAP7_75t_L g3289 ( 
.A1(n_2986),
.A2(n_3232),
.B1(n_3200),
.B2(n_3231),
.C1(n_3072),
.C2(n_3019),
.Y(n_3289)
);

NAND2x1p5_ASAP7_75t_L g3290 ( 
.A(n_3231),
.B(n_2692),
.Y(n_3290)
);

INVx2_ASAP7_75t_SL g3291 ( 
.A(n_2982),
.Y(n_3291)
);

OAI22xp33_ASAP7_75t_SL g3292 ( 
.A1(n_3131),
.A2(n_2621),
.B1(n_2609),
.B2(n_2941),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3139),
.B(n_2934),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3094),
.Y(n_3294)
);

HB1xp67_ASAP7_75t_L g3295 ( 
.A(n_3094),
.Y(n_3295)
);

OAI22xp5_ASAP7_75t_SL g3296 ( 
.A1(n_3152),
.A2(n_2646),
.B1(n_2637),
.B2(n_2704),
.Y(n_3296)
);

AND2x4_ASAP7_75t_L g3297 ( 
.A(n_2968),
.B(n_2692),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_SL g3298 ( 
.A1(n_3060),
.A2(n_3225),
.B1(n_3022),
.B2(n_3081),
.Y(n_3298)
);

OAI21xp5_ASAP7_75t_SL g3299 ( 
.A1(n_3033),
.A2(n_2726),
.B(n_2713),
.Y(n_3299)
);

AOI221xp5_ASAP7_75t_L g3300 ( 
.A1(n_3200),
.A2(n_3232),
.B1(n_2986),
.B2(n_2977),
.C(n_3072),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_3033),
.A2(n_2892),
.B1(n_2791),
.B2(n_2669),
.Y(n_3301)
);

INVx4_ASAP7_75t_SL g3302 ( 
.A(n_2965),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2998),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_3020),
.A2(n_2887),
.B1(n_2886),
.B2(n_2726),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3002),
.Y(n_3305)
);

CKINVDCx20_ASAP7_75t_R g3306 ( 
.A(n_2962),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3050),
.B(n_2686),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_3001),
.Y(n_3308)
);

NOR2x1_ASAP7_75t_R g3309 ( 
.A(n_2995),
.B(n_2880),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_R g3310 ( 
.A(n_3030),
.B(n_2694),
.Y(n_3310)
);

CKINVDCx20_ASAP7_75t_R g3311 ( 
.A(n_3030),
.Y(n_3311)
);

BUFx6f_ASAP7_75t_L g3312 ( 
.A(n_2965),
.Y(n_3312)
);

CKINVDCx8_ASAP7_75t_R g3313 ( 
.A(n_3037),
.Y(n_3313)
);

OAI22xp33_ASAP7_75t_L g3314 ( 
.A1(n_3161),
.A2(n_2935),
.B1(n_2939),
.B2(n_2918),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_SL g3315 ( 
.A1(n_3267),
.A2(n_2713),
.B1(n_2793),
.B2(n_2771),
.Y(n_3315)
);

CKINVDCx16_ASAP7_75t_R g3316 ( 
.A(n_3199),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_3034),
.A2(n_2793),
.B1(n_2814),
.B2(n_2799),
.Y(n_3317)
);

CKINVDCx20_ASAP7_75t_R g3318 ( 
.A(n_3224),
.Y(n_3318)
);

AND2x4_ASAP7_75t_L g3319 ( 
.A(n_3111),
.B(n_2981),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3051),
.B(n_2604),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_2997),
.A2(n_3214),
.B(n_3063),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_3005),
.A2(n_2799),
.B1(n_2814),
.B2(n_2878),
.Y(n_3322)
);

OR2x6_ASAP7_75t_L g3323 ( 
.A(n_3161),
.B(n_2824),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3053),
.B(n_2605),
.Y(n_3324)
);

CKINVDCx20_ASAP7_75t_R g3325 ( 
.A(n_3118),
.Y(n_3325)
);

CKINVDCx8_ASAP7_75t_R g3326 ( 
.A(n_3195),
.Y(n_3326)
);

INVx1_ASAP7_75t_SL g3327 ( 
.A(n_3236),
.Y(n_3327)
);

INVx4_ASAP7_75t_L g3328 ( 
.A(n_2993),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3005),
.A2(n_2746),
.B1(n_2939),
.B2(n_2935),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_3015),
.A2(n_2920),
.B1(n_2924),
.B2(n_2917),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3109),
.B(n_2918),
.Y(n_3331)
);

NOR2x1_ASAP7_75t_SL g3332 ( 
.A(n_3161),
.B(n_2663),
.Y(n_3332)
);

INVx2_ASAP7_75t_SL g3333 ( 
.A(n_3038),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3016),
.B(n_2648),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_2992),
.B(n_2987),
.Y(n_3335)
);

AOI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_3100),
.A2(n_2949),
.B1(n_2944),
.B2(n_2777),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_3052),
.A2(n_2685),
.B1(n_2947),
.B2(n_2615),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_2992),
.B(n_2711),
.Y(n_3338)
);

INVx2_ASAP7_75t_SL g3339 ( 
.A(n_3038),
.Y(n_3339)
);

BUFx2_ASAP7_75t_L g3340 ( 
.A(n_3044),
.Y(n_3340)
);

AOI221xp5_ASAP7_75t_L g3341 ( 
.A1(n_2977),
.A2(n_2685),
.B1(n_2753),
.B2(n_2778),
.C(n_2708),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3048),
.B(n_2648),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3138),
.B(n_523),
.Y(n_3343)
);

AOI22xp33_ASAP7_75t_L g3344 ( 
.A1(n_3052),
.A2(n_2947),
.B1(n_2937),
.B2(n_2929),
.Y(n_3344)
);

NOR3xp33_ASAP7_75t_SL g3345 ( 
.A(n_3121),
.B(n_2895),
.C(n_2817),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3106),
.B(n_524),
.Y(n_3346)
);

NOR2x1_ASAP7_75t_SL g3347 ( 
.A(n_3107),
.B(n_3140),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3009),
.Y(n_3348)
);

INVx1_ASAP7_75t_SL g3349 ( 
.A(n_3244),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_3017),
.A2(n_2701),
.B1(n_2846),
.B2(n_2829),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2963),
.B(n_2648),
.Y(n_3351)
);

OAI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_3265),
.A2(n_2764),
.B1(n_2729),
.B2(n_2738),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3097),
.A2(n_2860),
.B1(n_2855),
.B2(n_2714),
.Y(n_3353)
);

CKINVDCx5p33_ASAP7_75t_R g3354 ( 
.A(n_2996),
.Y(n_3354)
);

AOI222xp33_ASAP7_75t_L g3355 ( 
.A1(n_3206),
.A2(n_2717),
.B1(n_2710),
.B2(n_2718),
.C1(n_2715),
.C2(n_2703),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3006),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3007),
.Y(n_3357)
);

AOI21xp5_ASAP7_75t_SL g3358 ( 
.A1(n_3151),
.A2(n_2812),
.B(n_2787),
.Y(n_3358)
);

NAND3xp33_ASAP7_75t_SL g3359 ( 
.A(n_3190),
.B(n_2792),
.C(n_2768),
.Y(n_3359)
);

INVx1_ASAP7_75t_SL g3360 ( 
.A(n_3114),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3074),
.Y(n_3361)
);

BUFx2_ASAP7_75t_L g3362 ( 
.A(n_3206),
.Y(n_3362)
);

AOI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_3064),
.A2(n_2724),
.B1(n_2723),
.B2(n_2785),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_2989),
.B(n_525),
.Y(n_3364)
);

INVx5_ASAP7_75t_L g3365 ( 
.A(n_3123),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_3111),
.B(n_2668),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3064),
.A2(n_2806),
.B1(n_2798),
.B2(n_2620),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_3035),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_2989),
.B(n_526),
.Y(n_3369)
);

INVxp67_ASAP7_75t_SL g3370 ( 
.A(n_3104),
.Y(n_3370)
);

INVxp67_ASAP7_75t_L g3371 ( 
.A(n_2994),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_3042),
.B(n_2897),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3066),
.B(n_527),
.Y(n_3373)
);

OAI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3265),
.A2(n_2739),
.B1(n_2741),
.B2(n_2727),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3075),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3080),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2973),
.B(n_2805),
.Y(n_3377)
);

AND2x4_ASAP7_75t_L g3378 ( 
.A(n_2981),
.B(n_2668),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_SL g3379 ( 
.A1(n_2966),
.A2(n_2880),
.B1(n_2928),
.B2(n_2879),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3083),
.B(n_527),
.Y(n_3380)
);

CKINVDCx5p33_ASAP7_75t_R g3381 ( 
.A(n_3263),
.Y(n_3381)
);

BUFx12f_ASAP7_75t_L g3382 ( 
.A(n_3137),
.Y(n_3382)
);

OAI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3023),
.A2(n_2815),
.B1(n_2822),
.B2(n_2752),
.Y(n_3383)
);

OAI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3264),
.A2(n_2641),
.B1(n_2642),
.B2(n_2640),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3024),
.A2(n_3092),
.B1(n_3014),
.B2(n_3190),
.Y(n_3385)
);

OR2x2_ASAP7_75t_L g3386 ( 
.A(n_3143),
.B(n_2711),
.Y(n_3386)
);

BUFx10_ASAP7_75t_L g3387 ( 
.A(n_3150),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_3024),
.A2(n_2770),
.B1(n_2789),
.B2(n_2761),
.Y(n_3388)
);

OAI211xp5_ASAP7_75t_L g3389 ( 
.A1(n_3014),
.A2(n_2869),
.B(n_2853),
.C(n_2804),
.Y(n_3389)
);

OAI211xp5_ASAP7_75t_L g3390 ( 
.A1(n_3087),
.A2(n_2795),
.B(n_2676),
.C(n_2662),
.Y(n_3390)
);

CKINVDCx11_ASAP7_75t_R g3391 ( 
.A(n_3137),
.Y(n_3391)
);

INVx4_ASAP7_75t_SL g3392 ( 
.A(n_3123),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_3103),
.B(n_528),
.Y(n_3393)
);

OAI221xp5_ASAP7_75t_L g3394 ( 
.A1(n_3101),
.A2(n_2905),
.B1(n_2647),
.B2(n_2631),
.C(n_2882),
.Y(n_3394)
);

BUFx12f_ASAP7_75t_L g3395 ( 
.A(n_3227),
.Y(n_3395)
);

INVx3_ASAP7_75t_L g3396 ( 
.A(n_3079),
.Y(n_3396)
);

OR2x2_ASAP7_75t_L g3397 ( 
.A(n_3143),
.B(n_2711),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3103),
.B(n_529),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3043),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3099),
.B(n_2805),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_SL g3401 ( 
.A1(n_3197),
.A2(n_2880),
.B1(n_2928),
.B2(n_2879),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3086),
.Y(n_3402)
);

INVx4_ASAP7_75t_SL g3403 ( 
.A(n_3123),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_2976),
.B(n_2805),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3110),
.Y(n_3405)
);

INVx1_ASAP7_75t_SL g3406 ( 
.A(n_3188),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3116),
.Y(n_3407)
);

OAI22xp33_ASAP7_75t_L g3408 ( 
.A1(n_3264),
.A2(n_2956),
.B1(n_2957),
.B2(n_2677),
.Y(n_3408)
);

HB1xp67_ASAP7_75t_L g3409 ( 
.A(n_3104),
.Y(n_3409)
);

AND2x4_ASAP7_75t_L g3410 ( 
.A(n_3079),
.B(n_2677),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3126),
.B(n_2754),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3025),
.A2(n_2772),
.B(n_2750),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3021),
.A2(n_2956),
.B1(n_2750),
.B2(n_2818),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3046),
.B(n_2754),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3055),
.B(n_529),
.Y(n_3415)
);

AO22x2_ASAP7_75t_L g3416 ( 
.A1(n_3149),
.A2(n_2960),
.B1(n_2910),
.B2(n_2754),
.Y(n_3416)
);

CKINVDCx20_ASAP7_75t_R g3417 ( 
.A(n_3013),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3059),
.Y(n_3418)
);

BUFx2_ASAP7_75t_SL g3419 ( 
.A(n_3123),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_L g3420 ( 
.A(n_3067),
.B(n_530),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3125),
.A2(n_2818),
.B(n_2772),
.Y(n_3421)
);

BUFx2_ASAP7_75t_L g3422 ( 
.A(n_3011),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3133),
.B(n_531),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3119),
.Y(n_3424)
);

OR2x2_ASAP7_75t_L g3425 ( 
.A(n_2972),
.B(n_2910),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3085),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3165),
.B(n_531),
.Y(n_3427)
);

AOI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_3254),
.A2(n_2870),
.B1(n_2880),
.B2(n_2818),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3150),
.B(n_532),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3010),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_3125),
.A2(n_2880),
.B(n_2603),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3130),
.A2(n_2786),
.B1(n_2801),
.B2(n_2603),
.Y(n_3432)
);

AOI22xp33_ASAP7_75t_SL g3433 ( 
.A1(n_3197),
.A2(n_2960),
.B1(n_2910),
.B2(n_2786),
.Y(n_3433)
);

AND2x4_ASAP7_75t_L g3434 ( 
.A(n_2988),
.B(n_2960),
.Y(n_3434)
);

AOI22xp33_ASAP7_75t_L g3435 ( 
.A1(n_3032),
.A2(n_2786),
.B1(n_2801),
.B2(n_2603),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3010),
.Y(n_3436)
);

OAI21x1_ASAP7_75t_L g3437 ( 
.A1(n_2983),
.A2(n_2999),
.B(n_3091),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3093),
.A2(n_532),
.B(n_533),
.Y(n_3438)
);

OAI22xp5_ASAP7_75t_L g3439 ( 
.A1(n_3155),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_3439)
);

CKINVDCx5p33_ASAP7_75t_R g3440 ( 
.A(n_3070),
.Y(n_3440)
);

INVx1_ASAP7_75t_SL g3441 ( 
.A(n_3134),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3217),
.B(n_534),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3004),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_L g3444 ( 
.A1(n_3004),
.A2(n_540),
.B1(n_537),
.B2(n_539),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_3124),
.A2(n_541),
.B(n_542),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3089),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3098),
.B(n_541),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3089),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3101),
.A2(n_546),
.B1(n_544),
.B2(n_545),
.Y(n_3449)
);

AOI22xp33_ASAP7_75t_L g3450 ( 
.A1(n_2970),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_3450)
);

AO21x2_ASAP7_75t_L g3451 ( 
.A1(n_3237),
.A2(n_547),
.B(n_548),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_3168),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3169),
.B(n_550),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_3068),
.B(n_552),
.Y(n_3454)
);

OR2x6_ASAP7_75t_L g3455 ( 
.A(n_3218),
.B(n_553),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3164),
.Y(n_3456)
);

INVx3_ASAP7_75t_L g3457 ( 
.A(n_3054),
.Y(n_3457)
);

AOI22xp5_ASAP7_75t_L g3458 ( 
.A1(n_3108),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_R g3459 ( 
.A(n_3153),
.B(n_554),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3170),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_3460)
);

INVx3_ASAP7_75t_L g3461 ( 
.A(n_2985),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3202),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3169),
.B(n_560),
.Y(n_3463)
);

AO21x2_ASAP7_75t_L g3464 ( 
.A1(n_3237),
.A2(n_561),
.B(n_564),
.Y(n_3464)
);

AND2x6_ASAP7_75t_L g3465 ( 
.A(n_2971),
.B(n_564),
.Y(n_3465)
);

BUFx2_ASAP7_75t_L g3466 ( 
.A(n_3117),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_3077),
.Y(n_3467)
);

AOI22xp5_ASAP7_75t_L g3468 ( 
.A1(n_3070),
.A2(n_568),
.B1(n_565),
.B2(n_566),
.Y(n_3468)
);

BUFx6f_ASAP7_75t_L g3469 ( 
.A(n_2985),
.Y(n_3469)
);

O2A1O1Ixp33_ASAP7_75t_SL g3470 ( 
.A1(n_3095),
.A2(n_570),
.B(n_568),
.C(n_569),
.Y(n_3470)
);

AOI222xp33_ASAP7_75t_L g3471 ( 
.A1(n_3234),
.A2(n_569),
.B1(n_572),
.B2(n_573),
.C1(n_574),
.C2(n_575),
.Y(n_3471)
);

CKINVDCx20_ASAP7_75t_R g3472 ( 
.A(n_3047),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3210),
.B(n_3212),
.Y(n_3473)
);

OAI22xp33_ASAP7_75t_L g3474 ( 
.A1(n_3218),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3202),
.Y(n_3475)
);

INVx1_ASAP7_75t_SL g3476 ( 
.A(n_3056),
.Y(n_3476)
);

HB1xp67_ASAP7_75t_L g3477 ( 
.A(n_2991),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3204),
.B(n_578),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_L g3479 ( 
.A1(n_2970),
.A2(n_582),
.B1(n_578),
.B2(n_581),
.Y(n_3479)
);

AOI22xp33_ASAP7_75t_L g3480 ( 
.A1(n_2967),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3209),
.B(n_583),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_3056),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3211),
.B(n_3215),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3210),
.Y(n_3484)
);

NOR2x1_ASAP7_75t_SL g3485 ( 
.A(n_3107),
.B(n_584),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3212),
.Y(n_3486)
);

BUFx4f_ASAP7_75t_L g3487 ( 
.A(n_3222),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3179),
.Y(n_3488)
);

AOI21xp33_ASAP7_75t_L g3489 ( 
.A1(n_3031),
.A2(n_584),
.B(n_585),
.Y(n_3489)
);

AO31x2_ASAP7_75t_L g3490 ( 
.A1(n_3181),
.A2(n_587),
.A3(n_585),
.B(n_586),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3183),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_3142),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3192),
.Y(n_3493)
);

OAI22xp33_ASAP7_75t_L g3494 ( 
.A1(n_3222),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.Y(n_3494)
);

O2A1O1Ixp33_ASAP7_75t_L g3495 ( 
.A1(n_3026),
.A2(n_595),
.B(n_593),
.C(n_594),
.Y(n_3495)
);

BUFx3_ASAP7_75t_L g3496 ( 
.A(n_3090),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3246),
.Y(n_3497)
);

CKINVDCx16_ASAP7_75t_R g3498 ( 
.A(n_2971),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3220),
.B(n_3226),
.Y(n_3499)
);

INVx3_ASAP7_75t_L g3500 ( 
.A(n_2988),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_SL g3501 ( 
.A1(n_3172),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3239),
.B(n_3240),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3246),
.B(n_598),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3057),
.B(n_599),
.Y(n_3504)
);

OR2x2_ASAP7_75t_L g3505 ( 
.A(n_3012),
.B(n_3258),
.Y(n_3505)
);

OAI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3073),
.A2(n_3227),
.B1(n_3266),
.B2(n_3268),
.Y(n_3506)
);

OR2x2_ASAP7_75t_L g3507 ( 
.A(n_3012),
.B(n_599),
.Y(n_3507)
);

INVx2_ASAP7_75t_SL g3508 ( 
.A(n_3057),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3166),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3248),
.B(n_600),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_SL g3511 ( 
.A1(n_3029),
.A2(n_3076),
.B1(n_3112),
.B2(n_3234),
.Y(n_3511)
);

AO21x2_ASAP7_75t_L g3512 ( 
.A1(n_3173),
.A2(n_601),
.B(n_602),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3223),
.Y(n_3513)
);

AND2x4_ASAP7_75t_L g3514 ( 
.A(n_2980),
.B(n_603),
.Y(n_3514)
);

OAI22xp5_ASAP7_75t_L g3515 ( 
.A1(n_3216),
.A2(n_603),
.B1(n_605),
.B2(n_606),
.Y(n_3515)
);

AOI21xp33_ASAP7_75t_L g3516 ( 
.A1(n_3289),
.A2(n_3147),
.B(n_3144),
.Y(n_3516)
);

NOR2x1_ASAP7_75t_SL g3517 ( 
.A(n_3419),
.B(n_3102),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3300),
.A2(n_3102),
.B1(n_2967),
.B2(n_3167),
.Y(n_3518)
);

OAI22xp33_ASAP7_75t_L g3519 ( 
.A1(n_3328),
.A2(n_3243),
.B1(n_3216),
.B2(n_3230),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3467),
.B(n_3249),
.Y(n_3520)
);

AOI22xp33_ASAP7_75t_SL g3521 ( 
.A1(n_3332),
.A2(n_2980),
.B1(n_3176),
.B2(n_3153),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3376),
.B(n_3252),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3418),
.B(n_3008),
.Y(n_3523)
);

AOI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3301),
.A2(n_3230),
.B1(n_3058),
.B2(n_3061),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3331),
.A2(n_3274),
.B1(n_3296),
.B2(n_3314),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3441),
.B(n_3381),
.Y(n_3526)
);

AND2x2_ASAP7_75t_L g3527 ( 
.A(n_3276),
.B(n_3282),
.Y(n_3527)
);

OAI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_3280),
.A2(n_3180),
.B1(n_3189),
.B2(n_3113),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3278),
.B(n_3258),
.Y(n_3529)
);

AOI22xp33_ASAP7_75t_L g3530 ( 
.A1(n_3323),
.A2(n_3058),
.B1(n_3061),
.B2(n_3078),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_L g3531 ( 
.A1(n_3323),
.A2(n_3078),
.B1(n_3187),
.B2(n_3113),
.Y(n_3531)
);

INVx4_ASAP7_75t_L g3532 ( 
.A(n_3365),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3271),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3426),
.B(n_3008),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3335),
.B(n_3008),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3370),
.B(n_3158),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3315),
.A2(n_3187),
.B1(n_3186),
.B2(n_3171),
.Y(n_3537)
);

OAI222xp33_ASAP7_75t_L g3538 ( 
.A1(n_3298),
.A2(n_3000),
.B1(n_3062),
.B2(n_3189),
.C1(n_3157),
.C2(n_3069),
.Y(n_3538)
);

OAI22xp5_ASAP7_75t_L g3539 ( 
.A1(n_3487),
.A2(n_3173),
.B1(n_3221),
.B2(n_3207),
.Y(n_3539)
);

AOI221xp5_ASAP7_75t_L g3540 ( 
.A1(n_3287),
.A2(n_3256),
.B1(n_3148),
.B2(n_3156),
.C(n_3147),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_3275),
.A2(n_3186),
.B1(n_3235),
.B2(n_3171),
.Y(n_3541)
);

OAI22xp33_ASAP7_75t_L g3542 ( 
.A1(n_3328),
.A2(n_3259),
.B1(n_3069),
.B2(n_3178),
.Y(n_3542)
);

AOI22xp33_ASAP7_75t_L g3543 ( 
.A1(n_3506),
.A2(n_3281),
.B1(n_3385),
.B2(n_3304),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3359),
.A2(n_3235),
.B1(n_3140),
.B2(n_3256),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_SL g3545 ( 
.A1(n_3332),
.A2(n_3176),
.B1(n_3178),
.B2(n_3154),
.Y(n_3545)
);

OAI22xp33_ASAP7_75t_L g3546 ( 
.A1(n_3455),
.A2(n_3120),
.B1(n_3207),
.B2(n_3124),
.Y(n_3546)
);

OAI211xp5_ASAP7_75t_L g3547 ( 
.A1(n_3459),
.A2(n_3144),
.B(n_3156),
.C(n_3148),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3361),
.B(n_2964),
.Y(n_3548)
);

OAI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3487),
.A2(n_3129),
.B1(n_3120),
.B2(n_3191),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3279),
.Y(n_3550)
);

OAI221xp5_ASAP7_75t_L g3551 ( 
.A1(n_3330),
.A2(n_3355),
.B1(n_3299),
.B2(n_3468),
.C(n_3455),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_SL g3552 ( 
.A(n_3273),
.B(n_2991),
.Y(n_3552)
);

NAND3xp33_ASAP7_75t_L g3553 ( 
.A(n_3471),
.B(n_3182),
.C(n_3175),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_L g3554 ( 
.A1(n_3465),
.A2(n_3122),
.B1(n_2964),
.B2(n_3191),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3375),
.B(n_3184),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3283),
.B(n_3185),
.Y(n_3556)
);

OAI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3437),
.A2(n_2974),
.B(n_3062),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3303),
.Y(n_3558)
);

OA21x2_ASAP7_75t_L g3559 ( 
.A1(n_3321),
.A2(n_3203),
.B(n_3193),
.Y(n_3559)
);

HB1xp67_ASAP7_75t_L g3560 ( 
.A(n_3409),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3498),
.B(n_3262),
.Y(n_3561)
);

AOI22xp33_ASAP7_75t_L g3562 ( 
.A1(n_3465),
.A2(n_3198),
.B1(n_3245),
.B2(n_3233),
.Y(n_3562)
);

AOI22xp33_ASAP7_75t_L g3563 ( 
.A1(n_3286),
.A2(n_3198),
.B1(n_3245),
.B2(n_3233),
.Y(n_3563)
);

OR2x2_ASAP7_75t_L g3564 ( 
.A(n_3294),
.B(n_3163),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_SL g3565 ( 
.A1(n_3309),
.A2(n_3208),
.B(n_3027),
.Y(n_3565)
);

OR2x2_ASAP7_75t_SL g3566 ( 
.A(n_3316),
.B(n_3163),
.Y(n_3566)
);

BUFx6f_ASAP7_75t_L g3567 ( 
.A(n_3312),
.Y(n_3567)
);

BUFx5_ASAP7_75t_L g3568 ( 
.A(n_3297),
.Y(n_3568)
);

AND2x4_ASAP7_75t_L g3569 ( 
.A(n_3295),
.B(n_3071),
.Y(n_3569)
);

AOI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3372),
.A2(n_3071),
.B1(n_3115),
.B2(n_3247),
.Y(n_3570)
);

OR2x2_ASAP7_75t_L g3571 ( 
.A(n_3436),
.B(n_3166),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3308),
.Y(n_3572)
);

OAI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3395),
.A2(n_3255),
.B1(n_3242),
.B2(n_3201),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3305),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_SL g3575 ( 
.A1(n_3473),
.A2(n_3049),
.B1(n_3039),
.B2(n_3141),
.Y(n_3575)
);

AND2x4_ASAP7_75t_SL g3576 ( 
.A(n_3387),
.B(n_3105),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3360),
.B(n_3166),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3356),
.B(n_3049),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3317),
.A2(n_3242),
.B1(n_3229),
.B2(n_3219),
.Y(n_3579)
);

OAI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3501),
.A2(n_3228),
.B1(n_3241),
.B2(n_3238),
.Y(n_3580)
);

AOI221xp5_ASAP7_75t_L g3581 ( 
.A1(n_3284),
.A2(n_3039),
.B1(n_3160),
.B2(n_611),
.C(n_613),
.Y(n_3581)
);

OAI222xp33_ASAP7_75t_L g3582 ( 
.A1(n_3440),
.A2(n_3084),
.B1(n_3213),
.B2(n_3146),
.C1(n_3145),
.C2(n_3205),
.Y(n_3582)
);

AOI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_3341),
.A2(n_3196),
.B1(n_3253),
.B2(n_3251),
.Y(n_3583)
);

AOI222xp33_ASAP7_75t_L g3584 ( 
.A1(n_3277),
.A2(n_3261),
.B1(n_3260),
.B2(n_3257),
.C1(n_3194),
.C2(n_3177),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3413),
.A2(n_3065),
.B(n_3041),
.Y(n_3585)
);

AOI221xp5_ASAP7_75t_L g3586 ( 
.A1(n_3384),
.A2(n_607),
.B1(n_608),
.B2(n_613),
.C(n_617),
.Y(n_3586)
);

OR2x2_ASAP7_75t_L g3587 ( 
.A(n_3446),
.B(n_608),
.Y(n_3587)
);

OAI221xp5_ASAP7_75t_L g3588 ( 
.A1(n_3345),
.A2(n_3174),
.B1(n_3162),
.B2(n_3088),
.C(n_621),
.Y(n_3588)
);

A2O1A1Ixp33_ASAP7_75t_SL g3589 ( 
.A1(n_3420),
.A2(n_3036),
.B(n_3040),
.C(n_3136),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3357),
.B(n_2969),
.Y(n_3590)
);

INVx1_ASAP7_75t_SL g3591 ( 
.A(n_3340),
.Y(n_3591)
);

AOI22xp33_ASAP7_75t_L g3592 ( 
.A1(n_3285),
.A2(n_3346),
.B1(n_3383),
.B2(n_3515),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3466),
.B(n_617),
.Y(n_3593)
);

A2O1A1Ixp33_ASAP7_75t_L g3594 ( 
.A1(n_3495),
.A2(n_3003),
.B(n_620),
.C(n_622),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_3392),
.B(n_619),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3348),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3368),
.Y(n_3597)
);

AOI222xp33_ASAP7_75t_L g3598 ( 
.A1(n_3362),
.A2(n_620),
.B1(n_622),
.B2(n_624),
.C1(n_625),
.C2(n_626),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3288),
.B(n_627),
.Y(n_3599)
);

AOI211xp5_ASAP7_75t_L g3600 ( 
.A1(n_3292),
.A2(n_628),
.B(n_629),
.C(n_630),
.Y(n_3600)
);

OAI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3365),
.A2(n_628),
.B1(n_629),
.B2(n_632),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3272),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_L g3603 ( 
.A1(n_3329),
.A2(n_632),
.B1(n_633),
.B2(n_634),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_3371),
.B(n_634),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3352),
.A2(n_635),
.B(n_636),
.Y(n_3605)
);

AOI22xp5_ASAP7_75t_L g3606 ( 
.A1(n_3336),
.A2(n_635),
.B1(n_637),
.B2(n_638),
.Y(n_3606)
);

AO21x2_ASAP7_75t_L g3607 ( 
.A1(n_3489),
.A2(n_637),
.B(n_638),
.Y(n_3607)
);

OAI211xp5_ASAP7_75t_L g3608 ( 
.A1(n_3310),
.A2(n_639),
.B(n_640),
.C(n_641),
.Y(n_3608)
);

OAI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3290),
.A2(n_639),
.B1(n_640),
.B2(n_641),
.Y(n_3609)
);

NAND3xp33_ASAP7_75t_L g3610 ( 
.A(n_3433),
.B(n_642),
.C(n_643),
.Y(n_3610)
);

AOI221xp5_ASAP7_75t_L g3611 ( 
.A1(n_3453),
.A2(n_642),
.B1(n_644),
.B2(n_645),
.C(n_646),
.Y(n_3611)
);

OAI211xp5_ASAP7_75t_L g3612 ( 
.A1(n_3511),
.A2(n_645),
.B(n_646),
.C(n_647),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3399),
.Y(n_3613)
);

OR2x2_ASAP7_75t_L g3614 ( 
.A(n_3448),
.B(n_647),
.Y(n_3614)
);

INVx5_ASAP7_75t_SL g3615 ( 
.A(n_3312),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3293),
.A2(n_648),
.B1(n_649),
.B2(n_650),
.Y(n_3616)
);

OR2x6_ASAP7_75t_L g3617 ( 
.A(n_3431),
.B(n_651),
.Y(n_3617)
);

OAI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3514),
.A2(n_651),
.B1(n_652),
.B2(n_653),
.Y(n_3618)
);

HB1xp67_ASAP7_75t_L g3619 ( 
.A(n_3422),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3430),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3474),
.A2(n_652),
.B1(n_653),
.B2(n_654),
.Y(n_3621)
);

CKINVDCx14_ASAP7_75t_R g3622 ( 
.A(n_3311),
.Y(n_3622)
);

OAI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_3514),
.A2(n_654),
.B1(n_655),
.B2(n_656),
.Y(n_3623)
);

AOI22xp33_ASAP7_75t_SL g3624 ( 
.A1(n_3387),
.A2(n_655),
.B1(n_656),
.B2(n_657),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3483),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3494),
.A2(n_658),
.B1(n_659),
.B2(n_660),
.Y(n_3626)
);

BUFx12f_ASAP7_75t_L g3627 ( 
.A(n_3391),
.Y(n_3627)
);

OAI22xp5_ASAP7_75t_L g3628 ( 
.A1(n_3365),
.A2(n_658),
.B1(n_659),
.B2(n_662),
.Y(n_3628)
);

NAND4xp25_ASAP7_75t_L g3629 ( 
.A(n_3435),
.B(n_663),
.C(n_664),
.D(n_665),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3269),
.B(n_777),
.Y(n_3630)
);

AOI22xp33_ASAP7_75t_L g3631 ( 
.A1(n_3484),
.A2(n_663),
.B1(n_665),
.B2(n_666),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3393),
.B(n_777),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_L g3633 ( 
.A1(n_3486),
.A2(n_666),
.B1(n_667),
.B2(n_668),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3497),
.A2(n_667),
.B1(n_668),
.B2(n_670),
.Y(n_3634)
);

OR2x2_ASAP7_75t_L g3635 ( 
.A(n_3406),
.B(n_670),
.Y(n_3635)
);

OAI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3322),
.A2(n_671),
.B1(n_672),
.B2(n_673),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3439),
.A2(n_671),
.B1(n_674),
.B2(n_675),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3398),
.B(n_776),
.Y(n_3638)
);

OAI211xp5_ASAP7_75t_L g3639 ( 
.A1(n_3313),
.A2(n_674),
.B(n_675),
.C(n_676),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3402),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3499),
.Y(n_3641)
);

OAI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3458),
.A2(n_677),
.B1(n_678),
.B2(n_679),
.Y(n_3642)
);

OR3x1_ASAP7_75t_L g3643 ( 
.A(n_3302),
.B(n_775),
.C(n_681),
.Y(n_3643)
);

AND2x2_ASAP7_75t_L g3644 ( 
.A(n_3319),
.B(n_3405),
.Y(n_3644)
);

OAI211xp5_ASAP7_75t_L g3645 ( 
.A1(n_3429),
.A2(n_678),
.B(n_681),
.C(n_682),
.Y(n_3645)
);

BUFx4f_ASAP7_75t_L g3646 ( 
.A(n_3291),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3319),
.B(n_3407),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3452),
.A2(n_3460),
.B1(n_3374),
.B2(n_3504),
.Y(n_3648)
);

AOI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3504),
.A2(n_682),
.B1(n_683),
.B2(n_684),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3502),
.Y(n_3650)
);

OAI33xp33_ASAP7_75t_L g3651 ( 
.A1(n_3463),
.A2(n_684),
.A3(n_685),
.B1(n_686),
.B2(n_687),
.B3(n_688),
.Y(n_3651)
);

AOI22xp33_ASAP7_75t_SL g3652 ( 
.A1(n_3485),
.A2(n_685),
.B1(n_686),
.B2(n_687),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3424),
.Y(n_3653)
);

OAI22xp33_ASAP7_75t_SL g3654 ( 
.A1(n_3396),
.A2(n_3297),
.B1(n_3476),
.B2(n_3386),
.Y(n_3654)
);

OAI211xp5_ASAP7_75t_L g3655 ( 
.A1(n_3450),
.A2(n_689),
.B(n_690),
.C(n_691),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3462),
.B(n_3475),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3364),
.B(n_775),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_SL g3658 ( 
.A1(n_3347),
.A2(n_689),
.B1(n_690),
.B2(n_693),
.Y(n_3658)
);

AOI22xp33_ASAP7_75t_L g3659 ( 
.A1(n_3388),
.A2(n_694),
.B1(n_695),
.B2(n_696),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3449),
.A2(n_695),
.B1(n_697),
.B2(n_700),
.Y(n_3660)
);

INVx1_ASAP7_75t_SL g3661 ( 
.A(n_3327),
.Y(n_3661)
);

AO21x2_ASAP7_75t_L g3662 ( 
.A1(n_3509),
.A2(n_3408),
.B(n_3438),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3456),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3503),
.A2(n_697),
.B1(n_700),
.B2(n_701),
.Y(n_3664)
);

BUFx4f_ASAP7_75t_SL g3665 ( 
.A(n_3325),
.Y(n_3665)
);

AOI22xp5_ASAP7_75t_L g3666 ( 
.A1(n_3363),
.A2(n_701),
.B1(n_702),
.B2(n_703),
.Y(n_3666)
);

AND2x4_ASAP7_75t_L g3667 ( 
.A(n_3392),
.B(n_702),
.Y(n_3667)
);

INVx3_ASAP7_75t_L g3668 ( 
.A(n_3396),
.Y(n_3668)
);

OAI221xp5_ASAP7_75t_SL g3669 ( 
.A1(n_3480),
.A2(n_704),
.B1(n_707),
.B2(n_708),
.C(n_709),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_L g3670 ( 
.A1(n_3425),
.A2(n_704),
.B1(n_707),
.B2(n_708),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3505),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3411),
.Y(n_3672)
);

AOI221xp5_ASAP7_75t_L g3673 ( 
.A1(n_3307),
.A2(n_710),
.B1(n_711),
.B2(n_712),
.C(n_713),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3488),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3369),
.Y(n_3675)
);

BUFx4f_ASAP7_75t_SL g3676 ( 
.A(n_3472),
.Y(n_3676)
);

AOI22xp33_ASAP7_75t_L g3677 ( 
.A1(n_3434),
.A2(n_713),
.B1(n_714),
.B2(n_715),
.Y(n_3677)
);

AOI22xp33_ASAP7_75t_L g3678 ( 
.A1(n_3434),
.A2(n_714),
.B1(n_715),
.B2(n_716),
.Y(n_3678)
);

OR2x2_ASAP7_75t_L g3679 ( 
.A(n_3404),
.B(n_3338),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3397),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3454),
.B(n_774),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_SL g3682 ( 
.A1(n_3347),
.A2(n_716),
.B1(n_717),
.B2(n_718),
.Y(n_3682)
);

AOI222xp33_ASAP7_75t_L g3683 ( 
.A1(n_3427),
.A2(n_717),
.B1(n_719),
.B2(n_721),
.C1(n_722),
.C2(n_723),
.Y(n_3683)
);

AOI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3412),
.A2(n_719),
.B(n_722),
.Y(n_3684)
);

AOI21xp5_ASAP7_75t_L g3685 ( 
.A1(n_3421),
.A2(n_724),
.B(n_725),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3490),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3663),
.Y(n_3687)
);

INVx8_ASAP7_75t_L g3688 ( 
.A(n_3627),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3674),
.Y(n_3689)
);

AND4x1_ASAP7_75t_L g3690 ( 
.A(n_3552),
.B(n_3445),
.C(n_3479),
.D(n_3326),
.Y(n_3690)
);

BUFx2_ASAP7_75t_L g3691 ( 
.A(n_3566),
.Y(n_3691)
);

OAI211xp5_ASAP7_75t_L g3692 ( 
.A1(n_3525),
.A2(n_3543),
.B(n_3551),
.C(n_3516),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3550),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3558),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3574),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3560),
.Y(n_3696)
);

HB1xp67_ASAP7_75t_L g3697 ( 
.A(n_3619),
.Y(n_3697)
);

HB1xp67_ASAP7_75t_L g3698 ( 
.A(n_3564),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3620),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3529),
.B(n_3477),
.Y(n_3700)
);

HB1xp67_ASAP7_75t_L g3701 ( 
.A(n_3533),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3522),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3520),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3572),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3596),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3527),
.B(n_3500),
.Y(n_3706)
);

INVx5_ASAP7_75t_L g3707 ( 
.A(n_3532),
.Y(n_3707)
);

INVx2_ASAP7_75t_SL g3708 ( 
.A(n_3668),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3656),
.Y(n_3709)
);

BUFx12f_ASAP7_75t_L g3710 ( 
.A(n_3595),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3644),
.B(n_3500),
.Y(n_3711)
);

AND2x4_ASAP7_75t_L g3712 ( 
.A(n_3569),
.B(n_3680),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3647),
.B(n_3416),
.Y(n_3713)
);

INVx3_ASAP7_75t_SL g3714 ( 
.A(n_3576),
.Y(n_3714)
);

AOI22xp33_ASAP7_75t_SL g3715 ( 
.A1(n_3528),
.A2(n_3382),
.B1(n_3270),
.B2(n_3442),
.Y(n_3715)
);

INVxp67_ASAP7_75t_L g3716 ( 
.A(n_3617),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3597),
.Y(n_3717)
);

AOI22xp33_ASAP7_75t_SL g3718 ( 
.A1(n_3591),
.A2(n_3416),
.B1(n_3464),
.B2(n_3451),
.Y(n_3718)
);

INVx2_ASAP7_75t_SL g3719 ( 
.A(n_3668),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3547),
.B(n_3320),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3602),
.B(n_3432),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_3567),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3613),
.Y(n_3723)
);

OR2x2_ASAP7_75t_L g3724 ( 
.A(n_3671),
.B(n_3414),
.Y(n_3724)
);

OR2x2_ASAP7_75t_L g3725 ( 
.A(n_3679),
.B(n_3377),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3640),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3625),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3641),
.B(n_3334),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3535),
.B(n_3400),
.Y(n_3729)
);

AND2x2_ASAP7_75t_L g3730 ( 
.A(n_3675),
.B(n_3508),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3650),
.B(n_3342),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3653),
.B(n_3351),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3536),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3536),
.B(n_3378),
.Y(n_3734)
);

AND2x4_ASAP7_75t_L g3735 ( 
.A(n_3569),
.B(n_3403),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3672),
.B(n_3593),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3531),
.B(n_3378),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3555),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3556),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3548),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3577),
.Y(n_3741)
);

AOI22xp33_ASAP7_75t_L g3742 ( 
.A1(n_3540),
.A2(n_3510),
.B1(n_3343),
.B2(n_3344),
.Y(n_3742)
);

INVx4_ASAP7_75t_L g3743 ( 
.A(n_3532),
.Y(n_3743)
);

INVxp67_ASAP7_75t_L g3744 ( 
.A(n_3617),
.Y(n_3744)
);

INVx3_ASAP7_75t_L g3745 ( 
.A(n_3617),
.Y(n_3745)
);

HB1xp67_ASAP7_75t_L g3746 ( 
.A(n_3578),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3563),
.B(n_3312),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3590),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3534),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3530),
.B(n_3366),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3681),
.B(n_3366),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3523),
.B(n_3491),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3524),
.B(n_3507),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3661),
.B(n_3457),
.Y(n_3754)
);

AOI222xp33_ASAP7_75t_L g3755 ( 
.A1(n_3651),
.A2(n_3423),
.B1(n_3324),
.B2(n_3481),
.C1(n_3478),
.C2(n_3447),
.Y(n_3755)
);

OR2x2_ASAP7_75t_L g3756 ( 
.A(n_3571),
.B(n_3493),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3686),
.Y(n_3757)
);

HB1xp67_ASAP7_75t_L g3758 ( 
.A(n_3559),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3587),
.Y(n_3759)
);

BUFx3_ASAP7_75t_L g3760 ( 
.A(n_3646),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3559),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3614),
.Y(n_3762)
);

INVxp67_ASAP7_75t_L g3763 ( 
.A(n_3662),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3568),
.B(n_3513),
.Y(n_3764)
);

OR2x2_ASAP7_75t_L g3765 ( 
.A(n_3635),
.B(n_3349),
.Y(n_3765)
);

OR2x2_ASAP7_75t_SL g3766 ( 
.A(n_3622),
.B(n_3610),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3568),
.B(n_3333),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3524),
.B(n_3373),
.Y(n_3768)
);

OAI22xp5_ASAP7_75t_L g3769 ( 
.A1(n_3643),
.A2(n_3444),
.B1(n_3443),
.B2(n_3379),
.Y(n_3769)
);

NAND4xp25_ASAP7_75t_L g3770 ( 
.A(n_3600),
.B(n_3367),
.C(n_3353),
.D(n_3350),
.Y(n_3770)
);

INVx2_ASAP7_75t_SL g3771 ( 
.A(n_3568),
.Y(n_3771)
);

AND2x4_ASAP7_75t_L g3772 ( 
.A(n_3712),
.B(n_3517),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3725),
.B(n_3553),
.Y(n_3773)
);

OAI33xp33_ASAP7_75t_L g3774 ( 
.A1(n_3696),
.A2(n_3519),
.A3(n_3618),
.B1(n_3623),
.B2(n_3546),
.B3(n_3542),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3701),
.Y(n_3775)
);

INVx1_ASAP7_75t_SL g3776 ( 
.A(n_3714),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3770),
.A2(n_3629),
.B1(n_3592),
.B2(n_3648),
.Y(n_3777)
);

OAI33xp33_ASAP7_75t_L g3778 ( 
.A1(n_3703),
.A2(n_3539),
.A3(n_3609),
.B1(n_3601),
.B2(n_3636),
.B3(n_3549),
.Y(n_3778)
);

NOR2x1p5_ASAP7_75t_L g3779 ( 
.A(n_3760),
.B(n_3595),
.Y(n_3779)
);

NOR2x1_ASAP7_75t_L g3780 ( 
.A(n_3760),
.B(n_3667),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3693),
.Y(n_3781)
);

OAI22xp33_ASAP7_75t_SL g3782 ( 
.A1(n_3691),
.A2(n_3646),
.B1(n_3561),
.B2(n_3667),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3701),
.Y(n_3783)
);

OAI31xp33_ASAP7_75t_SL g3784 ( 
.A1(n_3715),
.A2(n_3608),
.A3(n_3521),
.B(n_3639),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3700),
.B(n_3526),
.Y(n_3785)
);

AOI221xp5_ASAP7_75t_L g3786 ( 
.A1(n_3692),
.A2(n_3604),
.B1(n_3586),
.B2(n_3611),
.C(n_3645),
.Y(n_3786)
);

AO21x2_ASAP7_75t_L g3787 ( 
.A1(n_3763),
.A2(n_3589),
.B(n_3573),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3694),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3757),
.Y(n_3789)
);

AOI221xp5_ASAP7_75t_L g3790 ( 
.A1(n_3720),
.A2(n_3669),
.B1(n_3642),
.B2(n_3654),
.C(n_3537),
.Y(n_3790)
);

AO21x2_ASAP7_75t_L g3791 ( 
.A1(n_3763),
.A2(n_3565),
.B(n_3582),
.Y(n_3791)
);

OAI322xp33_ASAP7_75t_L g3792 ( 
.A1(n_3720),
.A2(n_3753),
.A3(n_3768),
.B1(n_3744),
.B2(n_3716),
.C1(n_3721),
.C2(n_3740),
.Y(n_3792)
);

INVx3_ASAP7_75t_L g3793 ( 
.A(n_3743),
.Y(n_3793)
);

AOI22xp33_ASAP7_75t_L g3794 ( 
.A1(n_3715),
.A2(n_3598),
.B1(n_3683),
.B2(n_3657),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3695),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3687),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3698),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3698),
.B(n_3568),
.Y(n_3798)
);

INVxp67_ASAP7_75t_SL g3799 ( 
.A(n_3758),
.Y(n_3799)
);

INVxp67_ASAP7_75t_SL g3800 ( 
.A(n_3758),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3697),
.B(n_3599),
.Y(n_3801)
);

OAI21xp5_ASAP7_75t_L g3802 ( 
.A1(n_3716),
.A2(n_3682),
.B(n_3658),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3687),
.Y(n_3803)
);

AND2x4_ASAP7_75t_L g3804 ( 
.A(n_3712),
.B(n_3403),
.Y(n_3804)
);

O2A1O1Ixp5_ASAP7_75t_SL g3805 ( 
.A1(n_3697),
.A2(n_3612),
.B(n_3390),
.C(n_3579),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3731),
.B(n_3702),
.Y(n_3806)
);

AOI221xp5_ASAP7_75t_L g3807 ( 
.A1(n_3759),
.A2(n_3673),
.B1(n_3518),
.B2(n_3664),
.C(n_3628),
.Y(n_3807)
);

BUFx3_ASAP7_75t_L g3808 ( 
.A(n_3714),
.Y(n_3808)
);

NAND2xp33_ASAP7_75t_R g3809 ( 
.A(n_3745),
.B(n_3410),
.Y(n_3809)
);

OR2x2_ASAP7_75t_L g3810 ( 
.A(n_3724),
.B(n_3570),
.Y(n_3810)
);

HB1xp67_ASAP7_75t_L g3811 ( 
.A(n_3733),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3744),
.A2(n_3562),
.B1(n_3554),
.B2(n_3652),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3745),
.A2(n_3538),
.B(n_3585),
.Y(n_3813)
);

INVx3_ASAP7_75t_L g3814 ( 
.A(n_3743),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3689),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3699),
.Y(n_3816)
);

HB1xp67_ASAP7_75t_L g3817 ( 
.A(n_3733),
.Y(n_3817)
);

INVxp67_ASAP7_75t_L g3818 ( 
.A(n_3746),
.Y(n_3818)
);

OAI21xp5_ASAP7_75t_L g3819 ( 
.A1(n_3718),
.A2(n_3624),
.B(n_3605),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3689),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3746),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3727),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3729),
.B(n_3541),
.Y(n_3823)
);

AND2x6_ASAP7_75t_SL g3824 ( 
.A(n_3688),
.B(n_3676),
.Y(n_3824)
);

INVxp67_ASAP7_75t_SL g3825 ( 
.A(n_3761),
.Y(n_3825)
);

HB1xp67_ASAP7_75t_L g3826 ( 
.A(n_3704),
.Y(n_3826)
);

HB1xp67_ASAP7_75t_L g3827 ( 
.A(n_3705),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3766),
.A2(n_3678),
.B1(n_3677),
.B2(n_3545),
.Y(n_3828)
);

NOR4xp25_ASAP7_75t_SL g3829 ( 
.A(n_3710),
.B(n_3354),
.C(n_3492),
.D(n_3588),
.Y(n_3829)
);

BUFx3_ASAP7_75t_L g3830 ( 
.A(n_3707),
.Y(n_3830)
);

NAND3xp33_ASAP7_75t_L g3831 ( 
.A(n_3718),
.B(n_3690),
.C(n_3755),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3709),
.Y(n_3832)
);

AOI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_3742),
.A2(n_3638),
.B1(n_3632),
.B2(n_3649),
.Y(n_3833)
);

OAI21x1_ASAP7_75t_L g3834 ( 
.A1(n_3745),
.A2(n_3557),
.B(n_3761),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3738),
.Y(n_3835)
);

BUFx3_ASAP7_75t_L g3836 ( 
.A(n_3707),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3706),
.B(n_3713),
.Y(n_3837)
);

AND2x4_ASAP7_75t_L g3838 ( 
.A(n_3772),
.B(n_3735),
.Y(n_3838)
);

INVx3_ASAP7_75t_L g3839 ( 
.A(n_3830),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3823),
.B(n_3741),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3837),
.B(n_3712),
.Y(n_3841)
);

OR2x2_ASAP7_75t_L g3842 ( 
.A(n_3821),
.B(n_3749),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3811),
.B(n_3736),
.Y(n_3843)
);

NOR2xp33_ASAP7_75t_L g3844 ( 
.A(n_3808),
.B(n_3688),
.Y(n_3844)
);

OR2x2_ASAP7_75t_L g3845 ( 
.A(n_3821),
.B(n_3752),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3773),
.B(n_3739),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3826),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3826),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3811),
.B(n_3750),
.Y(n_3849)
);

OR2x2_ASAP7_75t_L g3850 ( 
.A(n_3797),
.B(n_3756),
.Y(n_3850)
);

HB1xp67_ASAP7_75t_L g3851 ( 
.A(n_3817),
.Y(n_3851)
);

HB1xp67_ASAP7_75t_L g3852 ( 
.A(n_3817),
.Y(n_3852)
);

HB1xp67_ASAP7_75t_L g3853 ( 
.A(n_3827),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3818),
.B(n_3737),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3827),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3799),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3818),
.B(n_3728),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_3772),
.B(n_3735),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3806),
.B(n_3711),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3810),
.B(n_3734),
.Y(n_3860)
);

OR2x2_ASAP7_75t_L g3861 ( 
.A(n_3775),
.B(n_3748),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3799),
.Y(n_3862)
);

HB1xp67_ASAP7_75t_L g3863 ( 
.A(n_3783),
.Y(n_3863)
);

HB1xp67_ASAP7_75t_L g3864 ( 
.A(n_3800),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3798),
.B(n_3754),
.Y(n_3865)
);

INVx3_ASAP7_75t_L g3866 ( 
.A(n_3830),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3800),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3832),
.B(n_3835),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3825),
.B(n_3764),
.Y(n_3869)
);

AND2x4_ASAP7_75t_L g3870 ( 
.A(n_3779),
.B(n_3735),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3822),
.B(n_3762),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3825),
.B(n_3732),
.Y(n_3872)
);

NOR2x1_ASAP7_75t_L g3873 ( 
.A(n_3808),
.B(n_3743),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3789),
.Y(n_3874)
);

AND2x4_ASAP7_75t_L g3875 ( 
.A(n_3793),
.B(n_3708),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3785),
.B(n_3730),
.Y(n_3876)
);

OR2x2_ASAP7_75t_L g3877 ( 
.A(n_3801),
.B(n_3803),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3815),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3781),
.B(n_3788),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3820),
.Y(n_3880)
);

INVxp67_ASAP7_75t_L g3881 ( 
.A(n_3776),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3796),
.Y(n_3882)
);

BUFx2_ASAP7_75t_L g3883 ( 
.A(n_3836),
.Y(n_3883)
);

NAND4xp25_ASAP7_75t_L g3884 ( 
.A(n_3784),
.B(n_3742),
.C(n_3769),
.D(n_3544),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3795),
.B(n_3816),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3834),
.B(n_3717),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3791),
.B(n_3723),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3791),
.B(n_3723),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3842),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3860),
.B(n_3831),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3872),
.Y(n_3891)
);

AOI32xp33_ASAP7_75t_L g3892 ( 
.A1(n_3873),
.A2(n_3780),
.A3(n_3828),
.B1(n_3777),
.B2(n_3812),
.Y(n_3892)
);

OR2x2_ASAP7_75t_L g3893 ( 
.A(n_3845),
.B(n_3726),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3872),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3842),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3845),
.Y(n_3896)
);

NOR2x1_ASAP7_75t_L g3897 ( 
.A(n_3873),
.B(n_3793),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3877),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3877),
.Y(n_3899)
);

AND2x2_ASAP7_75t_SL g3900 ( 
.A(n_3870),
.B(n_3814),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3870),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3885),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3849),
.B(n_3787),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3860),
.B(n_3767),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3853),
.Y(n_3905)
);

AOI21xp33_ASAP7_75t_L g3906 ( 
.A1(n_3881),
.A2(n_3819),
.B(n_3777),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3854),
.B(n_3813),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3849),
.B(n_3787),
.Y(n_3908)
);

BUFx2_ASAP7_75t_L g3909 ( 
.A(n_3883),
.Y(n_3909)
);

INVxp67_ASAP7_75t_L g3910 ( 
.A(n_3864),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3855),
.Y(n_3911)
);

OR2x2_ASAP7_75t_L g3912 ( 
.A(n_3846),
.B(n_3726),
.Y(n_3912)
);

NAND2x1p5_ASAP7_75t_L g3913 ( 
.A(n_3883),
.B(n_3814),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3854),
.B(n_3765),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3885),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3840),
.B(n_3790),
.Y(n_3916)
);

HB1xp67_ASAP7_75t_L g3917 ( 
.A(n_3851),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3868),
.Y(n_3918)
);

INVxp67_ASAP7_75t_SL g3919 ( 
.A(n_3852),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3868),
.Y(n_3920)
);

OR2x2_ASAP7_75t_L g3921 ( 
.A(n_3857),
.B(n_3850),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3861),
.Y(n_3922)
);

NAND4xp25_ASAP7_75t_SL g3923 ( 
.A(n_3884),
.B(n_3794),
.C(n_3833),
.D(n_3802),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3843),
.B(n_3782),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3857),
.B(n_3708),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3916),
.B(n_3843),
.Y(n_3926)
);

NAND2xp33_ASAP7_75t_SL g3927 ( 
.A(n_3909),
.B(n_3839),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3921),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3917),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3917),
.Y(n_3930)
);

NOR3xp33_ASAP7_75t_L g3931 ( 
.A(n_3923),
.B(n_3774),
.C(n_3778),
.Y(n_3931)
);

NAND2xp33_ASAP7_75t_R g3932 ( 
.A(n_3901),
.B(n_3829),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3900),
.B(n_3901),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3891),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3902),
.Y(n_3935)
);

NAND2xp33_ASAP7_75t_SL g3936 ( 
.A(n_3901),
.B(n_3839),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3890),
.B(n_3859),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3907),
.B(n_3859),
.Y(n_3938)
);

AOI22xp5_ASAP7_75t_L g3939 ( 
.A1(n_3906),
.A2(n_3809),
.B1(n_3794),
.B2(n_3844),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3915),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3900),
.B(n_3838),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3896),
.B(n_3856),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3891),
.Y(n_3943)
);

INVx1_ASAP7_75t_SL g3944 ( 
.A(n_3913),
.Y(n_3944)
);

AOI221xp5_ASAP7_75t_L g3945 ( 
.A1(n_3892),
.A2(n_3792),
.B1(n_3871),
.B2(n_3786),
.C(n_3833),
.Y(n_3945)
);

NOR2xp33_ASAP7_75t_R g3946 ( 
.A(n_3924),
.B(n_3824),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3894),
.B(n_3903),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3894),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3903),
.B(n_3865),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3918),
.Y(n_3950)
);

AOI21xp33_ASAP7_75t_L g3951 ( 
.A1(n_3910),
.A2(n_3888),
.B(n_3887),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3911),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3920),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3908),
.B(n_3914),
.Y(n_3954)
);

AND2x2_ASAP7_75t_SL g3955 ( 
.A(n_3908),
.B(n_3870),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3912),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3910),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3914),
.B(n_3904),
.Y(n_3958)
);

NOR2x1_ASAP7_75t_L g3959 ( 
.A(n_3897),
.B(n_3839),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3889),
.B(n_3865),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3895),
.A2(n_3710),
.B1(n_3807),
.B2(n_3887),
.Y(n_3961)
);

AND2x2_ASAP7_75t_L g3962 ( 
.A(n_3922),
.B(n_3841),
.Y(n_3962)
);

NOR2xp33_ASAP7_75t_L g3963 ( 
.A(n_3919),
.B(n_3879),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3927),
.A2(n_3688),
.B(n_3913),
.Y(n_3964)
);

INVx2_ASAP7_75t_SL g3965 ( 
.A(n_3946),
.Y(n_3965)
);

OAI22xp5_ASAP7_75t_L g3966 ( 
.A1(n_3939),
.A2(n_3919),
.B1(n_3866),
.B2(n_3925),
.Y(n_3966)
);

AOI321xp33_ASAP7_75t_L g3967 ( 
.A1(n_3931),
.A2(n_3888),
.A3(n_3905),
.B1(n_3867),
.B2(n_3862),
.C(n_3856),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3929),
.Y(n_3968)
);

OR2x2_ASAP7_75t_L g3969 ( 
.A(n_3928),
.B(n_3898),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3941),
.B(n_3899),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3952),
.Y(n_3971)
);

OA21x2_ASAP7_75t_L g3972 ( 
.A1(n_3957),
.A2(n_3905),
.B(n_3867),
.Y(n_3972)
);

OR2x2_ASAP7_75t_L g3973 ( 
.A(n_3926),
.B(n_3893),
.Y(n_3973)
);

AOI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3945),
.A2(n_3751),
.B1(n_3862),
.B2(n_3886),
.Y(n_3974)
);

OAI21xp33_ASAP7_75t_SL g3975 ( 
.A1(n_3955),
.A2(n_3841),
.B(n_3876),
.Y(n_3975)
);

INVx3_ASAP7_75t_L g3976 ( 
.A(n_3933),
.Y(n_3976)
);

XOR2x2_ASAP7_75t_L g3977 ( 
.A(n_3961),
.B(n_3339),
.Y(n_3977)
);

NAND3xp33_ASAP7_75t_L g3978 ( 
.A(n_3927),
.B(n_3805),
.C(n_3886),
.Y(n_3978)
);

AOI211xp5_ASAP7_75t_L g3979 ( 
.A1(n_3946),
.A2(n_3858),
.B(n_3838),
.C(n_3866),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3952),
.Y(n_3980)
);

OAI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3944),
.A2(n_3809),
.B1(n_3866),
.B2(n_3836),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3930),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3956),
.Y(n_3983)
);

NOR3xp33_ASAP7_75t_L g3984 ( 
.A(n_3936),
.B(n_3655),
.C(n_3660),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3934),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3955),
.B(n_3838),
.Y(n_3986)
);

INVx1_ASAP7_75t_SL g3987 ( 
.A(n_3936),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3942),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3935),
.B(n_3911),
.Y(n_3989)
);

AOI21xp33_ASAP7_75t_L g3990 ( 
.A1(n_3932),
.A2(n_3306),
.B(n_724),
.Y(n_3990)
);

AOI222xp33_ASAP7_75t_L g3991 ( 
.A1(n_3966),
.A2(n_3961),
.B1(n_3963),
.B2(n_3937),
.C1(n_3954),
.C2(n_3947),
.Y(n_3991)
);

OAI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3979),
.A2(n_3938),
.B1(n_3959),
.B2(n_3949),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3965),
.B(n_3958),
.Y(n_3993)
);

INVx2_ASAP7_75t_SL g3994 ( 
.A(n_3977),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3969),
.Y(n_3995)
);

OAI21xp33_ASAP7_75t_L g3996 ( 
.A1(n_3990),
.A2(n_3974),
.B(n_3966),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3973),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3988),
.B(n_3963),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3986),
.B(n_3949),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3983),
.Y(n_4000)
);

CKINVDCx14_ASAP7_75t_R g4001 ( 
.A(n_3976),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3972),
.Y(n_4002)
);

AOI222xp33_ASAP7_75t_L g4003 ( 
.A1(n_3974),
.A2(n_3987),
.B1(n_3968),
.B2(n_3982),
.C1(n_3978),
.C2(n_3976),
.Y(n_4003)
);

INVxp67_ASAP7_75t_L g4004 ( 
.A(n_3990),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3970),
.Y(n_4005)
);

AOI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_3984),
.A2(n_3932),
.B1(n_3950),
.B2(n_3940),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3989),
.Y(n_4007)
);

AOI322xp5_ASAP7_75t_L g4008 ( 
.A1(n_3975),
.A2(n_3960),
.A3(n_3951),
.B1(n_3962),
.B2(n_3953),
.C1(n_3948),
.C2(n_3943),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3964),
.B(n_3960),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3964),
.A2(n_3943),
.B(n_3934),
.Y(n_4010)
);

OR2x2_ASAP7_75t_L g4011 ( 
.A(n_3989),
.B(n_3948),
.Y(n_4011)
);

OAI21xp33_ASAP7_75t_L g4012 ( 
.A1(n_3996),
.A2(n_3984),
.B(n_3981),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3993),
.Y(n_4013)
);

XOR2xp5_ASAP7_75t_L g4014 ( 
.A(n_4001),
.B(n_3318),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_4002),
.Y(n_4015)
);

NOR2x1_ASAP7_75t_L g4016 ( 
.A(n_4000),
.B(n_3981),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_4011),
.Y(n_4017)
);

NAND4xp25_ASAP7_75t_L g4018 ( 
.A(n_4006),
.B(n_3967),
.C(n_3606),
.D(n_3626),
.Y(n_4018)
);

OAI221xp5_ASAP7_75t_SL g4019 ( 
.A1(n_3996),
.A2(n_3985),
.B1(n_3980),
.B2(n_3971),
.C(n_3666),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_4009),
.B(n_3999),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3997),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3994),
.B(n_3962),
.Y(n_4022)
);

XOR2x2_ASAP7_75t_L g4023 ( 
.A(n_4006),
.B(n_3998),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_4005),
.B(n_3972),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3995),
.Y(n_4025)
);

OAI221xp5_ASAP7_75t_L g4026 ( 
.A1(n_4010),
.A2(n_3621),
.B1(n_3603),
.B2(n_3670),
.C(n_3616),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_4007),
.Y(n_4027)
);

NOR2xp33_ASAP7_75t_L g4028 ( 
.A(n_4004),
.B(n_3665),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_4003),
.B(n_3876),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3992),
.B(n_3417),
.Y(n_4030)
);

O2A1O1Ixp33_ASAP7_75t_L g4031 ( 
.A1(n_4012),
.A2(n_3991),
.B(n_4008),
.C(n_3470),
.Y(n_4031)
);

NOR4xp25_ASAP7_75t_L g4032 ( 
.A(n_4012),
.B(n_4027),
.C(n_4019),
.D(n_4021),
.Y(n_4032)
);

XOR2x2_ASAP7_75t_L g4033 ( 
.A(n_4014),
.B(n_3838),
.Y(n_4033)
);

XNOR2x1_ASAP7_75t_L g4034 ( 
.A(n_4023),
.B(n_3858),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_4020),
.B(n_3847),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_4015),
.Y(n_4036)
);

NOR2x1_ASAP7_75t_L g4037 ( 
.A(n_4028),
.B(n_3607),
.Y(n_4037)
);

INVxp67_ASAP7_75t_L g4038 ( 
.A(n_4013),
.Y(n_4038)
);

NOR2x1_ASAP7_75t_L g4039 ( 
.A(n_4016),
.B(n_3607),
.Y(n_4039)
);

NOR3x1_ASAP7_75t_L g4040 ( 
.A(n_4018),
.B(n_3389),
.C(n_3847),
.Y(n_4040)
);

AOI211xp5_ASAP7_75t_SL g4041 ( 
.A1(n_4030),
.A2(n_3684),
.B(n_3685),
.C(n_3858),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_4022),
.B(n_3848),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_4017),
.B(n_3848),
.Y(n_4043)
);

O2A1O1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_4036),
.A2(n_4025),
.B(n_4029),
.C(n_4018),
.Y(n_4044)
);

OAI21xp33_ASAP7_75t_SL g4045 ( 
.A1(n_4034),
.A2(n_4024),
.B(n_4026),
.Y(n_4045)
);

NAND4xp25_ASAP7_75t_L g4046 ( 
.A(n_4031),
.B(n_3637),
.C(n_3633),
.D(n_3634),
.Y(n_4046)
);

NAND4xp25_ASAP7_75t_L g4047 ( 
.A(n_4038),
.B(n_3631),
.C(n_3659),
.D(n_3858),
.Y(n_4047)
);

AOI221x1_ASAP7_75t_SL g4048 ( 
.A1(n_4032),
.A2(n_3875),
.B1(n_3855),
.B2(n_3580),
.C(n_3882),
.Y(n_4048)
);

OAI21xp5_ASAP7_75t_SL g4049 ( 
.A1(n_4041),
.A2(n_3875),
.B(n_3804),
.Y(n_4049)
);

AOI221xp5_ASAP7_75t_L g4050 ( 
.A1(n_4043),
.A2(n_3594),
.B1(n_3875),
.B2(n_3863),
.C(n_3358),
.Y(n_4050)
);

NAND4xp25_ASAP7_75t_L g4051 ( 
.A(n_4040),
.B(n_3804),
.C(n_3581),
.D(n_3747),
.Y(n_4051)
);

AOI211xp5_ASAP7_75t_L g4052 ( 
.A1(n_4035),
.A2(n_3380),
.B(n_3394),
.C(n_3630),
.Y(n_4052)
);

OAI22xp5_ASAP7_75t_L g4053 ( 
.A1(n_4042),
.A2(n_3861),
.B1(n_3850),
.B2(n_3707),
.Y(n_4053)
);

INVxp67_ASAP7_75t_L g4054 ( 
.A(n_4046),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_4044),
.A2(n_4039),
.B(n_4033),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_SL g4056 ( 
.A(n_4049),
.B(n_4037),
.Y(n_4056)
);

INVx1_ASAP7_75t_SL g4057 ( 
.A(n_4053),
.Y(n_4057)
);

AOI211x1_ASAP7_75t_L g4058 ( 
.A1(n_4048),
.A2(n_3869),
.B(n_3882),
.C(n_3880),
.Y(n_4058)
);

OAI221xp5_ASAP7_75t_SL g4059 ( 
.A1(n_4057),
.A2(n_4045),
.B1(n_4050),
.B2(n_4051),
.C(n_4047),
.Y(n_4059)
);

AOI221xp5_ASAP7_75t_L g4060 ( 
.A1(n_4055),
.A2(n_4054),
.B1(n_4058),
.B2(n_4056),
.C(n_4052),
.Y(n_4060)
);

CKINVDCx5p33_ASAP7_75t_R g4061 ( 
.A(n_4057),
.Y(n_4061)
);

NOR2xp33_ASAP7_75t_L g4062 ( 
.A(n_4057),
.B(n_3302),
.Y(n_4062)
);

NAND2x1p5_ASAP7_75t_L g4063 ( 
.A(n_4057),
.B(n_3707),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_4061),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4063),
.Y(n_4065)
);

AOI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_4062),
.A2(n_3615),
.B1(n_3869),
.B2(n_3512),
.Y(n_4066)
);

NAND3xp33_ASAP7_75t_SL g4067 ( 
.A(n_4060),
.B(n_3415),
.C(n_3584),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_4064),
.B(n_4059),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_4065),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4069),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_4070),
.A2(n_4068),
.B1(n_4067),
.B2(n_4066),
.Y(n_4071)
);

OAI22xp5_ASAP7_75t_SL g4072 ( 
.A1(n_4070),
.A2(n_3567),
.B1(n_3401),
.B2(n_3719),
.Y(n_4072)
);

BUFx2_ASAP7_75t_L g4073 ( 
.A(n_4072),
.Y(n_4073)
);

AOI222xp33_ASAP7_75t_L g4074 ( 
.A1(n_4073),
.A2(n_4071),
.B1(n_3615),
.B2(n_3880),
.C1(n_3874),
.C2(n_3878),
.Y(n_4074)
);

AOI22xp33_ASAP7_75t_L g4075 ( 
.A1(n_4074),
.A2(n_3719),
.B1(n_3722),
.B2(n_3878),
.Y(n_4075)
);

AOI22xp5_ASAP7_75t_SL g4076 ( 
.A1(n_4075),
.A2(n_3771),
.B1(n_3482),
.B2(n_3461),
.Y(n_4076)
);

OAI221xp5_ASAP7_75t_R g4077 ( 
.A1(n_4076),
.A2(n_3337),
.B1(n_3428),
.B2(n_3583),
.C(n_3575),
.Y(n_4077)
);

AOI211xp5_ASAP7_75t_L g4078 ( 
.A1(n_4077),
.A2(n_3722),
.B(n_3469),
.C(n_3496),
.Y(n_4078)
);


endmodule