module fake_jpeg_3018_n_63 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_63);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_23),
.B(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_28),
.B1(n_24),
.B2(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_19),
.B1(n_18),
.B2(n_25),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_28),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_31),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_34),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_23),
.C(n_20),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_22),
.B(n_41),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_1),
.C(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_36),
.B1(n_33),
.B2(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_6),
.C(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_5),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_56),
.B1(n_7),
.B2(n_8),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_50),
.B(n_48),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.C(n_55),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_8),
.Y(n_62)
);

NAND4xp25_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_9),
.C(n_10),
.D(n_21),
.Y(n_63)
);


endmodule