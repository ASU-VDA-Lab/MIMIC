module fake_jpeg_32001_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_14),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_0),
.B(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_53),
.Y(n_94)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_87),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_53),
.B(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_56),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_52),
.B1(n_54),
.B2(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_57),
.B1(n_69),
.B2(n_70),
.Y(n_101)
);

AO22x2_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_71),
.B1(n_58),
.B2(n_67),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_71),
.B1(n_67),
.B2(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_1),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_111),
.Y(n_118)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_51),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_101),
.B1(n_110),
.B2(n_49),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_64),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_66),
.B(n_71),
.C(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_1),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_61),
.B1(n_83),
.B2(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_18),
.B1(n_36),
.B2(n_35),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_21),
.B1(n_47),
.B2(n_43),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_131),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_20),
.C(n_39),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_19),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_22),
.C(n_37),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_6),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_17),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_111),
.C(n_96),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_24),
.B(n_33),
.C(n_32),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_138),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_127),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_139),
.A2(n_145),
.B(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_13),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_124),
.C(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_129),
.B(n_118),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_150),
.C(n_136),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.C(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_136),
.C(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_138),
.Y(n_156)
);

XNOR2x2_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_135),
.C(n_152),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_140),
.A3(n_29),
.B1(n_25),
.B2(n_27),
.C1(n_28),
.C2(n_40),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_31),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_14),
.Y(n_162)
);


endmodule