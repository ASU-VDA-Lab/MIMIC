module fake_jpeg_5486_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_51),
.Y(n_80)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_57),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_18),
.B1(n_31),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_67),
.B1(n_29),
.B2(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_31),
.B1(n_34),
.B2(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_76),
.Y(n_110)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_45),
.B1(n_41),
.B2(n_48),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_39),
.B1(n_66),
.B2(n_30),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_45),
.B1(n_48),
.B2(n_40),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_66),
.B1(n_63),
.B2(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_87),
.Y(n_119)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_20),
.Y(n_122)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_31),
.B1(n_34),
.B2(n_17),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_97),
.B1(n_33),
.B2(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_40),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_43),
.A3(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_39),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_126),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_107),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_43),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_85),
.C(n_78),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_126),
.B1(n_74),
.B2(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_74),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_93),
.B1(n_99),
.B2(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_26),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_20),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_26),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_35),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_132),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_136),
.B1(n_150),
.B2(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_72),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_96),
.B1(n_77),
.B2(n_93),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_134),
.A2(n_141),
.B1(n_75),
.B2(n_123),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_27),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_71),
.B1(n_90),
.B2(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_85),
.B1(n_78),
.B2(n_88),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_27),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_19),
.Y(n_184)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_84),
.B(n_23),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_115),
.B(n_127),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_94),
.B(n_32),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_123),
.B(n_112),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_23),
.C(n_25),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_158),
.B(n_23),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_110),
.B1(n_103),
.B2(n_107),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_115),
.B1(n_111),
.B2(n_104),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_25),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_162),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_170),
.B1(n_190),
.B2(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_32),
.B(n_112),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_175),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_114),
.B1(n_32),
.B2(n_86),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_181),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_177),
.C(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_39),
.B1(n_111),
.B2(n_55),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_19),
.B(n_27),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_104),
.C(n_100),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_63),
.C(n_55),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_27),
.B(n_19),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_36),
.B1(n_24),
.B2(n_22),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_189),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_63),
.C(n_19),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_187),
.C(n_131),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_27),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_19),
.B(n_30),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_22),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_19),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_130),
.Y(n_213)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_141),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_197),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_135),
.B1(n_132),
.B2(n_151),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_210),
.B1(n_179),
.B2(n_174),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_36),
.B(n_24),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_216),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_160),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_207),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_212),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_162),
.A2(n_154),
.B1(n_152),
.B2(n_157),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_164),
.A2(n_168),
.B1(n_161),
.B2(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_22),
.B1(n_30),
.B2(n_36),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_221),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_222),
.C(n_178),
.Y(n_223)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

AO221x1_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_176),
.B1(n_186),
.B2(n_175),
.C(n_189),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_142),
.A3(n_158),
.B1(n_137),
.B2(n_22),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_142),
.C(n_150),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_227),
.C(n_233),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_225),
.A2(n_235),
.B1(n_236),
.B2(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_177),
.C(n_183),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_218),
.C(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_176),
.B1(n_185),
.B2(n_187),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_183),
.B1(n_163),
.B2(n_191),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_221),
.B1(n_15),
.B2(n_14),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_156),
.C(n_19),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_245),
.C(n_246),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_156),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_209),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_202),
.B1(n_220),
.B2(n_203),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_30),
.B1(n_36),
.B2(n_24),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_30),
.C(n_24),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_0),
.C(n_1),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_210),
.C(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_259),
.C(n_223),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_200),
.C(n_204),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_263),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_15),
.C(n_13),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_13),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_239),
.Y(n_277)
);

AO22x1_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_260),
.B1(n_254),
.B2(n_229),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_226),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_272),
.C(n_249),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_255),
.C(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_238),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_287),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_248),
.B(n_259),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_282),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_225),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_235),
.B1(n_248),
.B2(n_240),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_269),
.B1(n_268),
.B2(n_253),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_296),
.C(n_299),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_250),
.C(n_246),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_266),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_10),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_250),
.C(n_262),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_274),
.B(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_285),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_0),
.C(n_2),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_273),
.C(n_281),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_280),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_306),
.C(n_308),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_287),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_312),
.B(n_314),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_286),
.C(n_283),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_279),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_311),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_293),
.B(n_10),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_6),
.B(n_7),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_295),
.B(n_0),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_2),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_9),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_289),
.B(n_302),
.C(n_5),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_323),
.B(n_313),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_324),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_9),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_325),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.C(n_330),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_309),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_323),
.B(n_8),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_326),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_333),
.B(n_332),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_327),
.Y(n_337)
);

OAI31xp33_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_6),
.A3(n_8),
.B(n_9),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_6),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_8),
.B(n_323),
.Y(n_340)
);


endmodule