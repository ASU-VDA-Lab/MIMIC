module fake_jpeg_13743_n_601 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_601);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_60),
.Y(n_203)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_66),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_67),
.B(n_81),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_44),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_75),
.Y(n_144)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_32),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_82),
.B(n_83),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_1),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_85),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_87),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_21),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_91),
.B(n_100),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_92),
.Y(n_213)
);

HAxp5_ASAP7_75t_SL g93 ( 
.A(n_29),
.B(n_1),
.CON(n_93),
.SN(n_93)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_93),
.B(n_6),
.Y(n_215)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_4),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_23),
.B(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_103),
.B(n_105),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_23),
.B(n_4),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_108),
.B(n_123),
.Y(n_197)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_24),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_125),
.Y(n_178)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_34),
.B(n_4),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_35),
.B(n_5),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_60),
.A2(n_49),
.B1(n_52),
.B2(n_56),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_138),
.A2(n_205),
.B(n_24),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_67),
.B(n_33),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_139),
.B(n_156),
.Y(n_236)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_58),
.B1(n_54),
.B2(n_39),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_152),
.A2(n_167),
.B1(n_185),
.B2(n_201),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_33),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_36),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_160),
.B(n_208),
.Y(n_290)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_58),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_187),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_104),
.A2(n_31),
.B1(n_56),
.B2(n_55),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_59),
.Y(n_174)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_176),
.Y(n_254)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_84),
.Y(n_182)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_182),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_113),
.A2(n_54),
.B1(n_39),
.B2(n_57),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_78),
.B(n_28),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_79),
.Y(n_191)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_195),
.Y(n_286)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_68),
.Y(n_199)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_74),
.A2(n_57),
.B1(n_55),
.B2(n_31),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_98),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_204),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_112),
.A2(n_52),
.B1(n_49),
.B2(n_48),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_85),
.B(n_42),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_43),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_93),
.B(n_42),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_11),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_6),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_220),
.B(n_252),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_120),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_119),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_222),
.C(n_242),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_40),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_167),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_223),
.A2(n_228),
.B1(n_244),
.B2(n_260),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_225),
.B(n_235),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_36),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_227),
.B(n_277),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_89),
.B1(n_92),
.B2(n_48),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_144),
.A2(n_40),
.B1(n_43),
.B2(n_37),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_237),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_37),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_239),
.B(n_258),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_241),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_128),
.B(n_108),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_135),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_243),
.B(n_271),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_178),
.A2(n_75),
.B1(n_96),
.B2(n_66),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_155),
.Y(n_246)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_248),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_137),
.B(n_149),
.C(n_142),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_253),
.Y(n_315)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_158),
.Y(n_251)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_129),
.B(n_52),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_131),
.B(n_52),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_153),
.A2(n_52),
.B1(n_49),
.B2(n_24),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_255),
.A2(n_261),
.B1(n_272),
.B2(n_288),
.Y(n_303)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_256),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_193),
.B(n_49),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g259 ( 
.A(n_145),
.Y(n_259)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_259),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_157),
.A2(n_24),
.B1(n_7),
.B2(n_9),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_163),
.A2(n_172),
.B1(n_205),
.B2(n_138),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_132),
.B(n_6),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

AOI32xp33_ASAP7_75t_L g264 ( 
.A1(n_163),
.A2(n_24),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_264),
.B(n_214),
.CI(n_141),
.CON(n_309),
.SN(n_309)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

BUFx8_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_216),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_133),
.A2(n_17),
.B1(n_12),
.B2(n_13),
.Y(n_272)
);

OR2x4_ASAP7_75t_L g273 ( 
.A(n_134),
.B(n_11),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_273),
.A2(n_218),
.B(n_242),
.C(n_253),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_140),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_274),
.A2(n_278),
.B1(n_259),
.B2(n_287),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_275),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_144),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_143),
.B(n_14),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_170),
.A2(n_15),
.B1(n_17),
.B2(n_196),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_147),
.Y(n_282)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_172),
.B(n_173),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_283),
.B(n_273),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_184),
.Y(n_324)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_159),
.Y(n_285)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_151),
.A2(n_206),
.B1(n_181),
.B2(n_141),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_287),
.A2(n_278),
.B1(n_269),
.B2(n_217),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_190),
.A2(n_207),
.B1(n_198),
.B2(n_188),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_305),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_242),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_309),
.B(n_313),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_255),
.A2(n_213),
.B1(n_179),
.B2(n_200),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_311),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_226),
.B(n_175),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_202),
.B1(n_162),
.B2(n_130),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_227),
.B(n_164),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_337),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_257),
.A2(n_171),
.B1(n_169),
.B2(n_186),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_265),
.A2(n_184),
.B1(n_188),
.B2(n_272),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_222),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_325),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_220),
.A2(n_265),
.B1(n_277),
.B2(n_262),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_220),
.A2(n_277),
.B1(n_262),
.B2(n_218),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_331),
.Y(n_365)
);

NOR3xp33_ASAP7_75t_SL g337 ( 
.A(n_236),
.B(n_271),
.C(n_270),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_217),
.A2(n_266),
.B1(n_249),
.B2(n_291),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_346),
.B(n_314),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_221),
.B(n_285),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_320),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_231),
.Y(n_346)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_346),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_281),
.B1(n_282),
.B2(n_263),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_252),
.C(n_253),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_349),
.B(n_353),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_252),
.C(n_234),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_347),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_354),
.B(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_334),
.A2(n_230),
.B1(n_256),
.B2(n_251),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_322),
.A2(n_219),
.B(n_238),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_358),
.A2(n_368),
.B(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_303),
.A2(n_274),
.B1(n_280),
.B2(n_254),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_371),
.B1(n_372),
.B2(n_382),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_286),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_362),
.B(n_343),
.Y(n_404)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_366),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_295),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_232),
.B(n_229),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_334),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_369),
.A2(n_370),
.B1(n_383),
.B2(n_345),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_303),
.A2(n_224),
.B1(n_233),
.B2(n_247),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_326),
.A2(n_268),
.B1(n_279),
.B2(n_284),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_267),
.B1(n_284),
.B2(n_304),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_374),
.A2(n_387),
.B1(n_302),
.B2(n_318),
.Y(n_420)
);

FAx1_ASAP7_75t_SL g375 ( 
.A(n_300),
.B(n_339),
.CI(n_294),
.CON(n_375),
.SN(n_375)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_375),
.B(n_317),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_377),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_294),
.B(n_328),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_306),
.A2(n_331),
.B(n_328),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_313),
.B(n_327),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_384),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_306),
.A2(n_309),
.B1(n_311),
.B2(n_333),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_307),
.A2(n_342),
.B1(n_297),
.B2(n_293),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_310),
.B(n_309),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_312),
.A2(n_296),
.B1(n_297),
.B2(n_341),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_316),
.A2(n_330),
.B1(n_332),
.B2(n_337),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_342),
.B1(n_293),
.B2(n_308),
.Y(n_398)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_341),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_376),
.Y(n_423)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_301),
.C(n_307),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_343),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_390),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_393),
.B(n_407),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_398),
.A2(n_412),
.B1(n_422),
.B2(n_389),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_332),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_399),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_392),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_400),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_308),
.C(n_330),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_403),
.C(n_419),
.Y(n_461)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_343),
.C(n_317),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_425),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_299),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_408),
.B(n_417),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_420),
.B1(n_381),
.B2(n_373),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_318),
.B1(n_345),
.B2(n_302),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_354),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_413),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_391),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_292),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_418),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_378),
.A2(n_292),
.B(n_299),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_421),
.A2(n_368),
.B(n_358),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_371),
.B1(n_365),
.B2(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_377),
.B(n_375),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_359),
.Y(n_427)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_428),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_353),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_446),
.C(n_455),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_422),
.A2(n_384),
.B1(n_387),
.B2(n_374),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_433),
.A2(n_445),
.B1(n_449),
.B2(n_450),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_436),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_365),
.B1(n_381),
.B2(n_372),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_437),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_424),
.A2(n_365),
.B1(n_373),
.B2(n_386),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_457),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_349),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g474 ( 
.A1(n_440),
.A2(n_398),
.B(n_405),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_403),
.Y(n_442)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

BUFx5_ASAP7_75t_L g443 ( 
.A(n_426),
.Y(n_443)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_370),
.B1(n_389),
.B2(n_379),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_375),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_394),
.A2(n_389),
.B1(n_386),
.B2(n_352),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_414),
.A2(n_389),
.B1(n_355),
.B2(n_357),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_451),
.A2(n_452),
.B1(n_453),
.B2(n_410),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_402),
.A2(n_351),
.B1(n_360),
.B2(n_363),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_402),
.A2(n_351),
.B1(n_364),
.B2(n_400),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_454),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_404),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_416),
.B1(n_408),
.B2(n_414),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_458),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_416),
.A2(n_407),
.B(n_395),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_428),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_421),
.A2(n_395),
.B(n_409),
.Y(n_460)
);

AOI21xp33_ASAP7_75t_L g466 ( 
.A1(n_460),
.A2(n_413),
.B(n_417),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_419),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_464),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_401),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_465),
.B(n_482),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_466),
.B(n_487),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_423),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_469),
.B(n_474),
.Y(n_500)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_454),
.Y(n_470)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_470),
.Y(n_503)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_475),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_405),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_484),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_410),
.C(n_415),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_483),
.C(n_432),
.Y(n_492)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_432),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_431),
.B(n_415),
.C(n_426),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_412),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_397),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_474),
.Y(n_516)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_486),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_447),
.B(n_397),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_489),
.Y(n_499)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_443),
.Y(n_490)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_490),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_504),
.C(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_444),
.Y(n_494)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_480),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_496),
.B(n_463),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_444),
.Y(n_502)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_462),
.B(n_461),
.C(n_431),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_461),
.C(n_440),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_442),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_509),
.B(n_485),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_471),
.B(n_457),
.C(n_439),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_511),
.C(n_515),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_438),
.C(n_437),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_469),
.C(n_484),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_516),
.B(n_481),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_463),
.A2(n_456),
.B1(n_435),
.B2(n_436),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_473),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_502),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_527),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_505),
.Y(n_519)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_519),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_531),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_525),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_474),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_533),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_498),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_529),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_493),
.A2(n_473),
.B1(n_481),
.B2(n_491),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_530),
.A2(n_493),
.B1(n_513),
.B2(n_511),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_472),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_494),
.B(n_468),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_522),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_499),
.A2(n_456),
.B1(n_434),
.B2(n_472),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_537),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_497),
.B(n_491),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_536),
.B(n_497),
.Y(n_545)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_498),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_520),
.A2(n_506),
.B(n_492),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_542),
.Y(n_554)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_523),
.A2(n_508),
.B1(n_507),
.B2(n_460),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_545),
.B(n_546),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_501),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_549),
.C(n_552),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_526),
.B(n_501),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_515),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_500),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_521),
.C(n_533),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_541),
.A2(n_525),
.B1(n_547),
.B2(n_551),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_556),
.A2(n_561),
.B1(n_441),
.B2(n_503),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_544),
.A2(n_516),
.B(n_500),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_557),
.A2(n_558),
.B(n_559),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_541),
.A2(n_534),
.B(n_459),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_546),
.A2(n_530),
.B(n_517),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_550),
.A2(n_532),
.B(n_520),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_560),
.B(n_562),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_538),
.A2(n_507),
.B1(n_532),
.B2(n_531),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_509),
.C(n_450),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_565),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_543),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_433),
.C(n_445),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_566),
.B(n_543),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_562),
.B(n_527),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_568),
.B(n_572),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_554),
.A2(n_555),
.B(n_558),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_574),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_560),
.B(n_495),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_555),
.B(n_554),
.C(n_567),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_565),
.B(n_514),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_557),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_576),
.B(n_563),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_577),
.B(n_559),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_567),
.A2(n_512),
.B1(n_467),
.B2(n_478),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_556),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_579),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_580),
.B(n_581),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_574),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_585),
.C(n_586),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_570),
.A2(n_563),
.B(n_561),
.Y(n_585)
);

A2O1A1Ixp33_ASAP7_75t_L g587 ( 
.A1(n_579),
.A2(n_586),
.B(n_583),
.C(n_571),
.Y(n_587)
);

OAI21x1_ASAP7_75t_SL g595 ( 
.A1(n_587),
.A2(n_591),
.B(n_577),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_584),
.A2(n_573),
.B(n_571),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_588),
.B(n_578),
.Y(n_594)
);

INVx11_ASAP7_75t_L g591 ( 
.A(n_583),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_589),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_593),
.B(n_595),
.C(n_590),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_594),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_596),
.A2(n_591),
.B1(n_592),
.B2(n_587),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_597),
.B(n_564),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_566),
.C(n_549),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_545),
.B(n_548),
.Y(n_601)
);


endmodule