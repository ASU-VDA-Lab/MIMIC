module fake_jpeg_24262_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_26),
.B1(n_33),
.B2(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_16),
.B1(n_32),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_52),
.B1(n_32),
.B2(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_49),
.B(n_15),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_31),
.A3(n_19),
.B1(n_23),
.B2(n_37),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_16),
.B1(n_32),
.B2(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_38),
.B1(n_28),
.B2(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_33),
.B1(n_17),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_61),
.B1(n_19),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_27),
.B1(n_21),
.B2(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_78),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_21),
.B(n_29),
.C(n_22),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_80),
.B1(n_87),
.B2(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_70),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_0),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_52),
.B1(n_6),
.B2(n_8),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_81),
.B1(n_95),
.B2(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_96),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_11),
.B1(n_5),
.B2(n_9),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_4),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_101),
.Y(n_113)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_100),
.B1(n_114),
.B2(n_123),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_86),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_107),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_56),
.C(n_66),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_126),
.C(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_69),
.B1(n_14),
.B2(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_9),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_9),
.B1(n_11),
.B2(n_87),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_124),
.B1(n_126),
.B2(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_74),
.B(n_11),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

FAx1_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_93),
.CI(n_97),
.CON(n_123),
.SN(n_123)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_76),
.B1(n_88),
.B2(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_70),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_88),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_143),
.B1(n_137),
.B2(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_91),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_141),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_104),
.A3(n_118),
.B1(n_117),
.B2(n_111),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_147),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_105),
.B1(n_123),
.B2(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_102),
.C(n_111),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_152),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_160),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_155),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_171),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_134),
.B1(n_152),
.B2(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_169),
.B1(n_149),
.B2(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_119),
.B(n_122),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_154),
.B(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_109),
.B1(n_128),
.B2(n_119),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_169),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_144),
.C(n_147),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_165),
.C(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_172),
.CI(n_159),
.CON(n_190),
.SN(n_190)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_187),
.B1(n_188),
.B2(n_181),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_171),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_198),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_194),
.C(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_200),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_165),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_162),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_178),
.B(n_156),
.C(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_190),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_177),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_183),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_179),
.B(n_175),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_184),
.C(n_181),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_216),
.C(n_218),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_209),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_179),
.C(n_184),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_203),
.B(n_211),
.C(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_198),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_203),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_187),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_225),
.B(n_202),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_219),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_SL g229 ( 
.A(n_226),
.B(n_222),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_196),
.C(n_166),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.C(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_230),
.B(n_149),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_210),
.Y(n_232)
);


endmodule