module fake_netlist_6_1602_n_2743 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_788, n_325, n_767, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2743);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_788;
input n_325;
input n_767;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2743;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_822;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_1663;
wire n_2009;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_1165;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2319;
wire n_2519;
wire n_825;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_890;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_1992;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1397;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_876;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_875;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_735),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_674),
.Y(n_800)
);

CKINVDCx16_ASAP7_75t_R g801 ( 
.A(n_207),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_143),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_515),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_666),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_737),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_441),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_476),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_772),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_312),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_777),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_545),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_573),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_798),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_254),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_388),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_353),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_613),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_259),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_671),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_628),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_559),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_716),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_576),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_371),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_190),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_728),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_769),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_763),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_260),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_327),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_128),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_322),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_364),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_62),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_246),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_533),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_472),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_236),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_582),
.Y(n_839)
);

CKINVDCx14_ASAP7_75t_R g840 ( 
.A(n_449),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_445),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_192),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_597),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_542),
.Y(n_844)
);

BUFx10_ASAP7_75t_L g845 ( 
.A(n_692),
.Y(n_845)
);

BUFx10_ASAP7_75t_L g846 ( 
.A(n_767),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_169),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_446),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_619),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_755),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_668),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_263),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_107),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_722),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_271),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_424),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_746),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_739),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_742),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_781),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_677),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_709),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_218),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_426),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_531),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_733),
.Y(n_866)
);

INVxp33_ASAP7_75t_L g867 ( 
.A(n_688),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_721),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_165),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_506),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_726),
.Y(n_871)
);

CKINVDCx16_ASAP7_75t_R g872 ( 
.A(n_719),
.Y(n_872)
);

CKINVDCx16_ASAP7_75t_R g873 ( 
.A(n_637),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_284),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_681),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_88),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_240),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_35),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_481),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_254),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_395),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_105),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_459),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_147),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_797),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_691),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_320),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_715),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_490),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_698),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_562),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_675),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_252),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_756),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_603),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_138),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_717),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_712),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_31),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_26),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_247),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_779),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_219),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_790),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_239),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_232),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_90),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_551),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_565),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_774),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_724),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_121),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_363),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_795),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_759),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_743),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_235),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_444),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_762),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_249),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_684),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_648),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_703),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_540),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_157),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_114),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_251),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_303),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_778),
.Y(n_929)
);

BUFx10_ASAP7_75t_L g930 ( 
.A(n_694),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_161),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_734),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_249),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_569),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_687),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_682),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_784),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_268),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_594),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_757),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_760),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_794),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_157),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_793),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_650),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_376),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_685),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_705),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_467),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_493),
.Y(n_950)
);

CKINVDCx14_ASAP7_75t_R g951 ( 
.A(n_745),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_664),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_730),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_758),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_738),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_318),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_342),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_427),
.Y(n_958)
);

CKINVDCx16_ASAP7_75t_R g959 ( 
.A(n_9),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_696),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_665),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_773),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_348),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_663),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_783),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_732),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_339),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_221),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_255),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_486),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_100),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_747),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_706),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_189),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_690),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_699),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_62),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_34),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_780),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_516),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_770),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_18),
.Y(n_983)
);

BUFx5_ASAP7_75t_L g984 ( 
.A(n_302),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_186),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_212),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_639),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_65),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_544),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_398),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_765),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_736),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_494),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_141),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_792),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_649),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_776),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_142),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_557),
.Y(n_999)
);

BUFx8_ASAP7_75t_SL g1000 ( 
.A(n_282),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_340),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_475),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_464),
.Y(n_1003)
);

BUFx2_ASAP7_75t_SL g1004 ( 
.A(n_714),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_748),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_321),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_121),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_530),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_561),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_788),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_325),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_676),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_127),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_528),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_283),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_617),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_695),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_711),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_713),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_286),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_586),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_686),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_262),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_270),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_15),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_630),
.Y(n_1026)
);

BUFx8_ASAP7_75t_SL g1027 ( 
.A(n_49),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_318),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_356),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_701),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_702),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_622),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_376),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_114),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_741),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_680),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_631),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_725),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_25),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_541),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_727),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_501),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_754),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_624),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_115),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_113),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_429),
.Y(n_1047)
);

CKINVDCx14_ASAP7_75t_R g1048 ( 
.A(n_279),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_2),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_77),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_334),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_704),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_76),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_195),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_6),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_729),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_723),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_697),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_731),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_679),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_498),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_445),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_478),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_220),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_782),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_775),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_752),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_708),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_766),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_277),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_220),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_791),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_749),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_305),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_787),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_645),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_477),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_421),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_678),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_323),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_700),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_710),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_764),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_233),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_88),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_471),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_786),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_63),
.Y(n_1088)
);

BUFx2_ASAP7_75t_SL g1089 ( 
.A(n_331),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_744),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_170),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_422),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_151),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_720),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_750),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_222),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_564),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_347),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_672),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_585),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_217),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_740),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_176),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_604),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_442),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_618),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_707),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_127),
.Y(n_1108)
);

BUFx10_ASAP7_75t_L g1109 ( 
.A(n_761),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_771),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_316),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_479),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_11),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_753),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_409),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_693),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_454),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_768),
.Y(n_1118)
);

CKINVDCx16_ASAP7_75t_R g1119 ( 
.A(n_547),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_91),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_718),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_656),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_290),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_612),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_175),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_689),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_621),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_789),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_683),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_751),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_591),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_626),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_785),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_563),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_497),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_245),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_215),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_83),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_802),
.B(n_0),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_984),
.Y(n_1140)
);

BUFx8_ASAP7_75t_L g1141 ( 
.A(n_812),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_857),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_913),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_840),
.B(n_0),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_857),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_806),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_806),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_815),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1048),
.B(n_1),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_949),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_845),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_984),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_826),
.B(n_1),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_835),
.B(n_970),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_950),
.B(n_2),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_894),
.B(n_3),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_916),
.B(n_3),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_913),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_801),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_993),
.B(n_4),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_949),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_996),
.B(n_4),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_984),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_857),
.B(n_489),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_859),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_984),
.Y(n_1166)
);

BUFx8_ASAP7_75t_L g1167 ( 
.A(n_984),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_913),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_867),
.B(n_6),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_924),
.B(n_7),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_955),
.B(n_7),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_984),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_864),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1154),
.B(n_817),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1169),
.A2(n_951),
.B1(n_823),
.B2(n_873),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1143),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1144),
.B(n_872),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1154),
.B(n_960),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1143),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1159),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1145),
.B(n_1082),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1158),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1158),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1162),
.A2(n_834),
.B1(n_918),
.B2(n_841),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1151),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1148),
.B(n_959),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1168),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_SL g1188 ( 
.A(n_1153),
.Y(n_1188)
);

OAI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1149),
.A2(n_833),
.B1(n_977),
.B2(n_946),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1155),
.A2(n_887),
.B1(n_1089),
.B2(n_825),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1170),
.A2(n_1119),
.B1(n_1068),
.B2(n_822),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1171),
.A2(n_843),
.B1(n_861),
.B2(n_799),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1173),
.B(n_926),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1146),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1168),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1139),
.A2(n_831),
.B1(n_838),
.B2(n_832),
.Y(n_1196)
);

AO22x2_ASAP7_75t_L g1197 ( 
.A1(n_1139),
.A2(n_842),
.B1(n_855),
.B2(n_848),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1147),
.A2(n_945),
.B1(n_961),
.B2(n_886),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1140),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1145),
.B(n_1165),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1165),
.B(n_1112),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1156),
.A2(n_863),
.B1(n_878),
.B2(n_869),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1152),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1157),
.A2(n_1080),
.B1(n_905),
.B2(n_809),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_SL g1205 ( 
.A(n_1164),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1163),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1177),
.A2(n_1160),
.B(n_1166),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1175),
.B(n_1150),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1186),
.B(n_1161),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1199),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1185),
.B(n_1141),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1192),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1178),
.B(n_824),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1193),
.B(n_1142),
.Y(n_1214)
);

XNOR2x2_ASAP7_75t_L g1215 ( 
.A(n_1191),
.B(n_876),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1203),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1174),
.B(n_1167),
.Y(n_1217)
);

AND2x6_ASAP7_75t_L g1218 ( 
.A(n_1206),
.B(n_859),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1201),
.B(n_1166),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1200),
.B(n_1172),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1176),
.Y(n_1221)
);

XOR2x2_ASAP7_75t_L g1222 ( 
.A(n_1184),
.B(n_1023),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1181),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1179),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1182),
.Y(n_1225)
);

INVxp33_ASAP7_75t_SL g1226 ( 
.A(n_1198),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1187),
.B(n_1118),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1195),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1190),
.B(n_1025),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_1189),
.B(n_978),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1190),
.B(n_1039),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1196),
.B(n_1070),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1196),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1204),
.B(n_845),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1197),
.B(n_1103),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1194),
.B(n_1035),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1188),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1197),
.Y(n_1239)
);

INVxp33_ASAP7_75t_L g1240 ( 
.A(n_1202),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1202),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1205),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1199),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1199),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1177),
.B(n_800),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1199),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_1192),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1199),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1199),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1199),
.Y(n_1250)
);

INVxp33_ASAP7_75t_L g1251 ( 
.A(n_1180),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1199),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1199),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1213),
.B(n_998),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1224),
.B(n_804),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1227),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1245),
.B(n_808),
.Y(n_1257)
);

AND2x4_ASAP7_75t_SL g1258 ( 
.A(n_1238),
.B(n_964),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1248),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1220),
.A2(n_821),
.B(n_811),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1210),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1207),
.B(n_813),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1251),
.B(n_1096),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1253),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1228),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1228),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1221),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1242),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1240),
.B(n_1212),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1239),
.B(n_807),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1214),
.B(n_1098),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1209),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1216),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1241),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1223),
.B(n_1219),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1243),
.B(n_827),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1244),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1246),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1234),
.B(n_849),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1249),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1250),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1252),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1233),
.B(n_814),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1236),
.B(n_816),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1211),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1229),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1230),
.B(n_818),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1231),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1232),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1217),
.B(n_850),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1215),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1218),
.Y(n_1293)
);

AND2x2_ASAP7_75t_SL g1294 ( 
.A(n_1208),
.B(n_978),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1237),
.B(n_854),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1235),
.B(n_868),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1218),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1218),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1222),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1218),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1247),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1226),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1248),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1248),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1227),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_1224),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1253),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1224),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1224),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1245),
.B(n_871),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1213),
.B(n_829),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1213),
.B(n_830),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1227),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1239),
.B(n_1004),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1227),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1248),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1248),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1213),
.B(n_837),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1224),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1213),
.B(n_847),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1245),
.A2(n_973),
.B1(n_1081),
.B2(n_1059),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1248),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1245),
.B(n_1100),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1248),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1253),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1207),
.A2(n_897),
.B(n_875),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1213),
.B(n_852),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1248),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1248),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1253),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1224),
.B(n_909),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1253),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1227),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1253),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1245),
.B(n_910),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1224),
.B(n_914),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1213),
.B(n_853),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1245),
.B(n_919),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1245),
.B(n_929),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1248),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1213),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1248),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1248),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1251),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1245),
.B(n_934),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1213),
.B(n_856),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1251),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1213),
.B(n_874),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1245),
.B(n_941),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1227),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1253),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1245),
.B(n_942),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1245),
.B(n_1126),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1224),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1253),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1245),
.B(n_947),
.Y(n_1356)
);

NAND2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1306),
.B(n_858),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1344),
.B(n_1136),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1323),
.B(n_954),
.Y(n_1359)
);

AND2x2_ASAP7_75t_SL g1360 ( 
.A(n_1353),
.B(n_978),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1306),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1341),
.B(n_1128),
.Y(n_1362)
);

NAND2x1_ASAP7_75t_SL g1363 ( 
.A(n_1321),
.B(n_880),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1315),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1256),
.B(n_877),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1259),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1275),
.B(n_962),
.Y(n_1367)
);

BUFx4f_ASAP7_75t_L g1368 ( 
.A(n_1289),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1265),
.B(n_899),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1285),
.B(n_1000),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1347),
.B(n_1138),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1333),
.B(n_900),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1268),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1350),
.B(n_920),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1259),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1343),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1272),
.B(n_928),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1343),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1305),
.B(n_879),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1308),
.B(n_933),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1303),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1257),
.B(n_975),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1319),
.B(n_1009),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1309),
.B(n_943),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1304),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1354),
.B(n_958),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1289),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1294),
.B(n_1027),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1313),
.B(n_881),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1316),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1266),
.B(n_967),
.Y(n_1391)
);

NOR2xp67_ASAP7_75t_L g1392 ( 
.A(n_1302),
.B(n_803),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1279),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1272),
.Y(n_1394)
);

AND2x4_ASAP7_75t_SL g1395 ( 
.A(n_1319),
.B(n_846),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1269),
.B(n_1060),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1264),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1317),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1310),
.B(n_976),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1279),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1271),
.B(n_1090),
.Y(n_1401)
);

INVx5_ASAP7_75t_L g1402 ( 
.A(n_1314),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1290),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1263),
.Y(n_1404)
);

AND2x6_ASAP7_75t_L g1405 ( 
.A(n_1292),
.B(n_980),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1258),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1335),
.B(n_982),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1338),
.B(n_1339),
.Y(n_1408)
);

AND2x2_ASAP7_75t_SL g1409 ( 
.A(n_1301),
.B(n_1254),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1311),
.B(n_882),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1322),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1255),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1299),
.B(n_1312),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1307),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1345),
.B(n_1349),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1255),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1325),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1270),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1331),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1324),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1331),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1314),
.B(n_969),
.Y(n_1422)
);

AND2x2_ASAP7_75t_SL g1423 ( 
.A(n_1352),
.B(n_1024),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1318),
.B(n_1320),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1328),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1356),
.B(n_989),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1274),
.B(n_983),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1329),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1340),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1330),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1326),
.B(n_997),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1267),
.Y(n_1432)
);

BUFx4f_ASAP7_75t_L g1433 ( 
.A(n_1283),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1332),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1327),
.B(n_883),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1273),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1337),
.B(n_893),
.Y(n_1437)
);

BUFx5_ASAP7_75t_L g1438 ( 
.A(n_1342),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1288),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1346),
.B(n_896),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1334),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1348),
.B(n_901),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1336),
.B(n_985),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1284),
.B(n_903),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1336),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1262),
.B(n_1016),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1351),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1261),
.B(n_994),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1281),
.B(n_1003),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1298),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1277),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_SL g1452 ( 
.A(n_1291),
.B(n_846),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1278),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1280),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1355),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1298),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1282),
.B(n_1015),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1286),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1287),
.B(n_1020),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1296),
.Y(n_1460)
);

BUFx4f_ASAP7_75t_L g1461 ( 
.A(n_1293),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1276),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1295),
.B(n_1018),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1297),
.B(n_1022),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_SL g1465 ( 
.A(n_1300),
.B(n_930),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1260),
.B(n_859),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1256),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1259),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1323),
.B(n_1041),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1323),
.B(n_1044),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1341),
.B(n_906),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1323),
.B(n_1052),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1259),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1323),
.B(n_1056),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1259),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1259),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1259),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1344),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1259),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1323),
.B(n_1057),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1341),
.B(n_907),
.Y(n_1481)
);

BUFx8_ASAP7_75t_SL g1482 ( 
.A(n_1301),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1315),
.B(n_1053),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1326),
.A2(n_1076),
.B(n_1073),
.Y(n_1484)
);

NOR2x1_ASAP7_75t_SL g1485 ( 
.A(n_1275),
.B(n_1083),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1323),
.B(n_1095),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1323),
.B(n_1102),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1306),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1259),
.Y(n_1489)
);

NAND2x1_ASAP7_75t_L g1490 ( 
.A(n_1259),
.B(n_1164),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1315),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1306),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1259),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1306),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1272),
.B(n_1055),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1341),
.B(n_912),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1306),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1323),
.B(n_1107),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1341),
.B(n_925),
.Y(n_1499)
);

NAND2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1306),
.B(n_1110),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1259),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1259),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1344),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1315),
.B(n_1071),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1341),
.B(n_927),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1344),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1272),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1323),
.B(n_1116),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1506),
.Y(n_1509)
);

BUFx8_ASAP7_75t_L g1510 ( 
.A(n_1478),
.Y(n_1510)
);

BUFx12f_ASAP7_75t_L g1511 ( 
.A(n_1394),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_1507),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1503),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1376),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1387),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1378),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1387),
.B(n_1024),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1482),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1368),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1373),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1424),
.B(n_931),
.Y(n_1521)
);

INVxp33_ASAP7_75t_L g1522 ( 
.A(n_1358),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1364),
.Y(n_1523)
);

INVx5_ASAP7_75t_L g1524 ( 
.A(n_1377),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1491),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1359),
.A2(n_1132),
.B1(n_1121),
.B2(n_1164),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1403),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1406),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1439),
.Y(n_1529)
);

NAND2x1p5_ASAP7_75t_L g1530 ( 
.A(n_1361),
.B(n_1024),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1418),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1402),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1456),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1473),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1413),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1404),
.Y(n_1536)
);

INVx5_ASAP7_75t_L g1537 ( 
.A(n_1495),
.Y(n_1537)
);

NOR2xp67_ASAP7_75t_SL g1538 ( 
.A(n_1488),
.B(n_1124),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1408),
.B(n_805),
.Y(n_1539)
);

BUFx2_ASAP7_75t_SL g1540 ( 
.A(n_1416),
.Y(n_1540)
);

BUFx5_ASAP7_75t_L g1541 ( 
.A(n_1366),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1396),
.A2(n_1129),
.B1(n_1130),
.B2(n_1127),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1477),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1412),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1402),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1447),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1371),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1379),
.B(n_938),
.Y(n_1549)
);

CKINVDCx11_ASAP7_75t_R g1550 ( 
.A(n_1427),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1483),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1419),
.B(n_1086),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1467),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1493),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1445),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1412),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1415),
.B(n_810),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1421),
.Y(n_1558)
);

INVx5_ASAP7_75t_SL g1559 ( 
.A(n_1422),
.Y(n_1559)
);

BUFx4f_ASAP7_75t_SL g1560 ( 
.A(n_1409),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_SL g1561 ( 
.A(n_1504),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1380),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1492),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1501),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1401),
.B(n_956),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1494),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1393),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1469),
.B(n_819),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1497),
.Y(n_1569)
);

NOR2xp67_ASAP7_75t_L g1570 ( 
.A(n_1460),
.B(n_1432),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1362),
.Y(n_1571)
);

BUFx2_ASAP7_75t_SL g1572 ( 
.A(n_1393),
.Y(n_1572)
);

INVx6_ASAP7_75t_L g1573 ( 
.A(n_1384),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1386),
.Y(n_1574)
);

BUFx4_ASAP7_75t_SL g1575 ( 
.A(n_1422),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1433),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1372),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1395),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1365),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1374),
.Y(n_1580)
);

INVx8_ASAP7_75t_L g1581 ( 
.A(n_1449),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1363),
.Y(n_1582)
);

BUFx2_ASAP7_75t_SL g1583 ( 
.A(n_1400),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1450),
.Y(n_1584)
);

CKINVDCx11_ASAP7_75t_R g1585 ( 
.A(n_1443),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1502),
.Y(n_1586)
);

INVx5_ASAP7_75t_L g1587 ( 
.A(n_1405),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1470),
.B(n_820),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_SL g1589 ( 
.A(n_1405),
.Y(n_1589)
);

INVx5_ASAP7_75t_L g1590 ( 
.A(n_1405),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1410),
.B(n_957),
.Y(n_1591)
);

BUFx4_ASAP7_75t_SL g1592 ( 
.A(n_1451),
.Y(n_1592)
);

INVx5_ASAP7_75t_L g1593 ( 
.A(n_1455),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1448),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1455),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1472),
.A2(n_965),
.B1(n_979),
.B2(n_895),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1360),
.B(n_930),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1474),
.B(n_828),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1457),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1459),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1458),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1375),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1468),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1475),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1479),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1391),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1461),
.Y(n_1607)
);

INVx8_ASAP7_75t_L g1608 ( 
.A(n_1369),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1436),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1489),
.Y(n_1610)
);

BUFx2_ASAP7_75t_SL g1611 ( 
.A(n_1438),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1389),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1471),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1454),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_SL g1615 ( 
.A(n_1381),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1481),
.Y(n_1616)
);

BUFx12f_ASAP7_75t_L g1617 ( 
.A(n_1357),
.Y(n_1617)
);

BUFx12f_ASAP7_75t_L g1618 ( 
.A(n_1383),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1453),
.B(n_1385),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1500),
.Y(n_1620)
);

BUFx5_ASAP7_75t_L g1621 ( 
.A(n_1390),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1398),
.B(n_1091),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1496),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1397),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1480),
.A2(n_971),
.B1(n_974),
.B2(n_963),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1519),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1519),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1565),
.A2(n_1388),
.B1(n_1452),
.B2(n_1560),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1547),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1548),
.A2(n_1486),
.B1(n_1498),
.B2(n_1487),
.Y(n_1630)
);

INVx6_ASAP7_75t_L g1631 ( 
.A(n_1510),
.Y(n_1631)
);

INVx6_ASAP7_75t_L g1632 ( 
.A(n_1511),
.Y(n_1632)
);

BUFx10_ASAP7_75t_L g1633 ( 
.A(n_1615),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1619),
.A2(n_1508),
.B1(n_1431),
.B2(n_1367),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1553),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1525),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1571),
.A2(n_1423),
.B1(n_1435),
.B2(n_1444),
.Y(n_1638)
);

BUFx8_ASAP7_75t_SL g1639 ( 
.A(n_1518),
.Y(n_1639)
);

INVx6_ASAP7_75t_L g1640 ( 
.A(n_1593),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1625),
.A2(n_1597),
.B1(n_1616),
.B2(n_1613),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1617),
.A2(n_1465),
.B1(n_1370),
.B2(n_1442),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1623),
.A2(n_1437),
.B1(n_1440),
.B2(n_1499),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1539),
.B(n_1557),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

INVx6_ASAP7_75t_L g1646 ( 
.A(n_1520),
.Y(n_1646)
);

CKINVDCx11_ASAP7_75t_R g1647 ( 
.A(n_1532),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1579),
.A2(n_1392),
.B1(n_1505),
.B2(n_1462),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1610),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1612),
.A2(n_1420),
.B1(n_1425),
.B2(n_1411),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1602),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1604),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1568),
.B(n_1428),
.Y(n_1653)
);

CKINVDCx11_ASAP7_75t_R g1654 ( 
.A(n_1546),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1605),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1513),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1509),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1536),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1582),
.A2(n_1484),
.B1(n_1429),
.B2(n_1417),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1535),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1544),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1529),
.Y(n_1662)
);

INVx6_ASAP7_75t_L g1663 ( 
.A(n_1512),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1578),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1614),
.A2(n_1446),
.B1(n_1399),
.B2(n_1407),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1618),
.A2(n_1485),
.B1(n_1382),
.B2(n_1426),
.Y(n_1666)
);

CKINVDCx11_ASAP7_75t_R g1667 ( 
.A(n_1550),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1588),
.B(n_1438),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1527),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1591),
.A2(n_1414),
.B1(n_1434),
.B2(n_1430),
.Y(n_1670)
);

BUFx8_ASAP7_75t_L g1671 ( 
.A(n_1589),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1521),
.A2(n_1441),
.B1(n_1438),
.B2(n_1463),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1598),
.B(n_1464),
.Y(n_1673)
);

CKINVDCx11_ASAP7_75t_R g1674 ( 
.A(n_1585),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1545),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1576),
.Y(n_1676)
);

BUFx12f_ASAP7_75t_L g1677 ( 
.A(n_1528),
.Y(n_1677)
);

INVx4_ASAP7_75t_L g1678 ( 
.A(n_1545),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1522),
.A2(n_1133),
.B1(n_1134),
.B2(n_1131),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1514),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1595),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1516),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1533),
.Y(n_1683)
);

BUFx12f_ASAP7_75t_SL g1684 ( 
.A(n_1517),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1554),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1564),
.Y(n_1686)
);

OAI21xp33_ASAP7_75t_L g1687 ( 
.A1(n_1542),
.A2(n_988),
.B(n_986),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1523),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1580),
.A2(n_1622),
.B1(n_1577),
.B2(n_1552),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1570),
.A2(n_1490),
.B1(n_1466),
.B2(n_1032),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1534),
.A2(n_1109),
.B1(n_1066),
.B2(n_1069),
.Y(n_1691)
);

CKINVDCx11_ASAP7_75t_R g1692 ( 
.A(n_1531),
.Y(n_1692)
);

BUFx10_ASAP7_75t_L g1693 ( 
.A(n_1561),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1524),
.A2(n_1109),
.B1(n_1001),
.B2(n_1002),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1543),
.A2(n_1079),
.B1(n_981),
.B2(n_1115),
.Y(n_1695)
);

BUFx12f_ASAP7_75t_L g1696 ( 
.A(n_1524),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1586),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1624),
.A2(n_1137),
.B1(n_1092),
.B2(n_839),
.Y(n_1698)
);

BUFx12f_ASAP7_75t_L g1699 ( 
.A(n_1537),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1601),
.B(n_836),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1555),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1595),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1551),
.A2(n_1135),
.B1(n_851),
.B2(n_860),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1549),
.A2(n_862),
.B1(n_865),
.B2(n_844),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1594),
.A2(n_870),
.B1(n_885),
.B2(n_866),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1599),
.A2(n_888),
.B1(n_890),
.B2(n_889),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1600),
.A2(n_891),
.B1(n_898),
.B2(n_892),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1611),
.A2(n_902),
.B1(n_908),
.B2(n_904),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1515),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1558),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1567),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1573),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1562),
.Y(n_1713)
);

CKINVDCx6p67_ASAP7_75t_R g1714 ( 
.A(n_1537),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1609),
.Y(n_1715)
);

CKINVDCx11_ASAP7_75t_R g1716 ( 
.A(n_1581),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1608),
.A2(n_911),
.B1(n_921),
.B2(n_915),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1592),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1596),
.A2(n_923),
.B1(n_932),
.B2(n_922),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1569),
.B(n_935),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1559),
.A2(n_1006),
.B1(n_1007),
.B2(n_990),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1621),
.Y(n_1722)
);

BUFx4_ASAP7_75t_SL g1723 ( 
.A(n_1574),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1621),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1606),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1621),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1541),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1563),
.A2(n_937),
.B1(n_939),
.B2(n_936),
.Y(n_1728)
);

OAI22x1_ASAP7_75t_SL g1729 ( 
.A1(n_1587),
.A2(n_1013),
.B1(n_1028),
.B2(n_1011),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1566),
.A2(n_944),
.B1(n_948),
.B2(n_940),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1606),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1541),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1530),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1556),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1620),
.A2(n_953),
.B1(n_966),
.B2(n_952),
.Y(n_1735)
);

CKINVDCx6p67_ASAP7_75t_R g1736 ( 
.A(n_1587),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1607),
.Y(n_1737)
);

BUFx8_ASAP7_75t_L g1738 ( 
.A(n_1575),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1590),
.A2(n_1572),
.B1(n_1583),
.B2(n_1540),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1590),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1584),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1526),
.A2(n_1033),
.B1(n_1034),
.B2(n_1029),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1538),
.B(n_972),
.Y(n_1743)
);

INVx4_ASAP7_75t_L g1744 ( 
.A(n_1519),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1565),
.A2(n_991),
.B1(n_992),
.B2(n_987),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1519),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1547),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1603),
.Y(n_1748)
);

CKINVDCx11_ASAP7_75t_R g1749 ( 
.A(n_1511),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1619),
.A2(n_999),
.B1(n_1005),
.B2(n_995),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1519),
.Y(n_1751)
);

BUFx12f_ASAP7_75t_L g1752 ( 
.A(n_1585),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1657),
.Y(n_1753)
);

BUFx12f_ASAP7_75t_L g1754 ( 
.A(n_1749),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1687),
.A2(n_1046),
.B1(n_1047),
.B2(n_1045),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1651),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1630),
.A2(n_1010),
.B(n_1008),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1638),
.A2(n_1050),
.B1(n_1051),
.B2(n_1049),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1644),
.A2(n_1063),
.B1(n_1064),
.B2(n_1054),
.Y(n_1759)
);

BUFx4f_ASAP7_75t_SL g1760 ( 
.A(n_1696),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1652),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1643),
.A2(n_1077),
.B1(n_1078),
.B2(n_1074),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1635),
.A2(n_1085),
.B1(n_1088),
.B2(n_1084),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1628),
.B(n_1012),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1642),
.A2(n_1101),
.B1(n_1105),
.B2(n_1093),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1648),
.A2(n_1653),
.B1(n_1660),
.B2(n_1656),
.Y(n_1766)
);

NAND2xp33_ASAP7_75t_SL g1767 ( 
.A(n_1676),
.B(n_1741),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1694),
.A2(n_1111),
.B1(n_1113),
.B2(n_1108),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1655),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_SL g1770 ( 
.A1(n_1663),
.A2(n_1120),
.B1(n_1125),
.B2(n_1117),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1661),
.Y(n_1771)
);

OAI222xp33_ASAP7_75t_L g1772 ( 
.A1(n_1650),
.A2(n_1742),
.B1(n_1666),
.B2(n_1636),
.C1(n_1641),
.C2(n_1673),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_SL g1773 ( 
.A1(n_1663),
.A2(n_917),
.B1(n_968),
.B2(n_884),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1658),
.B(n_1645),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1681),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1649),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1640),
.Y(n_1777)
);

BUFx12f_ASAP7_75t_L g1778 ( 
.A(n_1647),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1745),
.A2(n_1017),
.B1(n_1019),
.B2(n_1014),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1721),
.A2(n_1123),
.B1(n_1062),
.B2(n_1026),
.Y(n_1780)
);

BUFx8_ASAP7_75t_SL g1781 ( 
.A(n_1639),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1748),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1665),
.A2(n_1099),
.B1(n_1061),
.B2(n_1030),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1685),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1680),
.B(n_1021),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1629),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1672),
.A2(n_1122),
.B1(n_1072),
.B2(n_1036),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1682),
.B(n_1031),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1669),
.B(n_1037),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1640),
.Y(n_1790)
);

NAND2xp33_ASAP7_75t_R g1791 ( 
.A(n_1662),
.B(n_1038),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1711),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1699),
.A2(n_1042),
.B1(n_1043),
.B2(n_1040),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1686),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1704),
.A2(n_1668),
.B1(n_1691),
.B2(n_1659),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1646),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1747),
.B(n_1058),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1631),
.A2(n_1067),
.B1(n_1075),
.B2(n_1065),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1646),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1627),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1689),
.A2(n_1094),
.B1(n_1104),
.B2(n_1087),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1670),
.A2(n_1106),
.B1(n_1114),
.B2(n_1097),
.Y(n_1802)
);

OAI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1714),
.A2(n_9),
.B1(n_5),
.B2(n_8),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1750),
.A2(n_10),
.B1(n_5),
.B2(n_8),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1631),
.A2(n_18),
.B1(n_26),
.B2(n_10),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1697),
.Y(n_1806)
);

OAI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1710),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1667),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1701),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1723),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1738),
.A2(n_23),
.B1(n_32),
.B2(n_14),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1698),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1812)
);

BUFx4f_ASAP7_75t_SL g1813 ( 
.A(n_1677),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1739),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_1814)
);

INVx4_ASAP7_75t_R g1815 ( 
.A(n_1626),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1679),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1713),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1705),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1709),
.Y(n_1819)
);

INVx5_ASAP7_75t_SL g1820 ( 
.A(n_1627),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1695),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1821)
);

OAI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1736),
.A2(n_1737),
.B1(n_1703),
.B2(n_1718),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1706),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1632),
.A2(n_35),
.B1(n_43),
.B2(n_27),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1674),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1708),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1707),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1722),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1728),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1730),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1724),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1726),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1727),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1735),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1709),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1700),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1732),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1740),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1734),
.B(n_491),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1715),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1688),
.Y(n_1841)
);

CKINVDCx8_ASAP7_75t_R g1842 ( 
.A(n_1681),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1816),
.A2(n_1743),
.B1(n_1684),
.B2(n_1632),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1780),
.A2(n_1733),
.B1(n_1692),
.B2(n_1752),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1765),
.A2(n_1717),
.B1(n_1720),
.B2(n_1725),
.C(n_1719),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1763),
.A2(n_1671),
.B1(n_1654),
.B2(n_1633),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1776),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1782),
.B(n_1731),
.Y(n_1848)
);

OA21x2_ASAP7_75t_L g1849 ( 
.A1(n_1828),
.A2(n_1690),
.B(n_1637),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1818),
.A2(n_1693),
.B1(n_1716),
.B2(n_1712),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1756),
.Y(n_1851)
);

OAI222xp33_ASAP7_75t_L g1852 ( 
.A1(n_1824),
.A2(n_1634),
.B1(n_1744),
.B2(n_1678),
.C1(n_1675),
.C2(n_1746),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1823),
.A2(n_1702),
.B1(n_1664),
.B2(n_1751),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_L g1854 ( 
.A(n_1834),
.B(n_1702),
.C(n_1741),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1836),
.A2(n_1729),
.B1(n_1683),
.B2(n_42),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1807),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.C(n_43),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1827),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1804),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1812),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1826),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1840),
.B(n_492),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1766),
.B(n_50),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1774),
.B(n_51),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1761),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1829),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1753),
.B(n_52),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1803),
.A2(n_55),
.B1(n_56),
.B2(n_54),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1757),
.B(n_53),
.C(n_54),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1830),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1806),
.B(n_57),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1814),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1821),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1822),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1768),
.A2(n_65),
.B1(n_61),
.B2(n_64),
.Y(n_1874)
);

OAI211xp5_ASAP7_75t_L g1875 ( 
.A1(n_1811),
.A2(n_1805),
.B(n_1838),
.C(n_1759),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1842),
.Y(n_1876)
);

AO22x1_ASAP7_75t_L g1877 ( 
.A1(n_1809),
.A2(n_1808),
.B1(n_1825),
.B2(n_1839),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1764),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1773),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1815),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1795),
.A2(n_1783),
.B1(n_1758),
.B2(n_1786),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1755),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1785),
.B(n_495),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1792),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1779),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1791),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1817),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1788),
.B(n_496),
.Y(n_1888)
);

NAND3xp33_ASAP7_75t_L g1889 ( 
.A(n_1770),
.B(n_75),
.C(n_78),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1772),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1801),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1762),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1797),
.A2(n_85),
.B1(n_82),
.B2(n_84),
.C(n_86),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1839),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1798),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1789),
.A2(n_91),
.B1(n_87),
.B2(n_89),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1767),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1771),
.B(n_92),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1793),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1802),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1769),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1784),
.B(n_96),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1841),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_SL g1904 ( 
.A1(n_1813),
.A2(n_1754),
.B1(n_1760),
.B2(n_1778),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1794),
.B(n_98),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1810),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1787),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1777),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1796),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1831),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1832),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1833),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1820),
.A2(n_116),
.B1(n_112),
.B2(n_115),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1837),
.B(n_499),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1790),
.A2(n_514),
.B(n_505),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1796),
.A2(n_118),
.B1(n_119),
.B2(n_117),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1799),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1819),
.A2(n_122),
.B1(n_119),
.B2(n_120),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_L g1919 ( 
.A(n_1868),
.B(n_1835),
.C(n_1799),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1847),
.B(n_1820),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1851),
.B(n_1775),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1890),
.A2(n_1800),
.B1(n_1775),
.B2(n_1781),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1864),
.B(n_1775),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1881),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1901),
.B(n_123),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1863),
.B(n_124),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1855),
.A2(n_128),
.B(n_126),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1862),
.B(n_125),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1898),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1902),
.B(n_125),
.Y(n_1930)
);

AOI211xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1867),
.A2(n_130),
.B(n_126),
.C(n_129),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1844),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1905),
.B(n_131),
.Y(n_1933)
);

NAND4xp25_ASAP7_75t_L g1934 ( 
.A(n_1886),
.B(n_134),
.C(n_132),
.D(n_133),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1876),
.B(n_132),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1875),
.B(n_133),
.C(n_134),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1873),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1870),
.B(n_135),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_L g1939 ( 
.A(n_1893),
.B(n_1889),
.C(n_1874),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1848),
.B(n_1861),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1914),
.B(n_136),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1866),
.B(n_137),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1896),
.B(n_139),
.Y(n_1943)
);

NAND3xp33_ASAP7_75t_L g1944 ( 
.A(n_1891),
.B(n_139),
.C(n_140),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1856),
.B(n_140),
.C(n_141),
.Y(n_1945)
);

AND4x1_ASAP7_75t_L g1946 ( 
.A(n_1846),
.B(n_144),
.C(n_142),
.D(n_143),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1883),
.B(n_144),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1888),
.B(n_145),
.Y(n_1948)
);

OAI221xp5_ASAP7_75t_SL g1949 ( 
.A1(n_1899),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1880),
.B(n_146),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1884),
.B(n_148),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1876),
.B(n_149),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1877),
.B(n_149),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1876),
.B(n_150),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1853),
.B(n_150),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1882),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_1956)
);

OA211x2_ASAP7_75t_L g1957 ( 
.A1(n_1897),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1910),
.B(n_155),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_L g1959 ( 
.A(n_1885),
.B(n_156),
.C(n_158),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1911),
.B(n_156),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1843),
.B(n_158),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1912),
.B(n_159),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1849),
.B(n_159),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1895),
.B(n_160),
.C(n_161),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1903),
.B(n_160),
.Y(n_1965)
);

OAI211xp5_ASAP7_75t_L g1966 ( 
.A1(n_1908),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1850),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1879),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1849),
.B(n_166),
.Y(n_1969)
);

OAI21xp33_ASAP7_75t_L g1970 ( 
.A1(n_1878),
.A2(n_167),
.B(n_168),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1916),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1894),
.B(n_171),
.Y(n_1972)
);

AND2x2_ASAP7_75t_SL g1973 ( 
.A(n_1871),
.B(n_172),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1918),
.B(n_172),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1906),
.B(n_173),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1892),
.B(n_173),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1854),
.B(n_500),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1900),
.B(n_174),
.Y(n_1978)
);

OA21x2_ASAP7_75t_L g1979 ( 
.A1(n_1857),
.A2(n_174),
.B(n_175),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1913),
.B(n_176),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1904),
.B(n_177),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1865),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1887),
.B(n_178),
.Y(n_1983)
);

NOR3xp33_ASAP7_75t_L g1984 ( 
.A(n_1845),
.B(n_179),
.C(n_180),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1860),
.B(n_180),
.Y(n_1985)
);

OAI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1907),
.A2(n_181),
.B(n_182),
.Y(n_1986)
);

OAI21xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1852),
.A2(n_183),
.B(n_182),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1869),
.B(n_181),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1858),
.B(n_183),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_R g1990 ( 
.A(n_1859),
.B(n_502),
.Y(n_1990)
);

NAND4xp25_ASAP7_75t_L g1991 ( 
.A(n_1872),
.B(n_186),
.C(n_184),
.D(n_185),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1909),
.B(n_184),
.Y(n_1992)
);

OAI21xp33_ASAP7_75t_L g1993 ( 
.A1(n_1917),
.A2(n_185),
.B(n_187),
.Y(n_1993)
);

OAI21xp5_ASAP7_75t_SL g1994 ( 
.A1(n_1915),
.A2(n_189),
.B(n_188),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1847),
.B(n_187),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1847),
.B(n_188),
.Y(n_1996)
);

OAI21xp33_ASAP7_75t_L g1997 ( 
.A1(n_1890),
.A2(n_190),
.B(n_191),
.Y(n_1997)
);

OA21x2_ASAP7_75t_L g1998 ( 
.A1(n_1868),
.A2(n_191),
.B(n_192),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_L g1999 ( 
.A(n_1868),
.B(n_193),
.C(n_194),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1847),
.B(n_193),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1868),
.B(n_194),
.C(n_195),
.Y(n_2001)
);

OAI221xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1886),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_2002)
);

OAI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1855),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_2003)
);

NOR2xp67_ASAP7_75t_L g2004 ( 
.A(n_1880),
.B(n_200),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1851),
.B(n_200),
.Y(n_2005)
);

OAI221xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1886),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1847),
.B(n_201),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1847),
.B(n_202),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1847),
.B(n_203),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1923),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1940),
.B(n_204),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_1984),
.B(n_205),
.C(n_206),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1929),
.B(n_205),
.Y(n_2013)
);

NAND4xp75_ASAP7_75t_L g2014 ( 
.A(n_1957),
.B(n_208),
.C(n_206),
.D(n_207),
.Y(n_2014)
);

AO21x2_ASAP7_75t_L g2015 ( 
.A1(n_1963),
.A2(n_208),
.B(n_209),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1952),
.B(n_209),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1920),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1936),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1921),
.B(n_210),
.Y(n_2019)
);

OA211x2_ASAP7_75t_L g2020 ( 
.A1(n_1919),
.A2(n_214),
.B(n_211),
.C(n_213),
.Y(n_2020)
);

NOR3xp33_ASAP7_75t_L g2021 ( 
.A(n_1939),
.B(n_213),
.C(n_214),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1954),
.B(n_215),
.Y(n_2022)
);

AO21x2_ASAP7_75t_L g2023 ( 
.A1(n_1969),
.A2(n_216),
.B(n_217),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1925),
.B(n_216),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_SL g2025 ( 
.A1(n_1973),
.A2(n_221),
.B1(n_218),
.B2(n_219),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1987),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1981),
.B(n_223),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1995),
.B(n_224),
.Y(n_2028)
);

NOR3xp33_ASAP7_75t_L g2029 ( 
.A(n_2002),
.B(n_225),
.C(n_226),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1996),
.B(n_225),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2005),
.B(n_1938),
.Y(n_2031)
);

NAND4xp75_ASAP7_75t_L g2032 ( 
.A(n_1998),
.B(n_228),
.C(n_226),
.D(n_227),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_L g2033 ( 
.A(n_2006),
.B(n_227),
.C(n_228),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1935),
.B(n_1950),
.Y(n_2034)
);

NOR3xp33_ASAP7_75t_L g2035 ( 
.A(n_1994),
.B(n_229),
.C(n_230),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2000),
.Y(n_2036)
);

NOR3xp33_ASAP7_75t_L g2037 ( 
.A(n_1999),
.B(n_229),
.C(n_230),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_1927),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.C(n_234),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1941),
.B(n_231),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_2009),
.B(n_234),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_2007),
.B(n_235),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1953),
.B(n_2008),
.Y(n_2042)
);

NOR3xp33_ASAP7_75t_L g2043 ( 
.A(n_2001),
.B(n_2003),
.C(n_1944),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1961),
.B(n_236),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_SL g2045 ( 
.A(n_1946),
.B(n_1931),
.C(n_1966),
.Y(n_2045)
);

NAND4xp75_ASAP7_75t_L g2046 ( 
.A(n_1998),
.B(n_239),
.C(n_237),
.D(n_238),
.Y(n_2046)
);

NAND4xp75_ASAP7_75t_L g2047 ( 
.A(n_1971),
.B(n_240),
.C(n_237),
.D(n_238),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1930),
.B(n_241),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_1956),
.B(n_241),
.C(n_242),
.Y(n_2049)
);

NOR2x1_ASAP7_75t_L g2050 ( 
.A(n_1933),
.B(n_242),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1926),
.B(n_243),
.Y(n_2051)
);

NAND3xp33_ASAP7_75t_L g2052 ( 
.A(n_1964),
.B(n_243),
.C(n_244),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1942),
.Y(n_2053)
);

NAND4xp75_ASAP7_75t_L g2054 ( 
.A(n_1968),
.B(n_246),
.C(n_244),
.D(n_245),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1947),
.B(n_247),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1948),
.B(n_248),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1997),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1928),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1979),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1943),
.B(n_250),
.Y(n_2060)
);

NAND3xp33_ASAP7_75t_L g2061 ( 
.A(n_1945),
.B(n_252),
.C(n_253),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1979),
.B(n_253),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1955),
.B(n_255),
.Y(n_2063)
);

AOI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_1949),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_1977),
.Y(n_2065)
);

NOR3xp33_ASAP7_75t_L g2066 ( 
.A(n_1937),
.B(n_256),
.C(n_257),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1983),
.Y(n_2067)
);

NOR2x1_ASAP7_75t_L g2068 ( 
.A(n_2004),
.B(n_258),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_1934),
.B(n_259),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_SL g2070 ( 
.A1(n_1990),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1991),
.A2(n_265),
.B1(n_261),
.B2(n_264),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1992),
.B(n_264),
.Y(n_2072)
);

AOI221x1_ASAP7_75t_L g2073 ( 
.A1(n_1993),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_1975),
.B(n_266),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1986),
.A2(n_270),
.B1(n_267),
.B2(n_269),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_R g2076 ( 
.A(n_1980),
.B(n_269),
.Y(n_2076)
);

BUFx2_ASAP7_75t_L g2077 ( 
.A(n_1972),
.Y(n_2077)
);

AO21x2_ASAP7_75t_L g2078 ( 
.A1(n_1976),
.A2(n_271),
.B(n_272),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1958),
.Y(n_2079)
);

BUFx12f_ASAP7_75t_L g2080 ( 
.A(n_1932),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1922),
.B(n_1951),
.Y(n_2081)
);

NOR3xp33_ASAP7_75t_L g2082 ( 
.A(n_1924),
.B(n_272),
.C(n_273),
.Y(n_2082)
);

AOI211x1_ASAP7_75t_L g2083 ( 
.A1(n_1967),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_L g2084 ( 
.A(n_1959),
.B(n_274),
.C(n_275),
.Y(n_2084)
);

AO21x2_ASAP7_75t_L g2085 ( 
.A1(n_1978),
.A2(n_276),
.B(n_277),
.Y(n_2085)
);

NOR3xp33_ASAP7_75t_L g2086 ( 
.A(n_1970),
.B(n_276),
.C(n_278),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_1974),
.Y(n_2087)
);

NAND3xp33_ASAP7_75t_L g2088 ( 
.A(n_1960),
.B(n_278),
.C(n_279),
.Y(n_2088)
);

NAND3xp33_ASAP7_75t_L g2089 ( 
.A(n_1962),
.B(n_1965),
.C(n_1985),
.Y(n_2089)
);

NAND3xp33_ASAP7_75t_L g2090 ( 
.A(n_1988),
.B(n_280),
.C(n_281),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1989),
.B(n_280),
.Y(n_2091)
);

OAI211xp5_ASAP7_75t_L g2092 ( 
.A1(n_1982),
.A2(n_289),
.B(n_297),
.C(n_281),
.Y(n_2092)
);

NAND3xp33_ASAP7_75t_L g2093 ( 
.A(n_1984),
.B(n_282),
.C(n_283),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_L g2094 ( 
.A(n_1919),
.B(n_284),
.Y(n_2094)
);

XNOR2x2_ASAP7_75t_L g2095 ( 
.A(n_1934),
.B(n_286),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1923),
.Y(n_2096)
);

NAND4xp75_ASAP7_75t_L g2097 ( 
.A(n_1957),
.B(n_288),
.C(n_285),
.D(n_287),
.Y(n_2097)
);

NAND3xp33_ASAP7_75t_L g2098 ( 
.A(n_1984),
.B(n_285),
.C(n_287),
.Y(n_2098)
);

NOR3xp33_ASAP7_75t_L g2099 ( 
.A(n_1984),
.B(n_288),
.C(n_289),
.Y(n_2099)
);

NOR3xp33_ASAP7_75t_L g2100 ( 
.A(n_1984),
.B(n_290),
.C(n_291),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1940),
.B(n_291),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_1929),
.B(n_292),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1940),
.B(n_292),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1923),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1921),
.Y(n_2105)
);

NAND4xp75_ASAP7_75t_L g2106 ( 
.A(n_1957),
.B(n_295),
.C(n_293),
.D(n_294),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2010),
.B(n_293),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2096),
.Y(n_2108)
);

XOR2x2_ASAP7_75t_L g2109 ( 
.A(n_2095),
.B(n_294),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_2017),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2104),
.B(n_295),
.Y(n_2111)
);

XOR2x2_ASAP7_75t_L g2112 ( 
.A(n_2034),
.B(n_296),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2105),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2036),
.Y(n_2114)
);

NAND4xp75_ASAP7_75t_SL g2115 ( 
.A(n_2069),
.B(n_298),
.C(n_296),
.D(n_297),
.Y(n_2115)
);

XOR2x2_ASAP7_75t_L g2116 ( 
.A(n_2045),
.B(n_298),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2059),
.Y(n_2117)
);

NAND4xp75_ASAP7_75t_SL g2118 ( 
.A(n_2081),
.B(n_301),
.C(n_299),
.D(n_300),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2042),
.B(n_300),
.Y(n_2119)
);

XNOR2xp5_ASAP7_75t_L g2120 ( 
.A(n_2016),
.B(n_301),
.Y(n_2120)
);

XOR2x2_ASAP7_75t_L g2121 ( 
.A(n_2068),
.B(n_302),
.Y(n_2121)
);

NAND4xp25_ASAP7_75t_L g2122 ( 
.A(n_2064),
.B(n_305),
.C(n_303),
.D(n_304),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2042),
.B(n_2077),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_2058),
.B(n_304),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2067),
.Y(n_2125)
);

NAND4xp75_ASAP7_75t_L g2126 ( 
.A(n_2073),
.B(n_308),
.C(n_306),
.D(n_307),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2053),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2087),
.B(n_307),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2079),
.B(n_308),
.Y(n_2129)
);

INVxp33_ASAP7_75t_L g2130 ( 
.A(n_2076),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_2015),
.Y(n_2131)
);

BUFx2_ASAP7_75t_L g2132 ( 
.A(n_2023),
.Y(n_2132)
);

OAI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2026),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2133)
);

NAND3xp33_ASAP7_75t_SL g2134 ( 
.A(n_2021),
.B(n_311),
.C(n_310),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2102),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2031),
.B(n_309),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2062),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2019),
.B(n_312),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2028),
.Y(n_2139)
);

NOR3xp33_ASAP7_75t_L g2140 ( 
.A(n_2012),
.B(n_313),
.C(n_314),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2030),
.B(n_313),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2040),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2011),
.B(n_314),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2013),
.Y(n_2144)
);

NOR4xp25_ASAP7_75t_L g2145 ( 
.A(n_2038),
.B(n_317),
.C(n_315),
.D(n_316),
.Y(n_2145)
);

NOR2x1_ASAP7_75t_L g2146 ( 
.A(n_2032),
.B(n_315),
.Y(n_2146)
);

XOR2xp5_ASAP7_75t_L g2147 ( 
.A(n_2089),
.B(n_503),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_2041),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_2065),
.B(n_317),
.Y(n_2149)
);

INVx2_ASAP7_75t_SL g2150 ( 
.A(n_2048),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2101),
.B(n_319),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2078),
.Y(n_2152)
);

NOR2x1_ASAP7_75t_R g2153 ( 
.A(n_2080),
.B(n_319),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2085),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_2051),
.Y(n_2155)
);

XOR2x2_ASAP7_75t_L g2156 ( 
.A(n_2022),
.B(n_320),
.Y(n_2156)
);

NAND4xp75_ASAP7_75t_L g2157 ( 
.A(n_2073),
.B(n_323),
.C(n_321),
.D(n_322),
.Y(n_2157)
);

NAND4xp75_ASAP7_75t_SL g2158 ( 
.A(n_2091),
.B(n_326),
.C(n_324),
.D(n_325),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2060),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2074),
.Y(n_2160)
);

AND2x2_ASAP7_75t_SL g2161 ( 
.A(n_2035),
.B(n_324),
.Y(n_2161)
);

NAND4xp75_ASAP7_75t_SL g2162 ( 
.A(n_2063),
.B(n_2044),
.C(n_2072),
.D(n_2027),
.Y(n_2162)
);

XNOR2xp5_ASAP7_75t_L g2163 ( 
.A(n_2103),
.B(n_326),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2024),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2050),
.Y(n_2165)
);

XOR2x2_ASAP7_75t_L g2166 ( 
.A(n_2054),
.B(n_327),
.Y(n_2166)
);

XOR2x2_ASAP7_75t_L g2167 ( 
.A(n_2029),
.B(n_328),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2046),
.Y(n_2168)
);

XNOR2xp5_ASAP7_75t_L g2169 ( 
.A(n_2039),
.B(n_2055),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2056),
.B(n_328),
.Y(n_2170)
);

NAND3xp33_ASAP7_75t_L g2171 ( 
.A(n_2043),
.B(n_329),
.C(n_330),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2099),
.B(n_329),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2100),
.B(n_330),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2037),
.B(n_331),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2090),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2088),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2052),
.B(n_332),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2020),
.Y(n_2178)
);

NAND4xp75_ASAP7_75t_L g2179 ( 
.A(n_2083),
.B(n_2033),
.C(n_2047),
.D(n_2093),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_2061),
.Y(n_2180)
);

XOR2xp5_ASAP7_75t_L g2181 ( 
.A(n_2025),
.B(n_504),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2084),
.B(n_2070),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2066),
.B(n_332),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2098),
.B(n_333),
.Y(n_2184)
);

NAND4xp75_ASAP7_75t_SL g2185 ( 
.A(n_2014),
.B(n_335),
.C(n_333),
.D(n_334),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2086),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2049),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2092),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2097),
.Y(n_2189)
);

NOR4xp25_ASAP7_75t_L g2190 ( 
.A(n_2018),
.B(n_338),
.C(n_336),
.D(n_337),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2082),
.B(n_338),
.Y(n_2191)
);

NAND4xp75_ASAP7_75t_SL g2192 ( 
.A(n_2106),
.B(n_341),
.C(n_339),
.D(n_340),
.Y(n_2192)
);

BUFx3_ASAP7_75t_L g2193 ( 
.A(n_2071),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2075),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2057),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_2017),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2010),
.Y(n_2197)
);

XNOR2xp5_ASAP7_75t_L g2198 ( 
.A(n_2034),
.B(n_341),
.Y(n_2198)
);

NAND4xp75_ASAP7_75t_L g2199 ( 
.A(n_2094),
.B(n_344),
.C(n_342),
.D(n_343),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2010),
.B(n_343),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2010),
.B(n_344),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2105),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2010),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_2042),
.B(n_345),
.Y(n_2204)
);

XNOR2x1_ASAP7_75t_L g2205 ( 
.A(n_2034),
.B(n_345),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2105),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2010),
.Y(n_2207)
);

CKINVDCx20_ASAP7_75t_R g2208 ( 
.A(n_2076),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2105),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2105),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2137),
.B(n_346),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2123),
.B(n_346),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2160),
.B(n_347),
.Y(n_2213)
);

XOR2xp5_ASAP7_75t_L g2214 ( 
.A(n_2205),
.B(n_348),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2117),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_2165),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2196),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2209),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2113),
.Y(n_2219)
);

XOR2x2_ASAP7_75t_L g2220 ( 
.A(n_2112),
.B(n_349),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2125),
.B(n_349),
.Y(n_2221)
);

XOR2x2_ASAP7_75t_L g2222 ( 
.A(n_2156),
.B(n_350),
.Y(n_2222)
);

INVxp67_ASAP7_75t_L g2223 ( 
.A(n_2204),
.Y(n_2223)
);

XNOR2xp5_ASAP7_75t_L g2224 ( 
.A(n_2120),
.B(n_350),
.Y(n_2224)
);

NOR2x1_ASAP7_75t_L g2225 ( 
.A(n_2131),
.B(n_351),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2202),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2206),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_2119),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2144),
.B(n_352),
.Y(n_2229)
);

XNOR2xp5_ASAP7_75t_L g2230 ( 
.A(n_2198),
.B(n_352),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2179),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_2231)
);

NOR2x1_ASAP7_75t_R g2232 ( 
.A(n_2193),
.B(n_2182),
.Y(n_2232)
);

INVx2_ASAP7_75t_SL g2233 ( 
.A(n_2110),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2210),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2208),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2127),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2164),
.B(n_354),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2108),
.Y(n_2238)
);

OAI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2126),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2114),
.Y(n_2240)
);

INVx1_ASAP7_75t_SL g2241 ( 
.A(n_2130),
.Y(n_2241)
);

XNOR2xp5_ASAP7_75t_L g2242 ( 
.A(n_2163),
.B(n_357),
.Y(n_2242)
);

XOR2x2_ASAP7_75t_L g2243 ( 
.A(n_2116),
.B(n_358),
.Y(n_2243)
);

XOR2x2_ASAP7_75t_L g2244 ( 
.A(n_2162),
.B(n_2109),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2154),
.B(n_358),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2152),
.Y(n_2246)
);

XNOR2x1_ASAP7_75t_L g2247 ( 
.A(n_2169),
.B(n_360),
.Y(n_2247)
);

XNOR2x1_ASAP7_75t_L g2248 ( 
.A(n_2121),
.B(n_360),
.Y(n_2248)
);

NOR2x1_ASAP7_75t_R g2249 ( 
.A(n_2180),
.B(n_2189),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2131),
.Y(n_2250)
);

INVx2_ASAP7_75t_SL g2251 ( 
.A(n_2197),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_SL g2252 ( 
.A1(n_2161),
.A2(n_362),
.B1(n_359),
.B2(n_361),
.Y(n_2252)
);

XOR2x2_ASAP7_75t_L g2253 ( 
.A(n_2167),
.B(n_359),
.Y(n_2253)
);

INVxp67_ASAP7_75t_L g2254 ( 
.A(n_2175),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2203),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2132),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2136),
.Y(n_2257)
);

XNOR2xp5_ASAP7_75t_L g2258 ( 
.A(n_2166),
.B(n_361),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2132),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2159),
.B(n_363),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2135),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2139),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_2150),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2142),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2207),
.Y(n_2265)
);

XOR2x2_ASAP7_75t_L g2266 ( 
.A(n_2185),
.B(n_364),
.Y(n_2266)
);

OA22x2_ASAP7_75t_L g2267 ( 
.A1(n_2168),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_2267)
);

XNOR2xp5_ASAP7_75t_L g2268 ( 
.A(n_2147),
.B(n_365),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2148),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2155),
.Y(n_2270)
);

XNOR2xp5_ASAP7_75t_L g2271 ( 
.A(n_2181),
.B(n_366),
.Y(n_2271)
);

AO22x1_ASAP7_75t_L g2272 ( 
.A1(n_2146),
.A2(n_2177),
.B1(n_2176),
.B2(n_2140),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2149),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2157),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2274)
);

XOR2x2_ASAP7_75t_L g2275 ( 
.A(n_2192),
.B(n_2115),
.Y(n_2275)
);

XOR2x2_ASAP7_75t_L g2276 ( 
.A(n_2199),
.B(n_2158),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2107),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2111),
.Y(n_2278)
);

XNOR2xp5_ASAP7_75t_L g2279 ( 
.A(n_2122),
.B(n_368),
.Y(n_2279)
);

XNOR2x1_ASAP7_75t_SL g2280 ( 
.A(n_2183),
.B(n_369),
.Y(n_2280)
);

XOR2x2_ASAP7_75t_L g2281 ( 
.A(n_2118),
.B(n_370),
.Y(n_2281)
);

INVx1_ASAP7_75t_SL g2282 ( 
.A(n_2128),
.Y(n_2282)
);

INVx1_ASAP7_75t_SL g2283 ( 
.A(n_2138),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2200),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2201),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2129),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2187),
.Y(n_2287)
);

CKINVDCx16_ASAP7_75t_R g2288 ( 
.A(n_2149),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2141),
.Y(n_2289)
);

XOR2x2_ASAP7_75t_L g2290 ( 
.A(n_2170),
.B(n_370),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_2143),
.Y(n_2291)
);

OA22x2_ASAP7_75t_L g2292 ( 
.A1(n_2188),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2151),
.B(n_372),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2134),
.A2(n_2171),
.B1(n_2133),
.B2(n_2145),
.Y(n_2294)
);

OAI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2186),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2178),
.Y(n_2296)
);

XNOR2x1_ASAP7_75t_L g2297 ( 
.A(n_2174),
.B(n_374),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2124),
.B(n_375),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2191),
.B(n_2194),
.Y(n_2299)
);

INVx2_ASAP7_75t_SL g2300 ( 
.A(n_2195),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2172),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_2301)
);

XOR2x2_ASAP7_75t_L g2302 ( 
.A(n_2173),
.B(n_377),
.Y(n_2302)
);

XOR2x2_ASAP7_75t_L g2303 ( 
.A(n_2153),
.B(n_2184),
.Y(n_2303)
);

XNOR2xp5_ASAP7_75t_L g2304 ( 
.A(n_2190),
.B(n_378),
.Y(n_2304)
);

XOR2xp5_ASAP7_75t_L g2305 ( 
.A(n_2205),
.B(n_379),
.Y(n_2305)
);

XNOR2xp5_ASAP7_75t_L g2306 ( 
.A(n_2112),
.B(n_380),
.Y(n_2306)
);

XNOR2xp5_ASAP7_75t_L g2307 ( 
.A(n_2112),
.B(n_380),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2117),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2117),
.Y(n_2309)
);

INVxp67_ASAP7_75t_L g2310 ( 
.A(n_2165),
.Y(n_2310)
);

XNOR2xp5_ASAP7_75t_L g2311 ( 
.A(n_2112),
.B(n_381),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_2165),
.Y(n_2312)
);

XOR2x2_ASAP7_75t_L g2313 ( 
.A(n_2112),
.B(n_381),
.Y(n_2313)
);

OA22x2_ASAP7_75t_L g2314 ( 
.A1(n_2180),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2117),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2117),
.Y(n_2316)
);

XNOR2xp5_ASAP7_75t_L g2317 ( 
.A(n_2112),
.B(n_382),
.Y(n_2317)
);

INVxp67_ASAP7_75t_SL g2318 ( 
.A(n_2125),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2117),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_R g2320 ( 
.A(n_2208),
.B(n_383),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_2196),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2308),
.Y(n_2322)
);

OA22x2_ASAP7_75t_L g2323 ( 
.A1(n_2231),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2241),
.B(n_385),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2319),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2219),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2226),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2227),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2240),
.Y(n_2329)
);

HB1xp67_ASAP7_75t_L g2330 ( 
.A(n_2250),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2234),
.Y(n_2331)
);

OA22x2_ASAP7_75t_L g2332 ( 
.A1(n_2294),
.A2(n_2304),
.B1(n_2258),
.B2(n_2279),
.Y(n_2332)
);

OA22x2_ASAP7_75t_L g2333 ( 
.A1(n_2279),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_2333)
);

OAI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2225),
.A2(n_390),
.B1(n_387),
.B2(n_389),
.Y(n_2334)
);

OA22x2_ASAP7_75t_L g2335 ( 
.A1(n_2252),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2228),
.B(n_391),
.Y(n_2336)
);

INVx4_ASAP7_75t_L g2337 ( 
.A(n_2212),
.Y(n_2337)
);

INVx2_ASAP7_75t_SL g2338 ( 
.A(n_2233),
.Y(n_2338)
);

OAI22xp33_ASAP7_75t_SL g2339 ( 
.A1(n_2288),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_2339)
);

OA22x2_ASAP7_75t_L g2340 ( 
.A1(n_2306),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2249),
.Y(n_2341)
);

AOI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2239),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_2263),
.Y(n_2343)
);

AOI22x1_ASAP7_75t_L g2344 ( 
.A1(n_2280),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_SL g2345 ( 
.A1(n_2272),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2255),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2274),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2246),
.Y(n_2348)
);

OAI22x1_ASAP7_75t_SL g2349 ( 
.A1(n_2235),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2349)
);

INVx2_ASAP7_75t_SL g2350 ( 
.A(n_2273),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2236),
.Y(n_2351)
);

OA22x2_ASAP7_75t_L g2352 ( 
.A1(n_2307),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2320),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2261),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2215),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_2256),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2238),
.Y(n_2357)
);

OA22x2_ASAP7_75t_L g2358 ( 
.A1(n_2311),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_2358)
);

OA22x2_ASAP7_75t_L g2359 ( 
.A1(n_2317),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_2359)
);

AOI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2276),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_2360)
);

HB1xp67_ASAP7_75t_L g2361 ( 
.A(n_2259),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2282),
.Y(n_2362)
);

AO22x2_ASAP7_75t_L g2363 ( 
.A1(n_2287),
.A2(n_411),
.B1(n_408),
.B2(n_410),
.Y(n_2363)
);

XNOR2x1_ASAP7_75t_L g2364 ( 
.A(n_2248),
.B(n_411),
.Y(n_2364)
);

OA22x2_ASAP7_75t_L g2365 ( 
.A1(n_2214),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2217),
.Y(n_2366)
);

INVxp33_ASAP7_75t_L g2367 ( 
.A(n_2232),
.Y(n_2367)
);

AOI22x1_ASAP7_75t_L g2368 ( 
.A1(n_2305),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_2368)
);

OA22x2_ASAP7_75t_L g2369 ( 
.A1(n_2216),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2309),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2315),
.Y(n_2371)
);

BUFx2_ASAP7_75t_L g2372 ( 
.A(n_2318),
.Y(n_2372)
);

OA22x2_ASAP7_75t_L g2373 ( 
.A1(n_2310),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2244),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_2374)
);

OA22x2_ASAP7_75t_L g2375 ( 
.A1(n_2312),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_2375)
);

OA22x2_ASAP7_75t_L g2376 ( 
.A1(n_2254),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2316),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_2321),
.Y(n_2378)
);

OA22x2_ASAP7_75t_L g2379 ( 
.A1(n_2268),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2300),
.Y(n_2380)
);

AOI22x1_ASAP7_75t_L g2381 ( 
.A1(n_2224),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2251),
.Y(n_2382)
);

OA22x2_ASAP7_75t_L g2383 ( 
.A1(n_2230),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_2383)
);

OA22x2_ASAP7_75t_L g2384 ( 
.A1(n_2299),
.A2(n_431),
.B1(n_428),
.B2(n_430),
.Y(n_2384)
);

OA22x2_ASAP7_75t_L g2385 ( 
.A1(n_2301),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_2385)
);

XOR2x2_ASAP7_75t_L g2386 ( 
.A(n_2243),
.B(n_432),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2265),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2218),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2275),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_2389)
);

INVx3_ASAP7_75t_SL g2390 ( 
.A(n_2303),
.Y(n_2390)
);

OA22x2_ASAP7_75t_L g2391 ( 
.A1(n_2271),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_2391)
);

XNOR2x1_ASAP7_75t_L g2392 ( 
.A(n_2253),
.B(n_436),
.Y(n_2392)
);

XOR2x2_ASAP7_75t_L g2393 ( 
.A(n_2222),
.B(n_437),
.Y(n_2393)
);

OA22x2_ASAP7_75t_L g2394 ( 
.A1(n_2242),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2262),
.Y(n_2395)
);

XOR2x2_ASAP7_75t_L g2396 ( 
.A(n_2220),
.B(n_438),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_2245),
.Y(n_2397)
);

AOI22x1_ASAP7_75t_L g2398 ( 
.A1(n_2286),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_2398)
);

AOI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2281),
.A2(n_443),
.B1(n_440),
.B2(n_442),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2264),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2289),
.Y(n_2401)
);

XNOR2xp5_ASAP7_75t_L g2402 ( 
.A(n_2313),
.B(n_443),
.Y(n_2402)
);

OA22x2_ASAP7_75t_L g2403 ( 
.A1(n_2257),
.A2(n_447),
.B1(n_444),
.B2(n_446),
.Y(n_2403)
);

XOR2x2_ASAP7_75t_L g2404 ( 
.A(n_2247),
.B(n_447),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_2269),
.Y(n_2405)
);

OA22x2_ASAP7_75t_L g2406 ( 
.A1(n_2283),
.A2(n_2291),
.B1(n_2223),
.B2(n_2278),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2270),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2295),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2267),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_2409)
);

BUFx2_ASAP7_75t_L g2410 ( 
.A(n_2284),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2277),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2285),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2221),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2213),
.B(n_452),
.Y(n_2414)
);

AOI22x1_ASAP7_75t_L g2415 ( 
.A1(n_2293),
.A2(n_2302),
.B1(n_2314),
.B2(n_2292),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2260),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2211),
.Y(n_2417)
);

OA22x2_ASAP7_75t_L g2418 ( 
.A1(n_2298),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_2418)
);

AOI22x1_ASAP7_75t_L g2419 ( 
.A1(n_2266),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_2419)
);

AOI22x1_ASAP7_75t_L g2420 ( 
.A1(n_2290),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_2420)
);

AOI22x1_ASAP7_75t_SL g2421 ( 
.A1(n_2297),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_2421)
);

BUFx3_ASAP7_75t_L g2422 ( 
.A(n_2229),
.Y(n_2422)
);

CKINVDCx16_ASAP7_75t_R g2423 ( 
.A(n_2237),
.Y(n_2423)
);

XNOR2x1_ASAP7_75t_L g2424 ( 
.A(n_2248),
.B(n_460),
.Y(n_2424)
);

OA22x2_ASAP7_75t_L g2425 ( 
.A1(n_2231),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2308),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2233),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_SL g2428 ( 
.A(n_2232),
.B(n_461),
.Y(n_2428)
);

XOR2x2_ASAP7_75t_L g2429 ( 
.A(n_2243),
.B(n_462),
.Y(n_2429)
);

XNOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2248),
.B(n_463),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_2233),
.Y(n_2431)
);

OA22x2_ASAP7_75t_L g2432 ( 
.A1(n_2231),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2308),
.Y(n_2433)
);

OA22x2_ASAP7_75t_L g2434 ( 
.A1(n_2231),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_2434)
);

AND2x4_ASAP7_75t_L g2435 ( 
.A(n_2216),
.B(n_468),
.Y(n_2435)
);

OA22x2_ASAP7_75t_L g2436 ( 
.A1(n_2231),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2308),
.Y(n_2437)
);

OA22x2_ASAP7_75t_L g2438 ( 
.A1(n_2231),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2308),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2308),
.Y(n_2440)
);

AOI22x1_ASAP7_75t_L g2441 ( 
.A1(n_2280),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2250),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2296),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2296),
.Y(n_2444)
);

OA22x2_ASAP7_75t_L g2445 ( 
.A1(n_2231),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_2445)
);

OA22x2_ASAP7_75t_L g2446 ( 
.A1(n_2231),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_2446)
);

AOI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_2294),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_2447)
);

BUFx2_ASAP7_75t_L g2448 ( 
.A(n_2263),
.Y(n_2448)
);

OA22x2_ASAP7_75t_L g2449 ( 
.A1(n_2231),
.A2(n_483),
.B1(n_480),
.B2(n_482),
.Y(n_2449)
);

OAI22xp5_ASAP7_75t_SL g2450 ( 
.A1(n_2214),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_2450)
);

INVx2_ASAP7_75t_SL g2451 ( 
.A(n_2233),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2308),
.Y(n_2452)
);

XOR2x2_ASAP7_75t_L g2453 ( 
.A(n_2243),
.B(n_485),
.Y(n_2453)
);

OAI22x1_ASAP7_75t_SL g2454 ( 
.A1(n_2241),
.A2(n_487),
.B1(n_488),
.B2(n_507),
.Y(n_2454)
);

OA22x2_ASAP7_75t_L g2455 ( 
.A1(n_2231),
.A2(n_487),
.B1(n_488),
.B2(n_508),
.Y(n_2455)
);

OA22x2_ASAP7_75t_L g2456 ( 
.A1(n_2231),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2294),
.A2(n_517),
.B1(n_512),
.B2(n_513),
.Y(n_2457)
);

OA22x2_ASAP7_75t_L g2458 ( 
.A1(n_2231),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_2458)
);

OA22x2_ASAP7_75t_L g2459 ( 
.A1(n_2231),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_2459)
);

XNOR2xp5_ASAP7_75t_L g2460 ( 
.A(n_2222),
.B(n_524),
.Y(n_2460)
);

OA22x2_ASAP7_75t_L g2461 ( 
.A1(n_2231),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.Y(n_2461)
);

BUFx3_ASAP7_75t_L g2462 ( 
.A(n_2233),
.Y(n_2462)
);

OAI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2294),
.A2(n_534),
.B1(n_529),
.B2(n_532),
.Y(n_2463)
);

OA22x2_ASAP7_75t_L g2464 ( 
.A1(n_2231),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_2464)
);

XNOR2x1_ASAP7_75t_L g2465 ( 
.A(n_2248),
.B(n_538),
.Y(n_2465)
);

OA22x2_ASAP7_75t_L g2466 ( 
.A1(n_2231),
.A2(n_546),
.B1(n_539),
.B2(n_543),
.Y(n_2466)
);

OAI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2294),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_2467)
);

OA22x2_ASAP7_75t_L g2468 ( 
.A1(n_2231),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.Y(n_2468)
);

OA22x2_ASAP7_75t_L g2469 ( 
.A1(n_2231),
.A2(n_558),
.B1(n_555),
.B2(n_556),
.Y(n_2469)
);

AOI22xp5_ASAP7_75t_L g2470 ( 
.A1(n_2294),
.A2(n_567),
.B1(n_560),
.B2(n_566),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_2233),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2308),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2233),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2233),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2294),
.A2(n_571),
.B1(n_568),
.B2(n_570),
.Y(n_2475)
);

OA22x2_ASAP7_75t_L g2476 ( 
.A1(n_2231),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2263),
.Y(n_2477)
);

OA22x2_ASAP7_75t_L g2478 ( 
.A1(n_2231),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2320),
.Y(n_2479)
);

AO22x2_ASAP7_75t_L g2480 ( 
.A1(n_2250),
.A2(n_583),
.B1(n_580),
.B2(n_581),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2366),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2322),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2325),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2326),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2378),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2327),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_2343),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2448),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2328),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2331),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2390),
.B(n_584),
.Y(n_2491)
);

HB1xp67_ASAP7_75t_L g2492 ( 
.A(n_2372),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2477),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2426),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2433),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2431),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2462),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2437),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2427),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2439),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2440),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2452),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2473),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2472),
.Y(n_2504)
);

INVx1_ASAP7_75t_SL g2505 ( 
.A(n_2353),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2351),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2338),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2479),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2354),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2348),
.Y(n_2510)
);

INVx4_ASAP7_75t_SL g2511 ( 
.A(n_2349),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2411),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2412),
.Y(n_2513)
);

INVxp67_ASAP7_75t_L g2514 ( 
.A(n_2428),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2401),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2395),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2451),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2400),
.Y(n_2518)
);

INVxp67_ASAP7_75t_SL g2519 ( 
.A(n_2341),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2355),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2471),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2370),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2474),
.Y(n_2523)
);

INVxp33_ASAP7_75t_L g2524 ( 
.A(n_2367),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2405),
.B(n_587),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2406),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2371),
.Y(n_2527)
);

OA22x2_ASAP7_75t_L g2528 ( 
.A1(n_2447),
.A2(n_590),
.B1(n_588),
.B2(n_589),
.Y(n_2528)
);

INVx2_ASAP7_75t_SL g2529 ( 
.A(n_2435),
.Y(n_2529)
);

INVx1_ASAP7_75t_SL g2530 ( 
.A(n_2362),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2357),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2377),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2388),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2330),
.Y(n_2534)
);

CKINVDCx16_ASAP7_75t_R g2535 ( 
.A(n_2421),
.Y(n_2535)
);

INVx2_ASAP7_75t_SL g2536 ( 
.A(n_2350),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2356),
.Y(n_2537)
);

INVxp67_ASAP7_75t_SL g2538 ( 
.A(n_2345),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2361),
.Y(n_2539)
);

INVxp33_ASAP7_75t_SL g2540 ( 
.A(n_2450),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2442),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2387),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2410),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2443),
.Y(n_2544)
);

BUFx4f_ASAP7_75t_SL g2545 ( 
.A(n_2414),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2444),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2329),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2346),
.Y(n_2548)
);

INVxp67_ASAP7_75t_SL g2549 ( 
.A(n_2454),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2380),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2382),
.Y(n_2551)
);

INVx1_ASAP7_75t_SL g2552 ( 
.A(n_2403),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2413),
.Y(n_2553)
);

HB1xp67_ASAP7_75t_L g2554 ( 
.A(n_2407),
.Y(n_2554)
);

BUFx2_ASAP7_75t_L g2555 ( 
.A(n_2337),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2416),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2417),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2397),
.Y(n_2558)
);

CKINVDCx20_ASAP7_75t_R g2559 ( 
.A(n_2423),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2363),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2422),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2332),
.A2(n_595),
.B1(n_592),
.B2(n_593),
.Y(n_2562)
);

HB1xp67_ASAP7_75t_L g2563 ( 
.A(n_2369),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2373),
.Y(n_2564)
);

XNOR2x2_ASAP7_75t_L g2565 ( 
.A(n_2376),
.B(n_596),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2340),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2415),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2344),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2375),
.Y(n_2569)
);

AOI322xp5_ASAP7_75t_L g2570 ( 
.A1(n_2399),
.A2(n_2374),
.A3(n_2360),
.B1(n_2409),
.B2(n_2389),
.C1(n_2324),
.C2(n_2336),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2441),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2480),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2480),
.Y(n_2573)
);

INVx4_ASAP7_75t_L g2574 ( 
.A(n_2393),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2384),
.Y(n_2575)
);

HB1xp67_ASAP7_75t_L g2576 ( 
.A(n_2418),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2334),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2333),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2385),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2335),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2339),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2323),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2425),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2432),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2391),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2434),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2436),
.Y(n_2587)
);

HB1xp67_ASAP7_75t_L g2588 ( 
.A(n_2379),
.Y(n_2588)
);

INVxp67_ASAP7_75t_L g2589 ( 
.A(n_2419),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2420),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2438),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2445),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2365),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2383),
.Y(n_2594)
);

INVx1_ASAP7_75t_SL g2595 ( 
.A(n_2559),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2492),
.Y(n_2596)
);

AOI221xp5_ASAP7_75t_L g2597 ( 
.A1(n_2567),
.A2(n_2402),
.B1(n_2467),
.B2(n_2475),
.C(n_2463),
.Y(n_2597)
);

AOI221xp5_ASAP7_75t_L g2598 ( 
.A1(n_2538),
.A2(n_2347),
.B1(n_2342),
.B2(n_2408),
.C(n_2460),
.Y(n_2598)
);

OAI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2535),
.A2(n_2449),
.B1(n_2446),
.B2(n_2457),
.Y(n_2599)
);

AOI22xp5_ASAP7_75t_L g2600 ( 
.A1(n_2519),
.A2(n_2455),
.B1(n_2458),
.B2(n_2456),
.Y(n_2600)
);

NAND4xp75_ASAP7_75t_L g2601 ( 
.A(n_2562),
.B(n_2470),
.C(n_2429),
.D(n_2453),
.Y(n_2601)
);

OAI222xp33_ASAP7_75t_L g2602 ( 
.A1(n_2526),
.A2(n_2358),
.B1(n_2359),
.B2(n_2352),
.C1(n_2394),
.C2(n_2459),
.Y(n_2602)
);

INVx3_ASAP7_75t_L g2603 ( 
.A(n_2496),
.Y(n_2603)
);

AND4x1_ASAP7_75t_L g2604 ( 
.A(n_2491),
.B(n_2396),
.C(n_2386),
.D(n_2404),
.Y(n_2604)
);

NAND4xp75_ASAP7_75t_L g2605 ( 
.A(n_2581),
.B(n_2392),
.C(n_2368),
.D(n_2381),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2487),
.Y(n_2606)
);

OA22x2_ASAP7_75t_L g2607 ( 
.A1(n_2549),
.A2(n_2424),
.B1(n_2430),
.B2(n_2364),
.Y(n_2607)
);

OA22x2_ASAP7_75t_L g2608 ( 
.A1(n_2566),
.A2(n_2465),
.B1(n_2461),
.B2(n_2464),
.Y(n_2608)
);

INVx1_ASAP7_75t_SL g2609 ( 
.A(n_2505),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2542),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2482),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2483),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2484),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2486),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2489),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2555),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2524),
.A2(n_2466),
.B1(n_2469),
.B2(n_2468),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2490),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2494),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2495),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2498),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2500),
.Y(n_2622)
);

AOI22xp5_ASAP7_75t_L g2623 ( 
.A1(n_2585),
.A2(n_2476),
.B1(n_2478),
.B2(n_2398),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2501),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2497),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2502),
.Y(n_2626)
);

NOR2x1_ASAP7_75t_L g2627 ( 
.A(n_2568),
.B(n_598),
.Y(n_2627)
);

OAI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2563),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2504),
.Y(n_2629)
);

OA22x2_ASAP7_75t_L g2630 ( 
.A1(n_2588),
.A2(n_606),
.B1(n_602),
.B2(n_605),
.Y(n_2630)
);

AOI221xp5_ASAP7_75t_L g2631 ( 
.A1(n_2540),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.C(n_610),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2506),
.Y(n_2632)
);

INVxp67_ASAP7_75t_L g2633 ( 
.A(n_2576),
.Y(n_2633)
);

AOI22x1_ASAP7_75t_L g2634 ( 
.A1(n_2574),
.A2(n_615),
.B1(n_611),
.B2(n_614),
.Y(n_2634)
);

AND4x1_ASAP7_75t_L g2635 ( 
.A(n_2580),
.B(n_623),
.C(n_616),
.D(n_620),
.Y(n_2635)
);

AOI31xp33_ASAP7_75t_L g2636 ( 
.A1(n_2589),
.A2(n_629),
.A3(n_625),
.B(n_627),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_2530),
.Y(n_2637)
);

OAI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2552),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2509),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2510),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2516),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2518),
.Y(n_2642)
);

OAI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2560),
.A2(n_638),
.B1(n_635),
.B2(n_636),
.Y(n_2643)
);

OA22x2_ASAP7_75t_L g2644 ( 
.A1(n_2571),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_2644)
);

OAI22xp33_ASAP7_75t_L g2645 ( 
.A1(n_2572),
.A2(n_646),
.B1(n_643),
.B2(n_644),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2512),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2513),
.Y(n_2647)
);

OAI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2573),
.A2(n_652),
.B1(n_647),
.B2(n_651),
.Y(n_2648)
);

OA22x2_ASAP7_75t_L g2649 ( 
.A1(n_2578),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.Y(n_2649)
);

INVx2_ASAP7_75t_SL g2650 ( 
.A(n_2481),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2520),
.Y(n_2651)
);

OAI322xp33_ASAP7_75t_L g2652 ( 
.A1(n_2582),
.A2(n_657),
.A3(n_658),
.B1(n_659),
.B2(n_660),
.C1(n_661),
.C2(n_662),
.Y(n_2652)
);

AOI221xp5_ASAP7_75t_L g2653 ( 
.A1(n_2574),
.A2(n_670),
.B1(n_667),
.B2(n_669),
.C(n_673),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2522),
.Y(n_2654)
);

OAI22x1_ASAP7_75t_L g2655 ( 
.A1(n_2600),
.A2(n_2623),
.B1(n_2606),
.B2(n_2604),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2595),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_2637),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2633),
.A2(n_2577),
.B1(n_2584),
.B2(n_2583),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2617),
.A2(n_2608),
.B1(n_2599),
.B2(n_2605),
.Y(n_2659)
);

OAI22x1_ASAP7_75t_L g2660 ( 
.A1(n_2609),
.A2(n_2594),
.B1(n_2593),
.B2(n_2569),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2596),
.Y(n_2661)
);

INVxp33_ASAP7_75t_SL g2662 ( 
.A(n_2607),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2601),
.A2(n_2511),
.B1(n_2488),
.B2(n_2493),
.Y(n_2663)
);

OAI22x1_ASAP7_75t_L g2664 ( 
.A1(n_2650),
.A2(n_2564),
.B1(n_2575),
.B2(n_2579),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2603),
.Y(n_2665)
);

OAI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2598),
.A2(n_2587),
.B1(n_2591),
.B2(n_2586),
.Y(n_2666)
);

OAI22x1_ASAP7_75t_L g2667 ( 
.A1(n_2616),
.A2(n_2592),
.B1(n_2514),
.B2(n_2590),
.Y(n_2667)
);

OAI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2597),
.A2(n_2536),
.B1(n_2485),
.B2(n_2503),
.Y(n_2668)
);

OAI221xp5_ASAP7_75t_L g2669 ( 
.A1(n_2625),
.A2(n_2570),
.B1(n_2558),
.B2(n_2543),
.C(n_2539),
.Y(n_2669)
);

OAI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2630),
.A2(n_2499),
.B1(n_2517),
.B2(n_2507),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2651),
.Y(n_2671)
);

A2O1A1Ixp33_ASAP7_75t_L g2672 ( 
.A1(n_2627),
.A2(n_2511),
.B(n_2537),
.C(n_2534),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2654),
.Y(n_2673)
);

INVxp33_ASAP7_75t_SL g2674 ( 
.A(n_2649),
.Y(n_2674)
);

AO22x2_ASAP7_75t_L g2675 ( 
.A1(n_2611),
.A2(n_2561),
.B1(n_2541),
.B2(n_2521),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2612),
.Y(n_2676)
);

OAI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2636),
.A2(n_2523),
.B1(n_2531),
.B2(n_2529),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2613),
.Y(n_2678)
);

OAI22x1_ASAP7_75t_L g2679 ( 
.A1(n_2635),
.A2(n_2551),
.B1(n_2550),
.B2(n_2525),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_2610),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2647),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2614),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2615),
.Y(n_2683)
);

OAI22x1_ASAP7_75t_L g2684 ( 
.A1(n_2634),
.A2(n_2525),
.B1(n_2553),
.B2(n_2565),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2618),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_SL g2686 ( 
.A1(n_2628),
.A2(n_2528),
.B1(n_2545),
.B2(n_2554),
.Y(n_2686)
);

INVx1_ASAP7_75t_SL g2687 ( 
.A(n_2644),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2657),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2681),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2656),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2661),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2675),
.Y(n_2692)
);

AO22x2_ASAP7_75t_L g2693 ( 
.A1(n_2658),
.A2(n_2620),
.B1(n_2621),
.B2(n_2619),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2662),
.B(n_2557),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2663),
.B(n_2556),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2687),
.B(n_2622),
.Y(n_2696)
);

AOI221xp5_ASAP7_75t_L g2697 ( 
.A1(n_2659),
.A2(n_2602),
.B1(n_2624),
.B2(n_2629),
.C(n_2626),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2665),
.Y(n_2698)
);

OAI22xp33_ASAP7_75t_SL g2699 ( 
.A1(n_2674),
.A2(n_2632),
.B1(n_2640),
.B2(n_2639),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2675),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2664),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2684),
.A2(n_2653),
.B1(n_2631),
.B2(n_2638),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2671),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2673),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2676),
.Y(n_2705)
);

NOR3xp33_ASAP7_75t_L g2706 ( 
.A(n_2666),
.B(n_2642),
.C(n_2641),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2702),
.A2(n_2655),
.B1(n_2686),
.B2(n_2669),
.Y(n_2707)
);

NOR2x1_ASAP7_75t_L g2708 ( 
.A(n_2692),
.B(n_2672),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2688),
.Y(n_2709)
);

NOR2x2_ASAP7_75t_L g2710 ( 
.A(n_2698),
.B(n_2667),
.Y(n_2710)
);

INVx1_ASAP7_75t_SL g2711 ( 
.A(n_2694),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2701),
.B(n_2660),
.Y(n_2712)
);

INVxp67_ASAP7_75t_L g2713 ( 
.A(n_2693),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2689),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2690),
.Y(n_2715)
);

OAI22x1_ASAP7_75t_L g2716 ( 
.A1(n_2700),
.A2(n_2508),
.B1(n_2680),
.B2(n_2678),
.Y(n_2716)
);

NOR2xp67_ASAP7_75t_L g2717 ( 
.A(n_2713),
.B(n_2679),
.Y(n_2717)
);

AND2x4_ASAP7_75t_L g2718 ( 
.A(n_2709),
.B(n_2706),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2714),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2707),
.A2(n_2697),
.B1(n_2708),
.B2(n_2677),
.Y(n_2720)
);

HB1xp67_ASAP7_75t_L g2721 ( 
.A(n_2711),
.Y(n_2721)
);

NOR4xp25_ASAP7_75t_L g2722 ( 
.A(n_2712),
.B(n_2696),
.C(n_2695),
.D(n_2691),
.Y(n_2722)
);

NOR2x1_ASAP7_75t_L g2723 ( 
.A(n_2715),
.B(n_2703),
.Y(n_2723)
);

NOR4xp25_ASAP7_75t_L g2724 ( 
.A(n_2710),
.B(n_2705),
.C(n_2704),
.D(n_2682),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2716),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2721),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2720),
.A2(n_2693),
.B1(n_2670),
.B2(n_2668),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2718),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2717),
.B(n_2683),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2725),
.Y(n_2730)
);

BUFx3_ASAP7_75t_L g2731 ( 
.A(n_2719),
.Y(n_2731)
);

OAI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2727),
.A2(n_2533),
.B1(n_2515),
.B2(n_2685),
.Y(n_2732)
);

OAI22x1_ASAP7_75t_L g2733 ( 
.A1(n_2729),
.A2(n_2728),
.B1(n_2730),
.B2(n_2726),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2731),
.B(n_2723),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2734),
.Y(n_2735)
);

AOI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2735),
.A2(n_2732),
.B1(n_2699),
.B2(n_2733),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2736),
.Y(n_2737)
);

OAI22xp33_ASAP7_75t_L g2738 ( 
.A1(n_2737),
.A2(n_2646),
.B1(n_2724),
.B2(n_2722),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2738),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2738),
.Y(n_2740)
);

AOI221xp5_ASAP7_75t_L g2741 ( 
.A1(n_2740),
.A2(n_2643),
.B1(n_2648),
.B2(n_2645),
.C(n_2652),
.Y(n_2741)
);

AOI221x1_ASAP7_75t_L g2742 ( 
.A1(n_2739),
.A2(n_2527),
.B1(n_2532),
.B2(n_2546),
.C(n_2544),
.Y(n_2742)
);

AOI211xp5_ASAP7_75t_L g2743 ( 
.A1(n_2741),
.A2(n_2742),
.B(n_2547),
.C(n_2548),
.Y(n_2743)
);


endmodule