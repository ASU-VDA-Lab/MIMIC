module fake_netlist_5_1745_n_1730 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1730);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1730;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_7),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_115),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_21),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_42),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_81),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_112),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_45),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_58),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_17),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_27),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_68),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_7),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_17),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_61),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_9),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_55),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_58),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_104),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_106),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_69),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_103),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_59),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_36),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_143),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_35),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_82),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_160),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_55),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_60),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_96),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_87),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_86),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_49),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_149),
.Y(n_226)
);

BUFx8_ASAP7_75t_SL g227 ( 
.A(n_113),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_2),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_91),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_56),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_41),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_1),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_39),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_140),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_13),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_85),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_5),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_120),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_41),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_32),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_30),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_43),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_57),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_161),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_92),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_44),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_83),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_146),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_3),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_8),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_162),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_70),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_30),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_88),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_95),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_52),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_62),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_157),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_76),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_77),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_93),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_73),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_65),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_3),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_2),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_99),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_141),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_121),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_14),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_49),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_51),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_45),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_25),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_32),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_46),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_24),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_39),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_102),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_47),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_105),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_26),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_116),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_119),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_108),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_53),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_53),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_14),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_20),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_125),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_4),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_21),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_109),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_100),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_111),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_54),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_16),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_150),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_114),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_5),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_25),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_67),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_142),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_12),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_74),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_16),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_156),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_185),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_199),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_227),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_269),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_164),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_260),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_201),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_170),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_207),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_207),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_171),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_189),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_257),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_218),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_172),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_214),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_173),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_218),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_276),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_180),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_214),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_181),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_289),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_177),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_177),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_184),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_232),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_289),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_232),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_186),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_193),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_194),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_196),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_237),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_163),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_201),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_237),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_165),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_248),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_192),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_198),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_248),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_251),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_200),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_205),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_251),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_256),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_256),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_287),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_287),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_296),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_175),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_206),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_188),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_296),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_300),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_166),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_192),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_302),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_209),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_167),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_210),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_242),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_167),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_168),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_330),
.B(n_242),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

CKINVDCx8_ASAP7_75t_R g408 ( 
.A(n_339),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_334),
.Y(n_409)
);

AND2x2_ASAP7_75t_SL g410 ( 
.A(n_383),
.B(n_195),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_321),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_176),
.B(n_168),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_337),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_353),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_R g424 ( 
.A(n_323),
.B(n_212),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_352),
.A2(n_280),
.B1(n_245),
.B2(n_314),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_341),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_357),
.A2(n_225),
.B1(n_293),
.B2(n_301),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_279),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_383),
.B(n_273),
.Y(n_438)
);

AND2x6_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_195),
.Y(n_439)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_346),
.B(n_279),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_397),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_398),
.B(n_202),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_335),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_322),
.A2(n_223),
.B1(n_319),
.B2(n_317),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_335),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_336),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_371),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_371),
.A2(n_202),
.B(n_268),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_348),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_347),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_336),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_359),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_340),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_340),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_344),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_344),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_364),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_375),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_361),
.B(n_270),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_362),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_374),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_345),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_401),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_410),
.A2(n_365),
.B1(n_333),
.B2(n_437),
.Y(n_474)
);

INVx8_ASAP7_75t_L g475 ( 
.A(n_439),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_417),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx8_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_382),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_405),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_428),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_428),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_440),
.A2(n_342),
.B1(n_329),
.B2(n_293),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_345),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_413),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_410),
.B(n_393),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_440),
.B(n_395),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_403),
.B(n_442),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_410),
.B(n_387),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_409),
.B(n_343),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_436),
.B(n_270),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_438),
.B(n_176),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_402),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_436),
.B(n_238),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_418),
.B(n_355),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_412),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_431),
.B(n_360),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_451),
.A2(n_234),
.B1(n_253),
.B2(n_252),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_404),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_439),
.B(n_203),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_414),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g526 ( 
.A1(n_451),
.A2(n_331),
.B1(n_342),
.B2(n_231),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_436),
.B(n_255),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_456),
.B(n_370),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_450),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_461),
.B(n_373),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_470),
.B(n_471),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_411),
.B(n_215),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_420),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_411),
.B(n_216),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_415),
.B(n_217),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_416),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_415),
.B(n_220),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_441),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_416),
.A2(n_301),
.B1(n_225),
.B2(n_449),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_457),
.B(n_367),
.Y(n_545)
);

CKINVDCx6p67_ASAP7_75t_R g546 ( 
.A(n_420),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_441),
.B(n_221),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_441),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_425),
.B(n_367),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_449),
.B(n_197),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_450),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_450),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_450),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_433),
.A2(n_294),
.B1(n_197),
.B2(n_204),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_446),
.B(n_204),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_416),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_427),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_424),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_453),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_453),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_453),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_416),
.A2(n_235),
.B1(n_315),
.B2(n_311),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_419),
.A2(n_219),
.B(n_213),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

OA22x2_ASAP7_75t_L g572 ( 
.A1(n_425),
.A2(n_392),
.B1(n_391),
.B2(n_390),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_453),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_421),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_L g577 ( 
.A(n_439),
.B(n_224),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_422),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_433),
.B(n_213),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_439),
.A2(n_236),
.B1(n_241),
.B2(n_239),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_464),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_422),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_464),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_408),
.Y(n_585)
);

INVxp33_ASAP7_75t_L g586 ( 
.A(n_423),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_423),
.B(n_226),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_464),
.Y(n_588)
);

AOI21x1_ASAP7_75t_L g589 ( 
.A1(n_426),
.A2(n_230),
.B(n_219),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_464),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_464),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_429),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_427),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_429),
.B(n_432),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_439),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_432),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_434),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_434),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_435),
.B(n_230),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_439),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_435),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_408),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_443),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_443),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_444),
.B(n_349),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_444),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_445),
.B(n_326),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_445),
.B(n_229),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_427),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_439),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_447),
.B(n_249),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_430),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_452),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_458),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_447),
.B(n_273),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_448),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_448),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_454),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_454),
.B(n_250),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_510),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_484),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_525),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_493),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_493),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_505),
.B(n_254),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_568),
.B(n_192),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_490),
.B(n_459),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_504),
.B(n_192),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_235),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_564),
.B(n_263),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_544),
.B(n_604),
.Y(n_634)
);

AND2x2_ASAP7_75t_SL g635 ( 
.A(n_550),
.B(n_240),
.Y(n_635)
);

O2A1O1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_501),
.A2(n_459),
.B(n_469),
.C(n_467),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_240),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_607),
.B(n_258),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_586),
.B(n_169),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_509),
.B(n_174),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_523),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_536),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_545),
.B(n_460),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_560),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_516),
.B(n_264),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_473),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_574),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_607),
.B(n_258),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_529),
.B(n_267),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_620),
.B(n_272),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_514),
.A2(n_474),
.B1(n_482),
.B2(n_490),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_620),
.B(n_277),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_621),
.B(n_476),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_558),
.A2(n_274),
.B(n_311),
.C(n_306),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_484),
.B(n_259),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_514),
.A2(n_259),
.B1(n_294),
.B2(n_290),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_487),
.B(n_460),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_621),
.B(n_262),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_476),
.B(n_262),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_580),
.B(n_278),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_473),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_477),
.B(n_266),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_549),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_526),
.B(n_246),
.C(n_243),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_477),
.B(n_266),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_580),
.A2(n_579),
.B1(n_522),
.B2(n_597),
.C(n_572),
.Y(n_667)
);

AND3x1_ASAP7_75t_L g668 ( 
.A(n_522),
.B(n_379),
.C(n_376),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_514),
.A2(n_312),
.B1(n_307),
.B2(n_308),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_478),
.B(n_274),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_478),
.B(n_290),
.Y(n_671)
);

AO22x1_ASAP7_75t_L g672 ( 
.A1(n_550),
.A2(n_208),
.B1(n_211),
.B2(n_222),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_479),
.B(n_599),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_574),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_550),
.B(n_306),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_558),
.B(n_315),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_578),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_599),
.B(n_178),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_578),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_587),
.B(n_292),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_558),
.A2(n_469),
.B(n_467),
.C(n_472),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_514),
.A2(n_309),
.B1(n_182),
.B2(n_183),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_599),
.B(n_179),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_479),
.B(n_458),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_608),
.Y(n_687)
);

OA22x2_ASAP7_75t_L g688 ( 
.A1(n_579),
.A2(n_376),
.B1(n_392),
.B2(n_391),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_484),
.B(n_458),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_489),
.B(n_462),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_491),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_611),
.B(n_295),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_614),
.B(n_187),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_595),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_582),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_489),
.B(n_462),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_489),
.B(n_492),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_492),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_539),
.A2(n_378),
.B(n_377),
.C(n_379),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_622),
.B(n_190),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_534),
.B(n_188),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_514),
.B(n_191),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_605),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_595),
.Y(n_705)
);

BUFx8_ASAP7_75t_L g706 ( 
.A(n_546),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_492),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_593),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_593),
.B(n_297),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_519),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_511),
.B(n_188),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_600),
.B(n_462),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_512),
.A2(n_550),
.B1(n_538),
.B2(n_537),
.Y(n_713)
);

BUFx6f_ASAP7_75t_SL g714 ( 
.A(n_579),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_546),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_595),
.Y(n_716)
);

O2A1O1Ixp5_ASAP7_75t_L g717 ( 
.A1(n_542),
.A2(n_472),
.B(n_465),
.C(n_463),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_600),
.B(n_228),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_519),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_601),
.B(n_233),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_601),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_596),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_606),
.B(n_463),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_606),
.B(n_463),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_609),
.B(n_247),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_609),
.B(n_465),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_556),
.A2(n_265),
.B1(n_261),
.B2(n_281),
.C(n_275),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_608),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_619),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_535),
.B(n_271),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_618),
.B(n_298),
.C(n_283),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_540),
.B(n_303),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_610),
.B(n_286),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_539),
.B(n_465),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_596),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_572),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_488),
.B(n_472),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_488),
.B(n_430),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_495),
.B(n_497),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_495),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_596),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_497),
.B(n_430),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_498),
.B(n_430),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_518),
.B(n_390),
.C(n_389),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_585),
.B(n_377),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_498),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_572),
.B(n_316),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_506),
.B(n_430),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_506),
.B(n_430),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_515),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_515),
.B(n_430),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_521),
.B(n_530),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_547),
.B(n_320),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_527),
.B(n_288),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_527),
.B(n_192),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_532),
.B(n_188),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_533),
.B(n_483),
.Y(n_758)
);

NOR2x1p5_ASAP7_75t_L g759 ( 
.A(n_533),
.B(n_291),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_543),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_543),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_579),
.B(n_378),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_548),
.B(n_192),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_SL g764 ( 
.A(n_519),
.B(n_299),
.Y(n_764)
);

INVx6_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_548),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_524),
.A2(n_602),
.B1(n_570),
.B2(n_577),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_602),
.A2(n_192),
.B1(n_273),
.B2(n_318),
.Y(n_768)
);

AND2x6_ASAP7_75t_SL g769 ( 
.A(n_579),
.B(n_380),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_553),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_542),
.B(n_192),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_598),
.B(n_318),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_598),
.B(n_318),
.Y(n_773)
);

AND2x4_ASAP7_75t_SL g774 ( 
.A(n_602),
.B(n_318),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_557),
.B(n_192),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_496),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_589),
.B(n_613),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_553),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_589),
.A2(n_313),
.B1(n_384),
.B2(n_389),
.Y(n_779)
);

NAND2x1p5_ASAP7_75t_L g780 ( 
.A(n_613),
.B(n_385),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_559),
.B(n_386),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_559),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_570),
.B(n_285),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_570),
.A2(n_386),
.B(n_385),
.C(n_384),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_557),
.B(n_380),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_630),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_635),
.B(n_481),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_627),
.B(n_551),
.Y(n_788)
);

BUFx8_ASAP7_75t_L g789 ( 
.A(n_714),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_624),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_663),
.B(n_481),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_624),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_630),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_635),
.A2(n_555),
.B1(n_554),
.B2(n_561),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_644),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_676),
.B(n_598),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_676),
.B(n_603),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_642),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_687),
.B(n_485),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_713),
.B(n_603),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_624),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_647),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_760),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_651),
.B(n_603),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_728),
.B(n_551),
.Y(n_805)
);

AO21x1_ASAP7_75t_L g806 ( 
.A1(n_783),
.A2(n_779),
.B(n_784),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_661),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_728),
.B(n_552),
.Y(n_809)
);

AND2x6_ASAP7_75t_L g810 ( 
.A(n_710),
.B(n_531),
.Y(n_810)
);

AO22x1_ASAP7_75t_L g811 ( 
.A1(n_702),
.A2(n_640),
.B1(n_666),
.B2(n_733),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_677),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_634),
.A2(n_575),
.B1(n_561),
.B2(n_554),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_693),
.B(n_486),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_736),
.A2(n_667),
.B1(n_677),
.B2(n_688),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_693),
.A2(n_555),
.B1(n_565),
.B2(n_566),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_700),
.B(n_486),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_626),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_697),
.A2(n_734),
.B(n_673),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_674),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_700),
.B(n_616),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_683),
.A2(n_717),
.B(n_767),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_627),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_727),
.B(n_350),
.C(n_351),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_625),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_736),
.B(n_552),
.Y(n_826)
);

BUFx8_ASAP7_75t_L g827 ( 
.A(n_714),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_624),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_761),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_730),
.B(n_616),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_730),
.B(n_617),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_641),
.B(n_617),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_766),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_675),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_643),
.B(n_499),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_678),
.B(n_499),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_698),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_679),
.B(n_681),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_688),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_695),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_639),
.B(n_565),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_698),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_704),
.B(n_513),
.Y(n_843)
);

CKINVDCx11_ASAP7_75t_R g844 ( 
.A(n_703),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_677),
.A2(n_556),
.B1(n_557),
.B2(n_231),
.Y(n_845)
);

AOI22x1_ASAP7_75t_SL g846 ( 
.A1(n_715),
.A2(n_285),
.B1(n_284),
.B2(n_244),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_708),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_710),
.B(n_603),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_698),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_721),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_698),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_729),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_740),
.B(n_513),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_747),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_639),
.B(n_566),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_640),
.B(n_567),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_677),
.A2(n_571),
.B1(n_573),
.B2(n_575),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_770),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_765),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_703),
.B(n_556),
.Y(n_860)
);

NOR2x2_ASAP7_75t_L g861 ( 
.A(n_632),
.B(n_231),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_623),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_632),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_751),
.B(n_513),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_653),
.B(n_528),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_677),
.A2(n_783),
.B1(n_629),
.B2(n_779),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_680),
.B(n_528),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_778),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_759),
.B(n_762),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_762),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_628),
.B(n_573),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_680),
.B(n_528),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_719),
.B(n_531),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_701),
.A2(n_285),
.B1(n_284),
.B2(n_244),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_719),
.B(n_531),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_762),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_685),
.B(n_528),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_782),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_707),
.B(n_613),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_703),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_702),
.A2(n_657),
.B(n_636),
.C(n_733),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_685),
.B(n_581),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_684),
.A2(n_557),
.B1(n_244),
.B2(n_284),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_712),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_623),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_668),
.B(n_581),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_765),
.A2(n_496),
.B1(n_520),
.B2(n_517),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_711),
.B(n_231),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_745),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_745),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_694),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_656),
.A2(n_664),
.B1(n_660),
.B2(n_662),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_718),
.B(n_581),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_723),
.Y(n_894)
);

AOI21xp33_ASAP7_75t_L g895 ( 
.A1(n_757),
.A2(n_475),
.B(n_480),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_745),
.B(n_583),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_718),
.B(n_720),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_724),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_720),
.B(n_244),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_765),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_753),
.B(n_583),
.Y(n_901)
);

NOR2x2_ASAP7_75t_L g902 ( 
.A(n_632),
.B(n_769),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_744),
.B(n_755),
.C(n_725),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_707),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_748),
.B(n_475),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_725),
.B(n_583),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_758),
.B(n_584),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_706),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_637),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_705),
.Y(n_910)
);

OR2x4_ASAP7_75t_L g911 ( 
.A(n_755),
.B(n_284),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_726),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_638),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_706),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_746),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_659),
.A2(n_557),
.B1(n_285),
.B2(n_507),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_746),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_776),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_648),
.B(n_584),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_737),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_658),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_739),
.B(n_584),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_633),
.B(n_588),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_744),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_717),
.A2(n_738),
.B(n_750),
.Y(n_925)
);

INVx3_ASAP7_75t_SL g926 ( 
.A(n_774),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_781),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_672),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_691),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_771),
.A2(n_592),
.B(n_588),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_665),
.B(n_588),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_716),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_764),
.B(n_613),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_722),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_669),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_735),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_670),
.B(n_591),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_671),
.B(n_591),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_686),
.B(n_591),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_655),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_699),
.B(n_592),
.Y(n_941)
);

AND2x6_ASAP7_75t_SL g942 ( 
.A(n_756),
.B(n_763),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_741),
.Y(n_943)
);

OAI21xp33_ASAP7_75t_SL g944 ( 
.A1(n_645),
.A2(n_592),
.B(n_502),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_785),
.A2(n_557),
.B1(n_500),
.B2(n_502),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_689),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_690),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_775),
.A2(n_557),
.B1(n_500),
.B2(n_507),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_731),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_696),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_649),
.A2(n_709),
.B1(n_754),
.B2(n_692),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_655),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_682),
.B(n_520),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_654),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_742),
.B(n_613),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_743),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_768),
.B(n_494),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_631),
.A2(n_475),
.B1(n_480),
.B2(n_613),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_732),
.B(n_494),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_749),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_SL g961 ( 
.A1(n_780),
.A2(n_0),
.B1(n_8),
.B2(n_10),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_752),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_650),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_652),
.B(n_494),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_772),
.B(n_494),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_915),
.A2(n_777),
.B(n_746),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_859),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_897),
.B(n_773),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_844),
.Y(n_969)
);

AND2x2_ASAP7_75t_SL g970 ( 
.A(n_883),
.B(n_10),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_823),
.B(n_494),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_915),
.A2(n_746),
.B(n_475),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_818),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_859),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_856),
.A2(n_569),
.B(n_563),
.C(n_562),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_915),
.A2(n_480),
.B(n_562),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_869),
.B(n_503),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_914),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_909),
.B(n_503),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_891),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_866),
.A2(n_503),
.B1(n_480),
.B2(n_562),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_915),
.A2(n_563),
.B(n_541),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_917),
.A2(n_563),
.B(n_541),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_795),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_859),
.Y(n_985)
);

OAI321xp33_ASAP7_75t_L g986 ( 
.A1(n_935),
.A2(n_11),
.A3(n_15),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_909),
.B(n_503),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_866),
.A2(n_503),
.B1(n_18),
.B2(n_22),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_924),
.B(n_503),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_798),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_903),
.A2(n_541),
.B(n_562),
.C(n_563),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_917),
.A2(n_569),
.B(n_541),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_911),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_815),
.A2(n_11),
.B1(n_22),
.B2(n_23),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_SL g995 ( 
.A1(n_856),
.A2(n_855),
.B(n_841),
.C(n_822),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_825),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_925),
.A2(n_569),
.B(n_72),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_917),
.A2(n_612),
.B(n_508),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_815),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_888),
.B(n_28),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_811),
.B(n_31),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_801),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_900),
.B(n_612),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_SL g1004 ( 
.A1(n_874),
.A2(n_885),
.B1(n_862),
.B2(n_961),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_900),
.B(n_612),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_SL g1006 ( 
.A(n_824),
.B(n_33),
.C(n_34),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_881),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_917),
.A2(n_612),
.B(n_508),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_810),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_802),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_881),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_800),
.A2(n_508),
.B(n_615),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_900),
.B(n_508),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_910),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_800),
.A2(n_615),
.B(n_594),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_820),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_845),
.A2(n_839),
.B1(n_892),
.B2(n_812),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_819),
.A2(n_615),
.B(n_594),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_834),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_845),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_900),
.B(n_928),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_927),
.B(n_44),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_804),
.A2(n_615),
.B(n_594),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_848),
.A2(n_615),
.B(n_594),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_910),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_804),
.A2(n_615),
.B(n_594),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_904),
.A2(n_80),
.B(n_135),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_869),
.B(n_79),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_791),
.B(n_47),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_913),
.B(n_50),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_921),
.B(n_50),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_904),
.A2(n_84),
.B(n_127),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_791),
.B(n_51),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_786),
.B(n_89),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_899),
.A2(n_52),
.B(n_54),
.C(n_56),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_841),
.A2(n_57),
.B(n_59),
.C(n_63),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_SL g1037 ( 
.A(n_926),
.B(n_71),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_SL g1038 ( 
.A(n_812),
.B(n_75),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_848),
.A2(n_78),
.B(n_90),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_932),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_840),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_867),
.A2(n_97),
.B(n_98),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_930),
.A2(n_101),
.B(n_107),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_963),
.A2(n_123),
.B1(n_124),
.B2(n_148),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_884),
.B(n_894),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_832),
.B(n_949),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_793),
.B(n_896),
.Y(n_1047)
);

CKINVDCx11_ASAP7_75t_R g1048 ( 
.A(n_914),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_932),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_880),
.B(n_908),
.Y(n_1050)
);

BUFx8_ASAP7_75t_L g1051 ( 
.A(n_880),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_798),
.B(n_889),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_943),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_839),
.A2(n_892),
.B1(n_812),
.B2(n_954),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_812),
.A2(n_954),
.B1(n_787),
.B2(n_838),
.Y(n_1055)
);

CKINVDCx16_ASAP7_75t_R g1056 ( 
.A(n_889),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_863),
.B(n_890),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_837),
.B(n_842),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_814),
.A2(n_817),
.B1(n_912),
.B2(n_920),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_898),
.B(n_855),
.Y(n_1060)
);

AO22x1_ASAP7_75t_L g1061 ( 
.A1(n_890),
.A2(n_876),
.B1(n_870),
.B2(n_926),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_870),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_L g1063 ( 
.A(n_951),
.B(n_847),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_872),
.A2(n_877),
.B(n_882),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_850),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_896),
.B(n_788),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_852),
.B(n_854),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_837),
.B(n_842),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_876),
.A2(n_886),
.B1(n_923),
.B2(n_901),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_805),
.B(n_809),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_953),
.A2(n_871),
.B(n_923),
.C(n_830),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_860),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_803),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_943),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_835),
.B(n_805),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_809),
.B(n_940),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_L g1077 ( 
.A1(n_806),
.A2(n_831),
.B(n_821),
.C(n_797),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_948),
.A2(n_945),
.B1(n_860),
.B2(n_868),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_796),
.A2(n_797),
.B(n_931),
.Y(n_1079)
);

AOI21x1_ASAP7_75t_L g1080 ( 
.A1(n_893),
.A2(n_906),
.B(n_907),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_801),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_799),
.B(n_826),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_860),
.B(n_886),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_803),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_826),
.B(n_946),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_801),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_829),
.B(n_833),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_789),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_829),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_948),
.A2(n_945),
.B1(n_878),
.B2(n_858),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_947),
.B(n_950),
.Y(n_1091)
);

AO21x2_ASAP7_75t_L g1092 ( 
.A1(n_887),
.A2(n_941),
.B(n_907),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_833),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_858),
.B(n_878),
.Y(n_1094)
);

AND2x6_ASAP7_75t_SL g1095 ( 
.A(n_846),
.B(n_905),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_796),
.A2(n_938),
.B(n_937),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_929),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_895),
.A2(n_865),
.B(n_939),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_789),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_934),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_965),
.A2(n_873),
.B(n_875),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_918),
.B(n_953),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_873),
.A2(n_875),
.B(n_959),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_810),
.Y(n_1104)
);

INVx4_ASAP7_75t_SL g1105 ( 
.A(n_810),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_936),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_916),
.A2(n_887),
.B1(n_883),
.B2(n_952),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_959),
.A2(n_922),
.B(n_879),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_871),
.A2(n_905),
.B1(n_964),
.B2(n_940),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_964),
.A2(n_956),
.B(n_962),
.C(n_960),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_960),
.B(n_952),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_807),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_808),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_836),
.A2(n_864),
.B(n_853),
.C(n_843),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_879),
.A2(n_955),
.B(n_919),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_911),
.B(n_942),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_1001),
.A2(n_902),
.B1(n_813),
.B2(n_861),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1089),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_L g1119 ( 
.A(n_990),
.B(n_851),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1077),
.A2(n_944),
.B(n_816),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1063),
.A2(n_916),
.B(n_794),
.C(n_857),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1046),
.B(n_827),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_973),
.B(n_790),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1071),
.A2(n_958),
.B(n_851),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1045),
.B(n_790),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_970),
.A2(n_828),
.B1(n_849),
.B2(n_792),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1000),
.B(n_792),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1052),
.B(n_828),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1047),
.B(n_828),
.Y(n_1129)
);

BUFx4f_ASAP7_75t_SL g1130 ( 
.A(n_1051),
.Y(n_1130)
);

CKINVDCx16_ASAP7_75t_R g1131 ( 
.A(n_969),
.Y(n_1131)
);

AO22x2_ASAP7_75t_L g1132 ( 
.A1(n_988),
.A2(n_957),
.B1(n_810),
.B2(n_933),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1047),
.B(n_849),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1108),
.A2(n_957),
.B(n_1096),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1062),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1059),
.A2(n_957),
.B(n_1060),
.Y(n_1136)
);

OAI21xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1091),
.A2(n_957),
.B(n_1022),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_1038),
.B(n_957),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1018),
.A2(n_1024),
.B(n_1015),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1101),
.A2(n_1026),
.B(n_1023),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1055),
.A2(n_1017),
.A3(n_1054),
.B(n_1079),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1082),
.B(n_1085),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1115),
.A2(n_1103),
.B(n_1012),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_984),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_981),
.A2(n_1110),
.B(n_1114),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1029),
.A2(n_1033),
.B(n_968),
.C(n_1011),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1080),
.A2(n_1043),
.B(n_976),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_980),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1035),
.B(n_1006),
.C(n_1007),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1055),
.A2(n_1102),
.B(n_1054),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1087),
.B(n_1094),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1017),
.A2(n_1069),
.B(n_1107),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1030),
.A2(n_1031),
.B(n_1067),
.Y(n_1153)
);

AOI211x1_ASAP7_75t_L g1154 ( 
.A1(n_994),
.A2(n_999),
.B(n_1020),
.C(n_1078),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1028),
.B(n_1056),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1111),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_991),
.A2(n_1090),
.B(n_1109),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1010),
.B(n_1016),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1039),
.A2(n_966),
.B(n_972),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1090),
.A2(n_982),
.B(n_992),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1048),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1050),
.Y(n_1162)
);

AOI221xp5_ASAP7_75t_L g1163 ( 
.A1(n_986),
.A2(n_1020),
.B1(n_999),
.B2(n_994),
.C(n_1116),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1038),
.A2(n_1009),
.B(n_1104),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_977),
.B(n_1028),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1075),
.B(n_1070),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1086),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1036),
.A2(n_1083),
.B1(n_1078),
.B2(n_1042),
.C(n_1004),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_L g1169 ( 
.A(n_986),
.B(n_1037),
.C(n_1061),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_989),
.A2(n_1093),
.A3(n_1084),
.B(n_1073),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1019),
.B(n_1041),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_975),
.A2(n_1032),
.B(n_1027),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1065),
.B(n_987),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_1076),
.B(n_1072),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_983),
.A2(n_1008),
.B(n_998),
.Y(n_1175)
);

CKINVDCx16_ASAP7_75t_R g1176 ( 
.A(n_1099),
.Y(n_1176)
);

CKINVDCx14_ASAP7_75t_R g1177 ( 
.A(n_993),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_979),
.A2(n_1049),
.B(n_1040),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_977),
.B(n_985),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1014),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1003),
.A2(n_1005),
.B(n_1013),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1057),
.B(n_971),
.Y(n_1182)
);

NAND3x1_ASAP7_75t_L g1183 ( 
.A(n_1044),
.B(n_1097),
.C(n_978),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1025),
.A2(n_1053),
.A3(n_1074),
.B(n_1106),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1051),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1092),
.A2(n_1100),
.A3(n_1113),
.B(n_1112),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1058),
.A2(n_1068),
.B(n_1066),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1021),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1088),
.A2(n_1034),
.B1(n_974),
.B2(n_967),
.C(n_985),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1009),
.A2(n_1104),
.B(n_1068),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1081),
.A2(n_1105),
.A3(n_1002),
.B(n_1058),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_993),
.B(n_967),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1002),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1105),
.A2(n_1095),
.B(n_1081),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1086),
.A2(n_967),
.B1(n_974),
.B2(n_1105),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1086),
.A2(n_974),
.B(n_978),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_997),
.A2(n_1018),
.B(n_1024),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1060),
.B(n_897),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_SL g1199 ( 
.A(n_970),
.B(n_1038),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1089),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_997),
.A2(n_1018),
.B(n_1024),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1077),
.A2(n_1071),
.B(n_1096),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1077),
.A2(n_1098),
.B(n_822),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_977),
.B(n_1047),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_997),
.A2(n_1018),
.B(n_1024),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1045),
.B(n_897),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1046),
.B(n_899),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1045),
.B(n_897),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1046),
.B(n_321),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1063),
.A2(n_897),
.B(n_903),
.C(n_881),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1060),
.B(n_897),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1108),
.A2(n_1080),
.B(n_1079),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1086),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_995),
.Y(n_1214)
);

INVx3_ASAP7_75t_SL g1215 ( 
.A(n_996),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1046),
.B(n_897),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_973),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1045),
.B(n_897),
.Y(n_1218)
);

O2A1O1Ixp5_ASAP7_75t_L g1219 ( 
.A1(n_968),
.A2(n_897),
.B(n_811),
.C(n_903),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1060),
.B(n_897),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_995),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_995),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_973),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_996),
.B(n_825),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1009),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_980),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1063),
.A2(n_897),
.B(n_903),
.C(n_881),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1060),
.B(n_897),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1055),
.A2(n_806),
.A3(n_1071),
.B(n_1098),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_970),
.A2(n_988),
.B1(n_1060),
.B2(n_866),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1051),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1055),
.A2(n_806),
.A3(n_1071),
.B(n_1098),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1055),
.A2(n_806),
.A3(n_1071),
.B(n_1098),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_969),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1107),
.A2(n_1071),
.B(n_988),
.Y(n_1235)
);

CKINVDCx16_ASAP7_75t_R g1236 ( 
.A(n_969),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_995),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1045),
.B(n_897),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1063),
.A2(n_897),
.B(n_903),
.C(n_881),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1055),
.A2(n_806),
.A3(n_1071),
.B(n_1098),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1046),
.B(n_899),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1045),
.B(n_897),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1108),
.A2(n_1080),
.B(n_1079),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1077),
.A2(n_1071),
.B(n_1096),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_995),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1089),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1089),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1077),
.A2(n_1071),
.B(n_1096),
.Y(n_1248)
);

AOI211x1_ASAP7_75t_L g1249 ( 
.A1(n_994),
.A2(n_999),
.B(n_1020),
.C(n_988),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_973),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_970),
.A2(n_988),
.B1(n_1060),
.B2(n_866),
.Y(n_1251)
);

OAI21xp33_ASAP7_75t_SL g1252 ( 
.A1(n_970),
.A2(n_866),
.B(n_676),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_980),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1064),
.A2(n_1098),
.B(n_995),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1167),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1138),
.A2(n_1134),
.B(n_1164),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1158),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1234),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1171),
.Y(n_1259)
);

OR2x6_ASAP7_75t_L g1260 ( 
.A(n_1235),
.B(n_1249),
.Y(n_1260)
);

OR2x6_ASAP7_75t_L g1261 ( 
.A(n_1154),
.B(n_1190),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1138),
.A2(n_1221),
.B(n_1214),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1144),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1206),
.B(n_1208),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1216),
.B(n_1250),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1218),
.B(n_1238),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1184),
.Y(n_1267)
);

OAI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1199),
.A2(n_1146),
.B1(n_1252),
.B2(n_1163),
.C(n_1153),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1199),
.A2(n_1251),
.B(n_1230),
.C(n_1152),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1180),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1170),
.Y(n_1271)
);

AO21x1_ASAP7_75t_L g1272 ( 
.A1(n_1230),
.A2(n_1251),
.B(n_1169),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1148),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1223),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1222),
.A2(n_1245),
.A3(n_1254),
.B(n_1237),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1219),
.A2(n_1227),
.B(n_1239),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1128),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1186),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1191),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1149),
.B(n_1168),
.C(n_1210),
.Y(n_1280)
);

INVx3_ASAP7_75t_SL g1281 ( 
.A(n_1162),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1191),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1242),
.B(n_1198),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1250),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1170),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1209),
.B(n_1207),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1159),
.A2(n_1139),
.B(n_1175),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1241),
.B(n_1198),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1211),
.B(n_1220),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1127),
.B(n_1155),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1131),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1147),
.A2(n_1143),
.B(n_1140),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1160),
.A2(n_1212),
.B(n_1243),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1226),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1151),
.B(n_1211),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1192),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1161),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1156),
.B(n_1204),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1220),
.B(n_1228),
.Y(n_1299)
);

OAI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1149),
.A2(n_1228),
.B1(n_1122),
.B2(n_1152),
.C(n_1137),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1177),
.B(n_1215),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1182),
.B(n_1136),
.C(n_1202),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1204),
.B(n_1179),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1142),
.B(n_1156),
.Y(n_1304)
);

AOI221xp5_ASAP7_75t_L g1305 ( 
.A1(n_1117),
.A2(n_1157),
.B1(n_1248),
.B2(n_1244),
.C(n_1145),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1120),
.A2(n_1124),
.B(n_1172),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1217),
.B(n_1166),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1253),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1120),
.A2(n_1172),
.B(n_1181),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1187),
.A2(n_1178),
.B(n_1150),
.Y(n_1310)
);

CKINVDCx16_ASAP7_75t_R g1311 ( 
.A(n_1236),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1179),
.B(n_1174),
.Y(n_1312)
);

NAND2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1225),
.B(n_1196),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1173),
.B(n_1118),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1176),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_SL g1316 ( 
.A1(n_1190),
.A2(n_1173),
.B(n_1178),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1200),
.Y(n_1317)
);

AOI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1157),
.A2(n_1247),
.B1(n_1246),
.B2(n_1135),
.C(n_1121),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1132),
.A2(n_1188),
.B1(n_1203),
.B2(n_1174),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1130),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1132),
.A2(n_1203),
.B1(n_1174),
.B2(n_1135),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1129),
.B(n_1225),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1126),
.A2(n_1195),
.B(n_1183),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1170),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1125),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1185),
.A2(n_1231),
.B1(n_1195),
.B2(n_1123),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1189),
.A2(n_1119),
.B(n_1193),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1224),
.A2(n_1213),
.B1(n_1141),
.B2(n_1229),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1194),
.A2(n_1229),
.B(n_1232),
.Y(n_1329)
);

AO32x2_ASAP7_75t_L g1330 ( 
.A1(n_1141),
.A2(n_1232),
.A3(n_1233),
.B1(n_1240),
.B2(n_1213),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1141),
.B(n_1216),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1234),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1223),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1219),
.A2(n_897),
.B(n_903),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1207),
.B(n_1241),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1158),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1199),
.A2(n_1138),
.B1(n_970),
.B2(n_897),
.Y(n_1337)
);

AOI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1209),
.A2(n_510),
.B(n_534),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1197),
.A2(n_1205),
.B(n_1201),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1158),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1223),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1234),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1199),
.A2(n_1138),
.B1(n_986),
.B2(n_988),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1163),
.A2(n_970),
.B1(n_897),
.B2(n_1230),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1225),
.B(n_1009),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1219),
.A2(n_897),
.B(n_903),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1167),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1223),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1167),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1199),
.B(n_1138),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1206),
.B(n_1208),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1234),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1197),
.A2(n_1205),
.B(n_1201),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1158),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1184),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1209),
.A2(n_322),
.B1(n_331),
.B2(n_321),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1206),
.B(n_1208),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1184),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1184),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1250),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1214),
.A2(n_1222),
.B(n_1221),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1207),
.B(n_1241),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1151),
.A2(n_897),
.B1(n_1208),
.B2(n_1206),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1184),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1206),
.B(n_1208),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1165),
.B(n_1133),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1199),
.B(n_1138),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1216),
.B(n_1250),
.Y(n_1368)
);

AO32x2_ASAP7_75t_L g1369 ( 
.A1(n_1230),
.A2(n_1251),
.A3(n_988),
.B1(n_1020),
.B2(n_999),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1219),
.A2(n_897),
.B(n_903),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1263),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1269),
.B(n_1331),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1344),
.A2(n_1337),
.B1(n_1268),
.B2(n_1343),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1264),
.B(n_1266),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1301),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1265),
.B(n_1368),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1277),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1335),
.B(n_1362),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1269),
.B(n_1330),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1351),
.B(n_1357),
.Y(n_1380)
);

OA22x2_ASAP7_75t_L g1381 ( 
.A1(n_1350),
.A2(n_1367),
.B1(n_1289),
.B2(n_1299),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1301),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1304),
.B(n_1257),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1365),
.B(n_1283),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1336),
.B(n_1340),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1258),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1330),
.B(n_1261),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1277),
.Y(n_1388)
);

O2A1O1Ixp5_ASAP7_75t_L g1389 ( 
.A1(n_1343),
.A2(n_1272),
.B(n_1367),
.C(n_1350),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1270),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1312),
.B(n_1323),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1348),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1288),
.B(n_1295),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1354),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1330),
.B(n_1261),
.Y(n_1395)
);

OA22x2_ASAP7_75t_L g1396 ( 
.A1(n_1260),
.A2(n_1276),
.B1(n_1295),
.B2(n_1363),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1345),
.A2(n_1280),
.B(n_1305),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_SL g1398 ( 
.A1(n_1334),
.A2(n_1346),
.B(n_1370),
.C(n_1344),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1324),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1284),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1271),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1256),
.A2(n_1262),
.B(n_1300),
.C(n_1306),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1326),
.A2(n_1286),
.B1(n_1338),
.B2(n_1260),
.Y(n_1403)
);

AO21x1_ASAP7_75t_L g1404 ( 
.A1(n_1327),
.A2(n_1314),
.B(n_1325),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1260),
.A2(n_1356),
.B1(n_1307),
.B2(n_1360),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1312),
.B(n_1322),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1330),
.B(n_1261),
.Y(n_1407)
);

NOR2xp67_ASAP7_75t_R g1408 ( 
.A(n_1297),
.B(n_1259),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1341),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1341),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1348),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1319),
.B(n_1321),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1307),
.B(n_1318),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1328),
.A2(n_1333),
.B1(n_1274),
.B2(n_1296),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1319),
.B(n_1321),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1328),
.A2(n_1274),
.B1(n_1333),
.B2(n_1312),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1311),
.B(n_1302),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1285),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1275),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1316),
.A2(n_1281),
.B(n_1294),
.C(n_1308),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1320),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1273),
.B(n_1366),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1309),
.A2(n_1293),
.B(n_1329),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1287),
.A2(n_1310),
.B(n_1292),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1291),
.A2(n_1315),
.B1(n_1342),
.B2(n_1303),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1291),
.A2(n_1315),
.B1(n_1342),
.B2(n_1332),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1275),
.B(n_1361),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1369),
.B(n_1275),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1348),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1317),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1258),
.B(n_1352),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1332),
.B(n_1352),
.Y(n_1432)
);

AOI21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1313),
.A2(n_1369),
.B(n_1281),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1267),
.A2(n_1364),
.B(n_1359),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1317),
.B(n_1255),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1355),
.A2(n_1364),
.B(n_1359),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1355),
.A2(n_1358),
.B(n_1278),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1279),
.B(n_1282),
.Y(n_1438)
);

AOI211xp5_ASAP7_75t_L g1439 ( 
.A1(n_1347),
.A2(n_1349),
.B(n_1353),
.C(n_1339),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1279),
.B(n_1282),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1347),
.B(n_1297),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1338),
.A2(n_897),
.B(n_1146),
.C(n_438),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1342),
.Y(n_1443)
);

O2A1O1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1338),
.A2(n_897),
.B(n_1146),
.C(n_438),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1338),
.A2(n_897),
.B(n_1146),
.C(n_438),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1290),
.B(n_1298),
.Y(n_1446)
);

OA22x2_ASAP7_75t_L g1447 ( 
.A1(n_1350),
.A2(n_935),
.B1(n_1367),
.B2(n_1117),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1338),
.A2(n_897),
.B(n_1146),
.C(n_438),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1399),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1373),
.A2(n_1398),
.B1(n_1448),
.B2(n_1445),
.C(n_1444),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1447),
.A2(n_1413),
.B1(n_1403),
.B2(n_1405),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1447),
.A2(n_1396),
.B1(n_1381),
.B2(n_1374),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1427),
.B(n_1419),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1442),
.A2(n_1402),
.B(n_1380),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1401),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1418),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1379),
.B(n_1387),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1391),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1434),
.A2(n_1436),
.B(n_1437),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1391),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1395),
.B(n_1407),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1393),
.B(n_1372),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1395),
.B(n_1407),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1428),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1372),
.B(n_1412),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1415),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1412),
.A2(n_1415),
.B(n_1371),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1398),
.A2(n_1397),
.B(n_1440),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1390),
.A2(n_1440),
.B(n_1438),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1394),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1384),
.B(n_1376),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1391),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1423),
.B(n_1381),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1396),
.B(n_1424),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1397),
.B(n_1406),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1439),
.Y(n_1476)
);

OR2x6_ASAP7_75t_L g1477 ( 
.A(n_1406),
.B(n_1420),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1385),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1417),
.B(n_1446),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1383),
.B(n_1410),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1409),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1422),
.A2(n_1414),
.B(n_1416),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1462),
.B(n_1377),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1449),
.Y(n_1485)
);

NOR4xp25_ASAP7_75t_SL g1486 ( 
.A(n_1450),
.B(n_1375),
.C(n_1382),
.D(n_1386),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1469),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1476),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1451),
.B(n_1386),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1463),
.B(n_1378),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1477),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1388),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1469),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1460),
.B(n_1430),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1453),
.B(n_1400),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1497)
);

CKINVDCx14_ASAP7_75t_R g1498 ( 
.A(n_1479),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1470),
.B(n_1435),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1455),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1460),
.B(n_1458),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1451),
.A2(n_1443),
.B1(n_1392),
.B2(n_1411),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1457),
.B(n_1464),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1453),
.B(n_1467),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_SL g1505 ( 
.A(n_1459),
.B(n_1433),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1455),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1456),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1459),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1467),
.B(n_1425),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1492),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1490),
.A2(n_1450),
.B1(n_1452),
.B2(n_1454),
.C(n_1476),
.Y(n_1511)
);

OAI211xp5_ASAP7_75t_L g1512 ( 
.A1(n_1489),
.A2(n_1452),
.B(n_1466),
.C(n_1471),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1502),
.A2(n_1475),
.B1(n_1477),
.B2(n_1466),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1486),
.A2(n_1477),
.B1(n_1475),
.B2(n_1466),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1485),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1502),
.A2(n_1489),
.B1(n_1481),
.B2(n_1471),
.C(n_1483),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1488),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1485),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1508),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1501),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1505),
.A2(n_1466),
.B1(n_1498),
.B2(n_1468),
.Y(n_1522)
);

OR2x2_ASAP7_75t_SL g1523 ( 
.A(n_1509),
.B(n_1466),
.Y(n_1523)
);

OAI31xp33_ASAP7_75t_L g1524 ( 
.A1(n_1509),
.A2(n_1474),
.A3(n_1426),
.B(n_1473),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1492),
.A2(n_1477),
.B1(n_1466),
.B2(n_1475),
.C(n_1480),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1495),
.A2(n_1475),
.B1(n_1477),
.B2(n_1482),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1503),
.B(n_1457),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1495),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1492),
.A2(n_1475),
.B1(n_1477),
.B2(n_1482),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1483),
.A2(n_1481),
.B1(n_1478),
.B2(n_1480),
.C(n_1473),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

OAI31xp33_ASAP7_75t_L g1532 ( 
.A1(n_1496),
.A2(n_1479),
.A3(n_1429),
.B(n_1392),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1495),
.A2(n_1475),
.B1(n_1477),
.B2(n_1482),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1501),
.B(n_1472),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_1479),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1516),
.Y(n_1536)
);

INVx5_ASAP7_75t_L g1537 ( 
.A(n_1520),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1514),
.B(n_1487),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1521),
.B(n_1487),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1516),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1518),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1523),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1519),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1519),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1520),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1520),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1520),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1530),
.B(n_1500),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1531),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1528),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1537),
.B(n_1521),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1548),
.B(n_1535),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1542),
.B(n_1528),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1542),
.B(n_1528),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1536),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1536),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1542),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1548),
.A2(n_1511),
.B(n_1522),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1548),
.B(n_1497),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1552),
.B(n_1421),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1536),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1542),
.B(n_1517),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1552),
.B(n_1421),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1549),
.B(n_1491),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1540),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1549),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1497),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1551),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1537),
.B(n_1534),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1552),
.B(n_1443),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1540),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1543),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1551),
.B(n_1491),
.Y(n_1577)
);

INVx8_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1551),
.B(n_1524),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1539),
.B(n_1552),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1537),
.A2(n_1513),
.B1(n_1533),
.B2(n_1529),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1543),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1584)
);

OAI33xp33_ASAP7_75t_L g1585 ( 
.A1(n_1544),
.A2(n_1499),
.A3(n_1496),
.B1(n_1515),
.B2(n_1506),
.B3(n_1507),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1551),
.Y(n_1586)
);

AOI211x1_ASAP7_75t_L g1587 ( 
.A1(n_1538),
.A2(n_1525),
.B(n_1484),
.C(n_1493),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1526),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1544),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1544),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1578),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1559),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1573),
.B(n_1537),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1557),
.B(n_1537),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1562),
.B(n_1550),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1590),
.B(n_1551),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1578),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1562),
.B(n_1550),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1570),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1590),
.B(n_1538),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1564),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1564),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1567),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1572),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1586),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1560),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1567),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1589),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1561),
.B(n_1532),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_SL g1613 ( 
.A(n_1578),
.B(n_1537),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1565),
.B(n_1541),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1589),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1538),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1584),
.B(n_1547),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1558),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1569),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1575),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1576),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1582),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1583),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1591),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1571),
.B(n_1550),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1554),
.B(n_1550),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1597),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1607),
.B(n_1563),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1609),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1597),
.B(n_1555),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1555),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1595),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1600),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1601),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1600),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1617),
.B(n_1573),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1604),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1604),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1594),
.B(n_1573),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1595),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1614),
.B(n_1618),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1612),
.B(n_1566),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1614),
.B(n_1618),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1604),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1593),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1595),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1593),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1606),
.B(n_1587),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1594),
.B(n_1556),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1652),
.A2(n_1646),
.B(n_1630),
.C(n_1639),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1628),
.B(n_1606),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1629),
.A2(n_1579),
.B(n_1613),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1645),
.A2(n_1613),
.B(n_1581),
.Y(n_1657)
);

O2A1O1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1635),
.A2(n_1645),
.B(n_1647),
.C(n_1608),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1633),
.Y(n_1659)
);

OAI211xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1647),
.A2(n_1592),
.B(n_1598),
.C(n_1608),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1653),
.B(n_1592),
.Y(n_1661)
);

AOI211x1_ASAP7_75t_SL g1662 ( 
.A1(n_1634),
.A2(n_1650),
.B(n_1644),
.C(n_1627),
.Y(n_1662)
);

OAI222xp33_ASAP7_75t_L g1663 ( 
.A1(n_1628),
.A2(n_1598),
.B1(n_1556),
.B2(n_1627),
.C1(n_1596),
.C2(n_1599),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1635),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1633),
.B(n_1616),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1631),
.B(n_1632),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

AOI32xp33_ASAP7_75t_L g1668 ( 
.A1(n_1631),
.A2(n_1580),
.A3(n_1594),
.B1(n_1616),
.B2(n_1602),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1640),
.A2(n_1588),
.B1(n_1537),
.B2(n_1577),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1632),
.B(n_1620),
.C(n_1619),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1649),
.A2(n_1578),
.B(n_1585),
.Y(n_1671)
);

NAND2x1_ASAP7_75t_L g1672 ( 
.A(n_1640),
.B(n_1594),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1636),
.Y(n_1673)
);

BUFx12f_ASAP7_75t_L g1674 ( 
.A(n_1665),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1664),
.B(n_1653),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1659),
.B(n_1640),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1640),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1656),
.B(n_1653),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1672),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1666),
.B(n_1653),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1655),
.B(n_1596),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1658),
.A2(n_1486),
.B1(n_1651),
.B2(n_1649),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1667),
.B(n_1658),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1643),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1668),
.B(n_1660),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1674),
.A2(n_1671),
.B1(n_1643),
.B2(n_1670),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1676),
.B(n_1654),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_L g1688 ( 
.A1(n_1683),
.A2(n_1671),
.B(n_1662),
.C(n_1673),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1681),
.B(n_1663),
.Y(n_1689)
);

OAI211xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1682),
.A2(n_1634),
.B(n_1644),
.C(n_1650),
.Y(n_1690)
);

OA211x2_ASAP7_75t_L g1691 ( 
.A1(n_1675),
.A2(n_1432),
.B(n_1431),
.C(n_1568),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1682),
.A2(n_1678),
.B(n_1675),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1679),
.A2(n_1677),
.B1(n_1680),
.B2(n_1669),
.C(n_1599),
.Y(n_1693)
);

AOI222xp33_ASAP7_75t_L g1694 ( 
.A1(n_1679),
.A2(n_1651),
.B1(n_1643),
.B2(n_1641),
.C1(n_1638),
.C2(n_1648),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1694),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1685),
.A2(n_1643),
.B(n_1637),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1687),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1686),
.A2(n_1626),
.B1(n_1546),
.B2(n_1545),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1688),
.A2(n_1537),
.B1(n_1547),
.B2(n_1553),
.Y(n_1699)
);

OAI322xp33_ASAP7_75t_L g1700 ( 
.A1(n_1689),
.A2(n_1648),
.A3(n_1642),
.B1(n_1641),
.B2(n_1638),
.C1(n_1637),
.C2(n_1636),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1692),
.A2(n_1642),
.B(n_1620),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_R g1702 ( 
.A(n_1695),
.B(n_1697),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1696),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1699),
.B(n_1690),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1698),
.B(n_1602),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1701),
.B(n_1693),
.C(n_1622),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1700),
.B(n_1580),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1703),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_SL g1709 ( 
.A1(n_1707),
.A2(n_1621),
.B(n_1623),
.C(n_1625),
.Y(n_1709)
);

NAND4xp75_ASAP7_75t_L g1710 ( 
.A(n_1704),
.B(n_1691),
.C(n_1615),
.D(n_1611),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1706),
.B(n_1619),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1705),
.A2(n_1621),
.B1(n_1623),
.B2(n_1625),
.Y(n_1712)
);

AOI222xp33_ASAP7_75t_L g1713 ( 
.A1(n_1709),
.A2(n_1702),
.B1(n_1622),
.B2(n_1624),
.C1(n_1603),
.C2(n_1610),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1711),
.B(n_1702),
.C(n_1411),
.Y(n_1714)
);

NAND4xp75_ASAP7_75t_L g1715 ( 
.A(n_1708),
.B(n_1605),
.C(n_1603),
.D(n_1610),
.Y(n_1715)
);

AND2x2_ASAP7_75t_SL g1716 ( 
.A(n_1714),
.B(n_1712),
.Y(n_1716)
);

AOI322xp5_ASAP7_75t_L g1717 ( 
.A1(n_1716),
.A2(n_1710),
.A3(n_1715),
.B1(n_1713),
.B2(n_1605),
.C1(n_1611),
.C2(n_1615),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1621),
.B1(n_1625),
.B2(n_1623),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1717),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1719),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1718),
.Y(n_1721)
);

AO22x2_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1624),
.B1(n_1626),
.B2(n_1553),
.Y(n_1722)
);

INVxp67_ASAP7_75t_SL g1723 ( 
.A(n_1721),
.Y(n_1723)
);

XNOR2xp5_ASAP7_75t_L g1724 ( 
.A(n_1723),
.B(n_1441),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1722),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1725),
.A2(n_1553),
.B1(n_1547),
.B2(n_1546),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1724),
.B(n_1408),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1727),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1546),
.B1(n_1545),
.B2(n_1547),
.Y(n_1729)
);

AOI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1441),
.B(n_1546),
.C(n_1545),
.Y(n_1730)
);


endmodule