module fake_jpeg_25910_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_6),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_6),
.A2(n_5),
.B1(n_2),
.B2(n_4),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_13),
.A2(n_0),
.B1(n_14),
.B2(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.C(n_8),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_21),
.C(n_15),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_10),
.B(n_8),
.C(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_9),
.B(n_8),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.C(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_25),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_21),
.Y(n_32)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_33),
.CI(n_35),
.CON(n_38),
.SN(n_38)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_24),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_23),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_23),
.A3(n_32),
.B1(n_35),
.B2(n_38),
.C1(n_39),
.C2(n_34),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_43),
.B(n_38),
.C(n_42),
.Y(n_45)
);


endmodule