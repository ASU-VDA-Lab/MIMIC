module fake_jpeg_2733_n_661 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_661);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_661;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_10),
.B(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_62),
.B(n_124),
.Y(n_170)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_63),
.Y(n_200)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_64),
.Y(n_132)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_68),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_71),
.Y(n_194)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_80),
.Y(n_142)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_74),
.Y(n_179)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_79),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_8),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_84),
.Y(n_186)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_31),
.B(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_89),
.B(n_92),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_10),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_95),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_21),
.Y(n_96)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_10),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_108),
.B(n_110),
.Y(n_208)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_32),
.B(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_111),
.B(n_122),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_21),
.Y(n_113)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_32),
.B(n_12),
.Y(n_122)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_34),
.Y(n_131)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_53),
.B1(n_34),
.B2(n_48),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_138),
.A2(n_162),
.B1(n_165),
.B2(n_185),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_60),
.B(n_52),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_140),
.B(n_144),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_77),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_143),
.A2(n_88),
.B1(n_97),
.B2(n_95),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_68),
.B(n_52),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_41),
.C(n_45),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_157),
.B(n_173),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_113),
.A2(n_34),
.B1(n_48),
.B2(n_45),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_61),
.A2(n_34),
.B1(n_48),
.B2(n_24),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_107),
.B(n_48),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_81),
.B(n_38),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_177),
.B(n_182),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_55),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_99),
.A2(n_24),
.B1(n_37),
.B2(n_47),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_184),
.A2(n_169),
.A3(n_164),
.B1(n_152),
.B2(n_156),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_82),
.A2(n_37),
.B1(n_49),
.B2(n_47),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_109),
.B(n_55),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_188),
.B(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_202),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_43),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_215),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_82),
.A2(n_43),
.B1(n_42),
.B2(n_38),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_206),
.A2(n_207),
.B1(n_159),
.B2(n_178),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_64),
.A2(n_42),
.B1(n_116),
.B2(n_103),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_101),
.B(n_12),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_102),
.A2(n_6),
.B1(n_18),
.B2(n_2),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_212),
.A2(n_138),
.B1(n_207),
.B2(n_162),
.Y(n_260)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_59),
.Y(n_214)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_214),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_105),
.B(n_19),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_66),
.Y(n_216)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_216),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_64),
.A2(n_6),
.B(n_18),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_15),
.B(n_19),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_220),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_70),
.B(n_6),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_223),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_71),
.B(n_6),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_76),
.B(n_19),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_0),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_159),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_229),
.B(n_256),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

INVx8_ASAP7_75t_L g369 ( 
.A(n_230),
.Y(n_369)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_231),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_234),
.A2(n_260),
.B1(n_181),
.B2(n_199),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_235),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_151),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_236),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_132),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_238),
.Y(n_354)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_239),
.Y(n_364)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_240),
.Y(n_352)
);

INVx3_ASAP7_75t_SL g241 ( 
.A(n_200),
.Y(n_241)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_241),
.Y(n_361)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_244),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_SL g314 ( 
.A1(n_246),
.A2(n_270),
.B(n_302),
.C(n_172),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_247),
.A2(n_172),
.B(n_192),
.Y(n_329)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_189),
.A2(n_98),
.B1(n_90),
.B2(n_86),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_249),
.A2(n_277),
.B1(n_288),
.B2(n_294),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_251),
.B(n_267),
.Y(n_323)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_139),
.Y(n_253)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_254),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_179),
.Y(n_255)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_255),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_178),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_257),
.Y(n_353)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_158),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_259),
.Y(n_366)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_261),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_262),
.Y(n_358)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_137),
.Y(n_264)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_264),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_170),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_265),
.B(n_276),
.Y(n_359)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_158),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_266),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_160),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_196),
.A2(n_13),
.B(n_19),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_268),
.B(n_274),
.Y(n_332)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_269),
.Y(n_363)
);

AOI211xp5_ASAP7_75t_SL g270 ( 
.A1(n_184),
.A2(n_84),
.B(n_79),
.C(n_2),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_206),
.A2(n_4),
.B1(n_15),
.B2(n_2),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_271),
.A2(n_194),
.B1(n_155),
.B2(n_175),
.Y(n_326)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_272),
.Y(n_367)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_273),
.Y(n_372)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_279),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_201),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_219),
.A2(n_179),
.B1(n_180),
.B2(n_200),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_184),
.A2(n_5),
.B1(n_15),
.B2(n_3),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_278),
.A2(n_307),
.B1(n_135),
.B2(n_161),
.Y(n_313)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_171),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_280),
.B(n_281),
.Y(n_368)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_150),
.B(n_4),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_282),
.B(n_285),
.Y(n_339)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_187),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_295),
.Y(n_315)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_284),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_208),
.B(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_225),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_286),
.A2(n_146),
.B1(n_191),
.B2(n_199),
.Y(n_321)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_134),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_287),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_147),
.A2(n_14),
.B1(n_16),
.B2(n_0),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_134),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_289),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_142),
.B(n_0),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_291),
.B(n_296),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_173),
.B(n_145),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_238),
.C(n_235),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_293),
.Y(n_350)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_136),
.B(n_1),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_141),
.B(n_1),
.Y(n_296)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_165),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_297),
.Y(n_371)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_166),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_167),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_300),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_228),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_133),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_306),
.Y(n_319)
);

CKINVDCx6p67_ASAP7_75t_R g302 ( 
.A(n_185),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_228),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_305),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_221),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_204),
.A2(n_1),
.B1(n_135),
.B2(n_161),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_190),
.B(n_193),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_310),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_181),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_269),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_313),
.A2(n_314),
.B1(n_338),
.B2(n_241),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_316),
.A2(n_326),
.B1(n_355),
.B2(n_255),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_330),
.B1(n_348),
.B2(n_365),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_191),
.C(n_194),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_289),
.C(n_287),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_329),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_302),
.A2(n_175),
.B1(n_176),
.B2(n_205),
.Y(n_330)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_176),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_336),
.B(n_342),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_302),
.A2(n_205),
.B1(n_155),
.B2(n_192),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_258),
.B(n_245),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_245),
.B(n_263),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_346),
.B(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_250),
.B(n_310),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_302),
.A2(n_234),
.B1(n_270),
.B2(n_292),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_243),
.A2(n_292),
.B1(n_247),
.B2(n_233),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_255),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_297),
.A2(n_286),
.B1(n_283),
.B2(n_264),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_341),
.B(n_308),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_375),
.B(n_376),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_339),
.B(n_248),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_359),
.B(n_237),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_377),
.B(n_383),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_390),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_356),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_392),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_381),
.A2(n_393),
.B1(n_371),
.B2(n_314),
.Y(n_422)
);

AO21x2_ASAP7_75t_L g382 ( 
.A1(n_329),
.A2(n_242),
.B(n_254),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_382),
.A2(n_385),
.B1(n_386),
.B2(n_388),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_315),
.B(n_232),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_361),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_348),
.A2(n_290),
.B1(n_312),
.B2(n_303),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_365),
.A2(n_252),
.B1(n_261),
.B2(n_298),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_322),
.A2(n_266),
.B1(n_259),
.B2(n_239),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_387),
.A2(n_316),
.B1(n_321),
.B2(n_335),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_322),
.A2(n_252),
.B1(n_284),
.B2(n_244),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_346),
.B(n_240),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_299),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_417),
.C(n_367),
.Y(n_449)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_315),
.B(n_274),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_407),
.Y(n_424)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_328),
.Y(n_403)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_403),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_328),
.Y(n_405)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_405),
.Y(n_456)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_336),
.B(n_281),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_409),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_318),
.Y(n_409)
);

AO21x2_ASAP7_75t_L g410 ( 
.A1(n_330),
.A2(n_273),
.B(n_253),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_415),
.B1(n_257),
.B2(n_333),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_411),
.Y(n_430)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_413),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_414),
.Y(n_454)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_314),
.A2(n_347),
.B1(n_371),
.B2(n_324),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_332),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_418),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_342),
.B(n_293),
.C(n_279),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_319),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_421),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_355),
.A2(n_267),
.B(n_251),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_420),
.A2(n_344),
.B(n_320),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_422),
.A2(n_427),
.B1(n_382),
.B2(n_393),
.Y(n_477)
);

FAx1_ASAP7_75t_SL g423 ( 
.A(n_397),
.B(n_360),
.CI(n_314),
.CON(n_423),
.SN(n_423)
);

OAI32xp33_ASAP7_75t_L g467 ( 
.A1(n_423),
.A2(n_378),
.A3(n_396),
.B1(n_415),
.B2(n_417),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_399),
.A2(n_314),
.B1(n_318),
.B2(n_370),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_428),
.A2(n_431),
.B1(n_438),
.B2(n_444),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_370),
.Y(n_429)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_380),
.A2(n_327),
.B1(n_350),
.B2(n_343),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_343),
.Y(n_432)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_374),
.A2(n_420),
.B(n_382),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_437),
.A2(n_441),
.B(n_447),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_380),
.A2(n_350),
.B1(n_334),
.B2(n_337),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_382),
.A2(n_334),
.B(n_354),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_397),
.A2(n_354),
.B(n_344),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_407),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_325),
.C(n_353),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_450),
.B(n_457),
.C(n_395),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_395),
.B(n_325),
.C(n_353),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_418),
.B(n_333),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_459),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_415),
.A2(n_236),
.B1(n_364),
.B2(n_373),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_387),
.B1(n_410),
.B2(n_382),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_442),
.B(n_396),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_463),
.B(n_453),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_464),
.B(n_467),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_469),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_435),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_470),
.B(n_472),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_392),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_471),
.B(n_478),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_434),
.B(n_389),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_474),
.B(n_475),
.C(n_480),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_449),
.C(n_450),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_477),
.A2(n_459),
.B1(n_430),
.B2(n_436),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_413),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_479),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_388),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_452),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_481),
.B(n_491),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_489),
.B1(n_428),
.B2(n_433),
.Y(n_508)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_484),
.Y(n_522)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_425),
.Y(n_485)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_404),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_486),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_394),
.C(n_385),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_493),
.C(n_440),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_406),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_488),
.B(n_496),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_460),
.A2(n_386),
.B1(n_410),
.B2(n_398),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_497),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_432),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_437),
.B(n_419),
.C(n_411),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_434),
.B(n_340),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_494),
.B(n_499),
.Y(n_534)
);

XOR2x2_ASAP7_75t_L g496 ( 
.A(n_423),
.B(n_372),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_461),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_461),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_500),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_453),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_501),
.B(n_511),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_441),
.B(n_462),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_504),
.A2(n_506),
.B(n_509),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_427),
.B(n_444),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_508),
.A2(n_513),
.B1(n_524),
.B2(n_483),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_424),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_473),
.A2(n_423),
.B1(n_424),
.B2(n_459),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_423),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_514),
.B(n_518),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_477),
.A2(n_431),
.B1(n_438),
.B2(n_433),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_515),
.A2(n_517),
.B1(n_519),
.B2(n_521),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_445),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_516),
.B(n_500),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_473),
.A2(n_452),
.B1(n_436),
.B2(n_426),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_463),
.B(n_459),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_443),
.Y(n_520)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_520),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_482),
.A2(n_445),
.B1(n_451),
.B2(n_446),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_466),
.A2(n_410),
.B1(n_456),
.B2(n_451),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_479),
.B(n_443),
.Y(n_525)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_525),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_493),
.B(n_440),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_476),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_489),
.A2(n_468),
.B1(n_466),
.B2(n_465),
.Y(n_528)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_528),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_468),
.A2(n_456),
.B1(n_446),
.B2(n_454),
.Y(n_529)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_529),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_464),
.C(n_480),
.Y(n_539)
);

XNOR2x1_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_496),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_537),
.B(n_520),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_539),
.B(n_548),
.C(n_561),
.Y(n_570)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_541),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_545),
.A2(n_552),
.B1(n_554),
.B2(n_560),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_495),
.C(n_465),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_515),
.A2(n_485),
.B1(n_495),
.B2(n_467),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_549),
.A2(n_555),
.B1(n_556),
.B2(n_503),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_557),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_506),
.A2(n_498),
.B1(n_497),
.B2(n_490),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_384),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_533),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_513),
.A2(n_410),
.B1(n_430),
.B2(n_454),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_517),
.A2(n_469),
.B1(n_414),
.B2(n_412),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_519),
.A2(n_504),
.B1(n_535),
.B2(n_505),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_525),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_530),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_559),
.Y(n_585)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_507),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_505),
.A2(n_535),
.B1(n_527),
.B2(n_524),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_526),
.B(n_272),
.C(n_262),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_562),
.Y(n_580)
);

CKINVDCx14_ASAP7_75t_R g587 ( 
.A(n_563),
.Y(n_587)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_509),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_523),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_SL g565 ( 
.A1(n_527),
.A2(n_358),
.B(n_372),
.C(n_363),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g572 ( 
.A1(n_565),
.A2(n_502),
.B(n_531),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_526),
.B(n_514),
.C(n_533),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_566),
.B(n_512),
.C(n_534),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_567),
.B(n_540),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_501),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_568),
.B(n_569),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_548),
.B(n_518),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_571),
.B(n_567),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_572),
.A2(n_560),
.B(n_565),
.Y(n_603)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_573),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_574),
.B(n_537),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_539),
.B(n_502),
.C(n_522),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_578),
.Y(n_597)
);

AOI21xp33_ASAP7_75t_L g577 ( 
.A1(n_563),
.A2(n_510),
.B(n_522),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_577),
.A2(n_543),
.B(n_565),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_541),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_545),
.A2(n_503),
.B1(n_408),
.B2(n_345),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_581),
.B(n_555),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_582),
.A2(n_586),
.B1(n_554),
.B2(n_552),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_358),
.C(n_352),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_584),
.B(n_589),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_544),
.A2(n_373),
.B1(n_366),
.B2(n_280),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_352),
.C(n_340),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_546),
.B(n_357),
.C(n_363),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_590),
.B(n_568),
.C(n_540),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_587),
.A2(n_556),
.B(n_549),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_591),
.A2(n_603),
.B(n_331),
.Y(n_624)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_592),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_598),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_595),
.B(n_601),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_574),
.B(n_575),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_596),
.B(n_600),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_576),
.A2(n_547),
.B1(n_538),
.B2(n_551),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_599),
.A2(n_582),
.B1(n_580),
.B2(n_579),
.Y(n_621)
);

AOI21x1_ASAP7_75t_L g623 ( 
.A1(n_604),
.A2(n_609),
.B(n_584),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_543),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_605),
.B(n_606),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_585),
.B(n_546),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_571),
.B(n_565),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_608),
.B(n_610),
.Y(n_613)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_572),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_366),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_596),
.B(n_589),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_615),
.B(n_618),
.Y(n_627)
);

INVx11_ASAP7_75t_L g616 ( 
.A(n_597),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_616),
.A2(n_594),
.B1(n_369),
.B2(n_306),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_610),
.B(n_570),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_590),
.C(n_569),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_625),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_621),
.A2(n_622),
.B1(n_230),
.B2(n_624),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_599),
.A2(n_586),
.B1(n_588),
.B2(n_572),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_623),
.B(n_608),
.Y(n_632)
);

OAI21xp33_ASAP7_75t_L g630 ( 
.A1(n_624),
.A2(n_592),
.B(n_603),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_593),
.B(n_357),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_591),
.A2(n_331),
.B(n_301),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_626),
.A2(n_595),
.B(n_598),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_612),
.B(n_602),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_630),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_600),
.C(n_593),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_631),
.B(n_635),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_632),
.B(n_633),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_634),
.A2(n_636),
.B1(n_638),
.B2(n_621),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_612),
.B(n_305),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_614),
.A2(n_231),
.B(n_294),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_615),
.B(n_230),
.C(n_620),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_637),
.B(n_611),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_627),
.B(n_619),
.Y(n_640)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_640),
.B(n_641),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_SL g641 ( 
.A(n_632),
.B(n_611),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_642),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_644),
.A2(n_645),
.B(n_647),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_631),
.B(n_617),
.C(n_613),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_629),
.B(n_616),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_639),
.A2(n_638),
.B(n_630),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_648),
.B(n_652),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_643),
.A2(n_637),
.B(n_622),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_650),
.B(n_645),
.Y(n_653)
);

AO21x1_ASAP7_75t_L g657 ( 
.A1(n_653),
.A2(n_654),
.B(n_651),
.Y(n_657)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_649),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_655),
.B(n_641),
.Y(n_656)
);

AO21x2_ASAP7_75t_L g658 ( 
.A1(n_656),
.A2(n_657),
.B(n_646),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_646),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_613),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_660),
.B(n_625),
.Y(n_661)
);


endmodule