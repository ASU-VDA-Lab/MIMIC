module fake_jpeg_8821_n_52 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_44;
wire n_28;
wire n_38;
wire n_24;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_15;

INVx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_8),
.B1(n_2),
.B2(n_5),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_34),
.B(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_35),
.B1(n_36),
.B2(n_21),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_31),
.C(n_37),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_42),
.Y(n_46)
);

AO221x1_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_20),
.B1(n_32),
.B2(n_35),
.C(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_29),
.Y(n_47)
);

AOI21x1_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_32),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

AOI31xp33_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_22),
.A3(n_17),
.B(n_19),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_48),
.A3(n_17),
.B1(n_19),
.B2(n_24),
.C1(n_26),
.C2(n_16),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_24),
.Y(n_52)
);


endmodule