module fake_jpeg_14366_n_640 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_640);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_640;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_60),
.B(n_61),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_69),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_25),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_81),
.Y(n_156)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_82),
.B(n_86),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_83),
.B(n_121),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_0),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_103),
.B(n_106),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_19),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_25),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_114),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_19),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_120),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_58),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_36),
.B(n_1),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_58),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_124),
.Y(n_135)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_29),
.B(n_32),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_125),
.B(n_53),
.Y(n_215)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_21),
.Y(n_127)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_39),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_39),
.Y(n_134)
);

INVx2_ASAP7_75t_R g129 ( 
.A(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_165),
.Y(n_221)
);

NAND2x1_ASAP7_75t_L g245 ( 
.A(n_134),
.B(n_46),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_76),
.A2(n_46),
.B1(n_35),
.B2(n_21),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_136),
.A2(n_211),
.B(n_41),
.Y(n_224)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_187),
.Y(n_218)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_117),
.Y(n_154)
);

BUFx4f_ASAP7_75t_SL g240 ( 
.A(n_154),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_163),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_30),
.Y(n_165)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_169),
.Y(n_283)
);

BUFx4f_ASAP7_75t_SL g171 ( 
.A(n_118),
.Y(n_171)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_87),
.Y(n_180)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_82),
.B(n_41),
.Y(n_187)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_119),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_30),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_144),
.Y(n_226)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_65),
.Y(n_193)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_59),
.Y(n_197)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_198),
.Y(n_279)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_64),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_127),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_208),
.Y(n_252)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_68),
.Y(n_203)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_66),
.Y(n_205)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_118),
.B(n_78),
.Y(n_206)
);

OR2x2_ASAP7_75t_SL g274 ( 
.A(n_206),
.B(n_212),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_75),
.A2(n_88),
.B1(n_84),
.B2(n_111),
.Y(n_211)
);

AND2x4_ASAP7_75t_SL g212 ( 
.A(n_92),
.B(n_46),
.Y(n_212)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_89),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_111),
.Y(n_255)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_223),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_224),
.A2(n_276),
.B1(n_286),
.B2(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_226),
.B(n_273),
.Y(n_313)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

CKINVDCx9p33_ASAP7_75t_R g231 ( 
.A(n_171),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_231),
.Y(n_352)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_151),
.Y(n_236)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_236),
.Y(n_351)
);

INVx6_ASAP7_75t_SL g237 ( 
.A(n_139),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_237),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_188),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_243),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_144),
.B(n_44),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_244),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_245),
.B(n_289),
.Y(n_315)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_166),
.A2(n_99),
.B1(n_77),
.B2(n_109),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_247),
.A2(n_253),
.B1(n_263),
.B2(n_145),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_133),
.Y(n_248)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_149),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_149),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_251),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_166),
.A2(n_116),
.B1(n_105),
.B2(n_102),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_140),
.Y(n_254)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_254),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_255),
.B(n_256),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_135),
.B(n_113),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_156),
.B(n_33),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_260),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_212),
.A2(n_98),
.B1(n_91),
.B2(n_73),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_258),
.A2(n_261),
.B1(n_56),
.B2(n_50),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_156),
.B(n_32),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_181),
.A2(n_69),
.B1(n_21),
.B2(n_35),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_131),
.B(n_31),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_262),
.B(n_266),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_189),
.A2(n_35),
.B1(n_56),
.B2(n_50),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_167),
.Y(n_265)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_265),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_131),
.B(n_129),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_153),
.Y(n_267)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_188),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_272),
.Y(n_339)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_269),
.Y(n_338)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_138),
.Y(n_271)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_185),
.B(n_113),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_29),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_277),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_160),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_176),
.B(n_31),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_162),
.B(n_33),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_284),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_134),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_162),
.B(n_40),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_290),
.Y(n_308)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_177),
.Y(n_286)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_196),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_217),
.B(n_53),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_245),
.C(n_206),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_217),
.B(n_44),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_184),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_187),
.B(n_43),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_293),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_143),
.B(n_40),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_292),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_146),
.B(n_43),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_274),
.B1(n_253),
.B2(n_247),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_294),
.A2(n_306),
.B1(n_312),
.B2(n_333),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_297),
.B(n_242),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_181),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_309),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_147),
.B1(n_145),
.B2(n_182),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_168),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_218),
.B(n_211),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_317),
.C(n_283),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_222),
.B(n_172),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_311),
.B(n_314),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_224),
.A2(n_164),
.B1(n_193),
.B2(n_203),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_232),
.B(n_210),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_139),
.C(n_136),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_271),
.A2(n_170),
.B1(n_142),
.B2(n_175),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_219),
.B(n_209),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_324),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_322),
.A2(n_328),
.B1(n_329),
.B2(n_341),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g324 ( 
.A1(n_225),
.A2(n_178),
.B1(n_202),
.B2(n_147),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_263),
.A2(n_182),
.B1(n_183),
.B2(n_196),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_261),
.A2(n_183),
.B1(n_201),
.B2(n_164),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_265),
.A2(n_204),
.B1(n_201),
.B2(n_174),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_237),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_240),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_259),
.B(n_204),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_337),
.B(n_340),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_220),
.B(n_173),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_163),
.B(n_186),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_345),
.Y(n_381)
);

AO22x1_ASAP7_75t_L g347 ( 
.A1(n_231),
.A2(n_163),
.B1(n_158),
.B2(n_132),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_347),
.B(n_324),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_290),
.A2(n_194),
.B1(n_155),
.B2(n_174),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_348),
.A2(n_227),
.B1(n_230),
.B2(n_104),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_319),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_354),
.B(n_365),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_355),
.B(n_356),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_296),
.B(n_221),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_294),
.A2(n_287),
.B1(n_286),
.B2(n_235),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_363),
.A2(n_367),
.B1(n_384),
.B2(n_352),
.Y(n_414)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_334),
.Y(n_364)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_240),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_316),
.A2(n_225),
.B1(n_228),
.B2(n_254),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_380),
.C(n_342),
.Y(n_430)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_323),
.B(n_234),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_398),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_314),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_378),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_238),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_372),
.B(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_310),
.B(n_141),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_387),
.B(n_345),
.Y(n_402)
);

INVx11_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_240),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_341),
.A2(n_304),
.B1(n_317),
.B2(n_297),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_379),
.A2(n_383),
.B1(n_306),
.B2(n_321),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_298),
.A2(n_282),
.B1(n_246),
.B2(n_236),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_382),
.A2(n_390),
.B1(n_396),
.B2(n_318),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_308),
.A2(n_228),
.B1(n_276),
.B2(n_250),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_315),
.A2(n_270),
.B1(n_223),
.B2(n_282),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_279),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_391),
.Y(n_428)
);

OR2x2_ASAP7_75t_SL g387 ( 
.A(n_344),
.B(n_242),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_305),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_388),
.Y(n_420)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_315),
.B(n_154),
.Y(n_391)
);

INVx13_ASAP7_75t_L g392 ( 
.A(n_298),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_392),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_241),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_311),
.B(n_309),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_346),
.Y(n_429)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_302),
.Y(n_396)
);

XNOR2x2_ASAP7_75t_SL g397 ( 
.A(n_325),
.B(n_299),
.Y(n_397)
);

XOR2x2_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_308),
.Y(n_399)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_326),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_400),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_308),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_402),
.A2(n_416),
.B(n_374),
.Y(n_450)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_407),
.A2(n_427),
.B1(n_373),
.B2(n_386),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_331),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_425),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

O2A1O1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_376),
.A2(n_347),
.B(n_324),
.C(n_343),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_359),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_375),
.A2(n_323),
.B(n_344),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_366),
.A2(n_324),
.B1(n_332),
.B2(n_330),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_417),
.A2(n_418),
.B1(n_432),
.B2(n_362),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_366),
.A2(n_327),
.B1(n_305),
.B2(n_303),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_361),
.B(n_301),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_423),
.B(n_386),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_343),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_342),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_431),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_379),
.A2(n_333),
.B1(n_248),
.B2(n_327),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_429),
.B(n_393),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_430),
.A2(n_374),
.B(n_354),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_351),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_363),
.A2(n_303),
.B1(n_349),
.B2(n_351),
.Y(n_432)
);

OAI32xp33_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_349),
.A3(n_295),
.B1(n_52),
.B2(n_53),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_383),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_372),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_360),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_437),
.B(n_431),
.C(n_408),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_404),
.A2(n_381),
.B1(n_395),
.B2(n_367),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_439),
.A2(n_462),
.B(n_410),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_442),
.A2(n_450),
.B(n_453),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_425),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_452),
.Y(n_489)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_445),
.A2(n_457),
.B1(n_459),
.B2(n_465),
.Y(n_490)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_422),
.Y(n_446)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_447),
.Y(n_491)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_448),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_449),
.B(n_460),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_423),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_454),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_357),
.Y(n_455)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_455),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_353),
.Y(n_456)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_404),
.A2(n_381),
.B(n_395),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_407),
.A2(n_362),
.B1(n_391),
.B2(n_353),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_356),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_466),
.B1(n_413),
.B2(n_405),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_402),
.A2(n_387),
.B(n_318),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_413),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_463),
.B(n_464),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_423),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_427),
.A2(n_396),
.B1(n_390),
.B2(n_364),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_417),
.A2(n_397),
.B1(n_369),
.B2(n_358),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_409),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_467),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_398),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_468),
.Y(n_498)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_401),
.Y(n_469)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_405),
.B(n_433),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_471),
.B(n_419),
.Y(n_473)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_474),
.A2(n_496),
.B(n_463),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_400),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_476),
.B(n_477),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_440),
.B(n_430),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_462),
.A2(n_439),
.B(n_410),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_479),
.B(n_495),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_483),
.A2(n_451),
.B1(n_442),
.B2(n_464),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_440),
.B(n_426),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_435),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_459),
.A2(n_414),
.B1(n_418),
.B2(n_428),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_486),
.A2(n_503),
.B1(n_451),
.B2(n_445),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_412),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_492),
.B(n_497),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_441),
.C(n_450),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_468),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_458),
.B(n_413),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_SL g497 ( 
.A(n_438),
.B(n_416),
.C(n_412),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_454),
.B(n_399),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_499),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_460),
.B(n_399),
.Y(n_500)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_500),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_433),
.Y(n_501)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_501),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_457),
.A2(n_432),
.B1(n_421),
.B2(n_415),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_489),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_506),
.B(n_514),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_451),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_507),
.A2(n_522),
.B(n_496),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_508),
.A2(n_516),
.B1(n_498),
.B2(n_472),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_509),
.B(n_491),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_441),
.C(n_438),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_511),
.C(n_513),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_455),
.C(n_471),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_443),
.C(n_456),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_420),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_515),
.A2(n_517),
.B1(n_503),
.B2(n_486),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_490),
.A2(n_453),
.B1(n_461),
.B2(n_452),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_483),
.A2(n_465),
.B1(n_453),
.B2(n_449),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_475),
.B(n_448),
.Y(n_519)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_519),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_397),
.C(n_453),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_521),
.C(n_524),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_420),
.C(n_421),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_444),
.C(n_447),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_528),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_488),
.B(n_424),
.Y(n_527)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_527),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_446),
.Y(n_528)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_534),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_401),
.C(n_295),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_485),
.C(n_481),
.Y(n_539)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_504),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_539),
.B(n_542),
.C(n_551),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_519),
.B(n_498),
.Y(n_540)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_541),
.A2(n_507),
.B1(n_525),
.B2(n_521),
.Y(n_562)
);

XNOR2x1_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_513),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_522),
.A2(n_472),
.B(n_479),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_544),
.A2(n_526),
.B(n_520),
.Y(n_563)
);

AO21x1_ASAP7_75t_L g565 ( 
.A1(n_545),
.A2(n_546),
.B(n_470),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_507),
.A2(n_482),
.B(n_474),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_529),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_389),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_549),
.A2(n_392),
.B1(n_56),
.B2(n_52),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_517),
.A2(n_502),
.B1(n_480),
.B2(n_488),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_550),
.A2(n_559),
.B1(n_516),
.B2(n_523),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_502),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_509),
.B(n_485),
.C(n_487),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_556),
.C(n_558),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_518),
.A2(n_530),
.B1(n_508),
.B2(n_531),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_550),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_512),
.B(n_424),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_555),
.B(n_547),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_505),
.B(n_491),
.C(n_487),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_515),
.A2(n_481),
.B1(n_470),
.B2(n_478),
.Y(n_559)
);

INVx13_ASAP7_75t_L g560 ( 
.A(n_552),
.Y(n_560)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_560),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_561),
.A2(n_567),
.B1(n_574),
.B2(n_576),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_562),
.A2(n_570),
.B1(n_571),
.B2(n_536),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_563),
.B(n_565),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_524),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_568),
.A2(n_569),
.B(n_572),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_557),
.B(n_533),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_511),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_478),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_546),
.A2(n_505),
.B(n_470),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_575),
.B(n_577),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_549),
.A2(n_470),
.B1(n_469),
.B2(n_406),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_551),
.B(n_553),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_559),
.A2(n_470),
.B1(n_406),
.B2(n_301),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_578),
.B(n_579),
.Y(n_584)
);

BUFx24_ASAP7_75t_SL g583 ( 
.A(n_570),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_595),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_573),
.B(n_535),
.C(n_556),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_585),
.B(n_588),
.Y(n_600)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_586),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_535),
.C(n_537),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_542),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_589),
.B(n_596),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_564),
.B(n_537),
.C(n_558),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_590),
.B(n_592),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_564),
.B(n_538),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_544),
.B1(n_545),
.B2(n_539),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_594),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_566),
.A2(n_538),
.B1(n_392),
.B2(n_281),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_562),
.B(n_281),
.C(n_159),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_568),
.B(n_281),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_591),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_597),
.B(n_602),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_588),
.A2(n_563),
.B(n_567),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_601),
.A2(n_159),
.B(n_3),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_561),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_585),
.B(n_574),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_581),
.Y(n_612)
);

AOI21x1_ASAP7_75t_L g604 ( 
.A1(n_595),
.A2(n_566),
.B(n_569),
.Y(n_604)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_590),
.A2(n_571),
.B(n_565),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_605),
.A2(n_589),
.B(n_571),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_565),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_608),
.B(n_609),
.C(n_584),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_580),
.B(n_576),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_611),
.B(n_615),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_612),
.B(n_613),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_600),
.B(n_582),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_614),
.A2(n_616),
.B(n_617),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_606),
.B(n_596),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_L g616 ( 
.A(n_610),
.B(n_560),
.C(n_578),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_597),
.B(n_602),
.Y(n_617)
);

AOI31xp67_ASAP7_75t_L g620 ( 
.A1(n_608),
.A2(n_560),
.A3(n_584),
.B(n_579),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_620),
.B(n_1),
.C(n_4),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_621),
.A2(n_619),
.B(n_4),
.Y(n_628)
);

AOI322xp5_ASAP7_75t_L g623 ( 
.A1(n_618),
.A2(n_599),
.A3(n_598),
.B1(n_609),
.B2(n_607),
.C1(n_104),
.C2(n_93),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_624),
.C(n_8),
.Y(n_631)
);

AOI322xp5_ASAP7_75t_L g624 ( 
.A1(n_619),
.A2(n_607),
.A3(n_93),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_624)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_625),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_628),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g629 ( 
.A(n_626),
.B(n_1),
.C(n_4),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_629),
.A2(n_630),
.B(n_631),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_622),
.A2(n_7),
.B(n_8),
.Y(n_630)
);

AOI322xp5_ASAP7_75t_L g635 ( 
.A1(n_632),
.A2(n_627),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_16),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_635),
.B(n_633),
.C(n_10),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_636),
.A2(n_634),
.B(n_11),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_637),
.A2(n_9),
.B(n_11),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_9),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_13),
.Y(n_640)
);


endmodule