module fake_jpeg_16218_n_288 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_16),
.CON(n_52),
.SN(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_19),
.B1(n_15),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_15),
.B1(n_19),
.B2(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_16),
.A3(n_20),
.B1(n_25),
.B2(n_31),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_30),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_67),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_63),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_66),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_25),
.B(n_20),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_15),
.B1(n_29),
.B2(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_30),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_78),
.Y(n_97)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_40),
.B1(n_26),
.B2(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_77),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_36),
.B(n_21),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_90),
.B(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_50),
.B1(n_27),
.B2(n_37),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_93),
.B1(n_75),
.B2(n_73),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_21),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_100),
.B1(n_69),
.B2(n_28),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_71),
.B1(n_72),
.B2(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_62),
.Y(n_110)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_45),
.B(n_30),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_34),
.C(n_37),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_112),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_69),
.B1(n_50),
.B2(n_73),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_98),
.B1(n_84),
.B2(n_101),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_105),
.B1(n_88),
.B2(n_89),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_57),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_132),
.B1(n_98),
.B2(n_84),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_31),
.B(n_27),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_90),
.B(n_87),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_128),
.Y(n_138)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_56),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_56),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_27),
.B1(n_8),
.B2(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_56),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_153),
.B(n_131),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_158),
.B(n_130),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_92),
.B1(n_93),
.B2(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_149),
.B1(n_116),
.B2(n_1),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_126),
.B1(n_113),
.B2(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_92),
.C(n_101),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_152),
.C(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_89),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_99),
.B(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_162),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_0),
.B(n_1),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_53),
.C(n_6),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_53),
.C(n_6),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_114),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_167),
.B(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_110),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_180),
.Y(n_200)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_127),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_189),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_176),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_123),
.B1(n_109),
.B2(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_125),
.B1(n_115),
.B2(n_133),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_177),
.B1(n_186),
.B2(n_151),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_138),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_139),
.B(n_143),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_147),
.Y(n_180)
);

XNOR2x2_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_113),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_145),
.B1(n_161),
.B2(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_195),
.C(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_167),
.B1(n_170),
.B2(n_173),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_138),
.C(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_137),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_137),
.C(n_135),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_159),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_175),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_159),
.C(n_160),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_164),
.C(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_178),
.B(n_140),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_154),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_116),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_204),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_223),
.B1(n_205),
.B2(n_198),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_172),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_217),
.C(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_165),
.C(n_183),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_182),
.C(n_170),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_179),
.B1(n_168),
.B2(n_7),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_203),
.C(n_202),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_194),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_196),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_190),
.B(n_205),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_209),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_240),
.C(n_241),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_224),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_210),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_201),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_228),
.B(n_207),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_253),
.B(n_232),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_225),
.C(n_218),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_255),
.C(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_200),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_231),
.A2(n_211),
.B(n_214),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_211),
.C(n_1),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_251),
.B(n_255),
.Y(n_256)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_245),
.B(n_9),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_262),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_230),
.B(n_7),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_263),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_5),
.B1(n_10),
.B2(n_9),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_8),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_258),
.C(n_259),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_12),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_9),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_273),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_10),
.B(n_12),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_0),
.Y(n_277)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_279),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_2),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_280),
.A2(n_275),
.B(n_272),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_281),
.B(n_282),
.Y(n_284)
);

AOI321xp33_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_278),
.A3(n_274),
.B1(n_4),
.B2(n_3),
.C(n_2),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_286),
.A2(n_2),
.B(n_4),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_2),
.B(n_4),
.Y(n_288)
);


endmodule