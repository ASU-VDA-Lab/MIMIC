module fake_jpeg_26978_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_13),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_21),
.B1(n_35),
.B2(n_31),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_48),
.B1(n_34),
.B2(n_30),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_21),
.B1(n_26),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_23),
.B1(n_20),
.B2(n_25),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_35),
.B1(n_20),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_58),
.B1(n_25),
.B2(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_42),
.B1(n_46),
.B2(n_39),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_60),
.B1(n_43),
.B2(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_27),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_28),
.C(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_76),
.C(n_63),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_49),
.B(n_43),
.C(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_40),
.C(n_22),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_18),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

OAI211xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_65),
.B(n_63),
.C(n_55),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_61),
.B(n_53),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_87),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_89),
.B1(n_77),
.B2(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_75),
.B1(n_72),
.B2(n_63),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_95),
.B(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_101),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_70),
.B(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_88),
.C(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_89),
.C(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_110),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_117),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_100),
.B(n_73),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_115),
.B(n_110),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_25),
.B(n_24),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_8),
.B(n_11),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_123),
.C(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

AOI31xp67_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_104),
.A3(n_24),
.B(n_16),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_4),
.B(n_5),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_51),
.B1(n_74),
.B2(n_56),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_0),
.C(n_2),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_43),
.C(n_1),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_130),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_127),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_2),
.B(n_3),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_131),
.B(n_3),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_131),
.Y(n_135)
);


endmodule