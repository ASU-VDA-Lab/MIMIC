module fake_jpeg_13296_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_27),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

OR2x4_ASAP7_75t_SL g38 ( 
.A(n_12),
.B(n_0),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_20),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_12),
.Y(n_51)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_55),
.Y(n_75)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_19),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_24),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_28),
.A2(n_25),
.B(n_20),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_24),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_25),
.B1(n_13),
.B2(n_21),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_13),
.B1(n_22),
.B2(n_3),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_22),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_62),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_85),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_13),
.B1(n_2),
.B2(n_4),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_8),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_76),
.C(n_70),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_109),
.C(n_110),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_76),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_90),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_92),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_74),
.C(n_83),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_84),
.C(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_113),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_87),
.B(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_88),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_105),
.B(n_88),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_114),
.B(n_111),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_123),
.B(n_124),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_69),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_50),
.B(n_93),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_114),
.C(n_72),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.C(n_121),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_93),
.A3(n_73),
.B1(n_71),
.B2(n_2),
.C1(n_6),
.C2(n_69),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_93),
.B1(n_71),
.B2(n_48),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_72),
.C(n_50),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_131),
.B(n_48),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_6),
.B(n_53),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_6),
.B(n_63),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_45),
.Y(n_137)
);


endmodule