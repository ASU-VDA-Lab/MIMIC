module fake_jpeg_23026_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_17),
.B1(n_16),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_15),
.B1(n_25),
.B2(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_29),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_53),
.B1(n_25),
.B2(n_36),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_16),
.B1(n_17),
.B2(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_45),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_0),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_26),
.B(n_21),
.C(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_30),
.B1(n_18),
.B2(n_41),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_48),
.B(n_58),
.C(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_79),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_43),
.B1(n_37),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_82),
.B1(n_87),
.B2(n_59),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_84),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_85),
.Y(n_91)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_38),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_42),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_93),
.B1(n_77),
.B2(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_62),
.B1(n_38),
.B2(n_55),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_42),
.B(n_2),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_97),
.B(n_81),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_103),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_8),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_70),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_9),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_69),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_90),
.C(n_107),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_96),
.B(n_89),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_116),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_84),
.B(n_76),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_74),
.B1(n_87),
.B2(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_91),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_70),
.B1(n_4),
.B2(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_130),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_118),
.Y(n_142)
);

OAI221xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_90),
.B1(n_100),
.B2(n_107),
.C(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_100),
.C(n_101),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_140),
.C(n_116),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_102),
.A3(n_101),
.B1(n_8),
.B2(n_12),
.C(n_13),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_101),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_149),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_123),
.B1(n_114),
.B2(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_134),
.B1(n_130),
.B2(n_128),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_148),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_121),
.C(n_112),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_141),
.B1(n_127),
.B2(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_138),
.B(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_147),
.C(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_78),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_166),
.C(n_138),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_143),
.B(n_150),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_160),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_168),
.B(n_170),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_160),
.C(n_158),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_171),
.C(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_164),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_13),
.B(n_14),
.Y(n_177)
);

OAI21x1_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_176),
.B(n_14),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_113),
.Y(n_179)
);


endmodule