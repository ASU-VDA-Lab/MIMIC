module fake_jpeg_3933_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_40),
.B1(n_38),
.B2(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_35),
.C(n_41),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_27),
.C(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_59),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_18),
.B1(n_30),
.B2(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_77),
.B1(n_26),
.B2(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_78),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_25),
.B1(n_24),
.B2(n_28),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_22),
.B1(n_17),
.B2(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_83),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_17),
.B(n_24),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_26),
.B(n_31),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_69),
.B1(n_77),
.B2(n_60),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_90),
.B1(n_21),
.B2(n_19),
.Y(n_124)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_50),
.B1(n_22),
.B2(n_17),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_21),
.B1(n_19),
.B2(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_99),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_84),
.B(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_103),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_45),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_27),
.B(n_34),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_74),
.Y(n_105)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_46),
.C(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_113),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_98),
.B(n_104),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_118),
.C(n_122),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_116),
.B(n_93),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_90),
.B(n_88),
.C(n_96),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_68),
.B1(n_65),
.B2(n_75),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_34),
.C(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_34),
.C(n_64),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_126),
.B1(n_106),
.B2(n_99),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_21),
.B1(n_19),
.B2(n_34),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_101),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_104),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_142),
.B(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_141),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_120),
.B(n_118),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_155),
.B(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_144),
.Y(n_167)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_100),
.B1(n_97),
.B2(n_86),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_126),
.B(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_112),
.C(n_106),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_117),
.C(n_119),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_158),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_157),
.B1(n_61),
.B2(n_15),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_103),
.B(n_94),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_SL g180 ( 
.A(n_154),
.B(n_3),
.C(n_4),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_0),
.B(n_2),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_89),
.B1(n_72),
.B2(n_61),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_174),
.C(n_176),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_129),
.B1(n_108),
.B2(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_180),
.B1(n_141),
.B2(n_136),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_108),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_169),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_148),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_175),
.B1(n_150),
.B2(n_134),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_94),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_61),
.C(n_27),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_14),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_152),
.B1(n_151),
.B2(n_133),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_178),
.A2(n_146),
.B1(n_7),
.B2(n_8),
.Y(n_195)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_186),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_153),
.B(n_157),
.C(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_195),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_166),
.C(n_162),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_192),
.C(n_9),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_147),
.C(n_138),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_143),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_196),
.B(n_9),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_6),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_178),
.B1(n_160),
.B2(n_174),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_201),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_176),
.C(n_163),
.Y(n_201)
);

BUFx12_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_210),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_208),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_13),
.C(n_14),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_10),
.B1(n_11),
.B2(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_10),
.C(n_11),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_190),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_209),
.A2(n_204),
.B1(n_201),
.B2(n_199),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_218),
.B(n_212),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_189),
.CI(n_195),
.CON(n_215),
.SN(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_219),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_193),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_183),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_223),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_183),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_213),
.C(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_200),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_227),
.B(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_196),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_198),
.Y(n_231)
);

OAI221xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_207),
.B1(n_217),
.B2(n_215),
.C(n_219),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_222),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_225),
.B(n_202),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_235),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_224),
.B(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_10),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_233),
.B1(n_236),
.B2(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_242),
.B(n_238),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_247),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_245),
.Y(n_249)
);


endmodule