module fake_jpeg_23338_n_19 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_19;

wire n_13;
wire n_10;
wire n_14;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

OAI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_3),
.A2(n_9),
.B1(n_7),
.B2(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_14),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_11),
.B1(n_12),
.B2(n_6),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_15),
.B(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_1),
.Y(n_19)
);


endmodule