module fake_jpeg_23803_n_30 (n_3, n_2, n_1, n_0, n_4, n_5, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx13_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

HAxp5_ASAP7_75t_SL g11 ( 
.A(n_3),
.B(n_4),
.CON(n_11),
.SN(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_14),
.Y(n_18)
);

OAI21xp33_ASAP7_75t_SL g13 ( 
.A1(n_11),
.A2(n_0),
.B(n_2),
.Y(n_13)
);

MAJx2_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_8),
.C(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_15),
.B1(n_6),
.B2(n_17),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.C(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_8),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_14),
.B1(n_10),
.B2(n_4),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_18),
.B(n_21),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_25),
.B(n_20),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);


endmodule