module fake_jpeg_17163_n_33 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_3),
.B(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_0),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_25),
.B(n_20),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_1),
.B1(n_12),
.B2(n_17),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_26),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_15),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_18),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_21),
.B(n_23),
.Y(n_30)
);

OA21x2_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B(n_28),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_19),
.Y(n_33)
);


endmodule