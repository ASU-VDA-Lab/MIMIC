module fake_jpeg_11577_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_7),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_59),
.Y(n_110)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_16),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_68),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_65),
.Y(n_113)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_17),
.B(n_7),
.Y(n_66)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_15),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_17),
.B1(n_18),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_73),
.A2(n_94),
.B1(n_100),
.B2(n_28),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_29),
.B1(n_37),
.B2(n_32),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_36),
.B1(n_20),
.B2(n_37),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_78),
.A2(n_114),
.B1(n_24),
.B2(n_31),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_29),
.B1(n_37),
.B2(n_36),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_36),
.B1(n_20),
.B2(n_37),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_109),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_17),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_18),
.B1(n_35),
.B2(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_40),
.A2(n_35),
.B1(n_33),
.B2(n_27),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_36),
.C(n_20),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_61),
.C(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_33),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_19),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_141),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_117),
.C(n_139),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_31),
.B(n_24),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_122),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_78),
.B1(n_63),
.B2(n_26),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_131),
.B1(n_133),
.B2(n_136),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_148),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_71),
.B1(n_67),
.B2(n_41),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_135),
.B1(n_152),
.B2(n_156),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_27),
.B1(n_26),
.B2(n_50),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_49),
.B1(n_45),
.B2(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_72),
.C(n_62),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_43),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_77),
.B(n_15),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_150),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_84),
.B(n_42),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_84),
.B(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_86),
.B(n_38),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_38),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_91),
.A2(n_24),
.B1(n_31),
.B2(n_25),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_107),
.B1(n_93),
.B2(n_99),
.Y(n_181)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_91),
.A2(n_38),
.B1(n_52),
.B2(n_31),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_99),
.B(n_96),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_178),
.B(n_81),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_166),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_169),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_95),
.B(n_24),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_132),
.B1(n_142),
.B2(n_129),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_39),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_123),
.B(n_97),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_123),
.B(n_97),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_101),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_60),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_120),
.A2(n_96),
.B1(n_82),
.B2(n_101),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_130),
.B1(n_156),
.B2(n_134),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_115),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_197),
.B(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_116),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_210),
.C(n_229),
.Y(n_241)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_142),
.B1(n_132),
.B2(n_145),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_148),
.B1(n_119),
.B2(n_154),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_120),
.B1(n_150),
.B2(n_107),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_215),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_120),
.B1(n_126),
.B2(n_146),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_151),
.B1(n_153),
.B2(n_144),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_208),
.B1(n_225),
.B2(n_231),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_151),
.B1(n_146),
.B2(n_126),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_209),
.A2(n_226),
.B(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_143),
.C(n_138),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_173),
.A2(n_80),
.B1(n_81),
.B2(n_155),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_228),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_214),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_173),
.A2(n_80),
.B1(n_138),
.B2(n_55),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_179),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_159),
.Y(n_238)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_125),
.B1(n_128),
.B2(n_55),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_125),
.B(n_65),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_0),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_163),
.B(n_65),
.C(n_0),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_169),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_163),
.A2(n_6),
.B(n_1),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_239),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_197),
.B(n_162),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_251),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_162),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_246),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_165),
.C(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_254),
.C(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_201),
.B(n_185),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_165),
.C(n_194),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_159),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_172),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_160),
.C(n_164),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_267),
.C(n_9),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_206),
.A2(n_164),
.B1(n_180),
.B2(n_177),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_203),
.B1(n_223),
.B2(n_222),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_180),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_262),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_234),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_264),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_170),
.B(n_167),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_268),
.B(n_267),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_170),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_192),
.C(n_187),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_232),
.A2(n_186),
.B(n_184),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_208),
.B1(n_207),
.B2(n_205),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_271),
.A2(n_273),
.B1(n_282),
.B2(n_268),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_215),
.B(n_212),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_220),
.B1(n_224),
.B2(n_219),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_277),
.B1(n_280),
.B2(n_284),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_213),
.B1(n_217),
.B2(n_211),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_SL g278 ( 
.A1(n_240),
.A2(n_219),
.B(n_200),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_278),
.A2(n_270),
.B1(n_259),
.B2(n_249),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_225),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_296),
.C(n_297),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_199),
.B1(n_233),
.B2(n_157),
.Y(n_280)
);

AO22x1_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_184),
.B1(n_186),
.B2(n_188),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_233),
.B1(n_188),
.B2(n_157),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_176),
.B1(n_187),
.B2(n_231),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_286),
.A2(n_287),
.B1(n_248),
.B2(n_258),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_254),
.B1(n_265),
.B2(n_256),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_257),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_235),
.A2(n_176),
.B1(n_214),
.B2(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_290),
.Y(n_314)
);

OAI32xp33_ASAP7_75t_L g293 ( 
.A1(n_253),
.A2(n_214),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_214),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_241),
.B(n_9),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_250),
.C(n_252),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_0),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_272),
.Y(n_309)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_310),
.A2(n_319),
.B1(n_323),
.B2(n_286),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_244),
.B(n_257),
.Y(n_329)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_255),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_316),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_271),
.A2(n_274),
.B1(n_279),
.B2(n_282),
.Y(n_319)
);

XOR2x2_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_259),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_283),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_297),
.C(n_281),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_252),
.B1(n_249),
.B2(n_263),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_14),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_272),
.B1(n_300),
.B2(n_276),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_336),
.B1(n_311),
.B2(n_322),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_332),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_331),
.B1(n_342),
.B2(n_343),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_319),
.A2(n_287),
.B1(n_275),
.B2(n_284),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_340),
.C(n_346),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_293),
.C(n_294),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_306),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_263),
.C(n_0),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_310),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_306),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_343)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_3),
.C(n_4),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_9),
.C(n_10),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_321),
.C(n_324),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_344),
.Y(n_350)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_307),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_353),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_365),
.B1(n_342),
.B2(n_320),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_338),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_333),
.B(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_357),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_312),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_317),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_360),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_359),
.A2(n_336),
.B1(n_348),
.B2(n_305),
.Y(n_369)
);

AO22x1_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_326),
.B1(n_305),
.B2(n_323),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_363),
.Y(n_377)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_334),
.C(n_304),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_364),
.B(n_328),
.C(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_366),
.B(n_367),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_334),
.C(n_337),
.Y(n_367)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_331),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_378),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_340),
.C(n_330),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_373),
.A2(n_356),
.B(n_361),
.Y(n_385)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_350),
.A2(n_343),
.B1(n_301),
.B2(n_314),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_376),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_347),
.Y(n_378)
);

OAI221xp5_ASAP7_75t_L g379 ( 
.A1(n_349),
.A2(n_357),
.B1(n_358),
.B2(n_356),
.C(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_374),
.A2(n_349),
.B1(n_361),
.B2(n_360),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_388),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_385),
.B(n_387),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_367),
.A2(n_360),
.B(n_362),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_373),
.B(n_371),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_318),
.Y(n_387)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_380),
.Y(n_391)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_391),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_396),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_389),
.B(n_377),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_394),
.A2(n_371),
.B1(n_12),
.B2(n_14),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_368),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_395),
.B(n_397),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_378),
.B(n_390),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_381),
.A2(n_366),
.B(n_383),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_390),
.C(n_387),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_400),
.B(n_401),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_14),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_404),
.Y(n_408)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_400),
.B(n_395),
.CI(n_398),
.CON(n_406),
.SN(n_406)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_407),
.Y(n_411)
);

OAI211xp5_ASAP7_75t_L g407 ( 
.A1(n_405),
.A2(n_399),
.B(n_12),
.C(n_14),
.Y(n_407)
);

AOI21x1_ASAP7_75t_L g410 ( 
.A1(n_409),
.A2(n_403),
.B(n_402),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_410),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_411),
.B(n_402),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g414 ( 
.A1(n_413),
.A2(n_408),
.B(n_10),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_414),
.B(n_12),
.Y(n_415)
);


endmodule