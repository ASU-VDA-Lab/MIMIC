module fake_jpeg_13649_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g85 ( 
.A(n_39),
.Y(n_85)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_38),
.Y(n_81)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_59),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_17),
.B1(n_21),
.B2(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_84),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_45),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_77),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_33),
.B(n_25),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_88),
.B(n_96),
.C(n_85),
.D(n_71),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_28),
.B1(n_37),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_34),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_34),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_50),
.Y(n_116)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_102),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_109),
.Y(n_166)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_37),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_50),
.B1(n_42),
.B2(n_24),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_126),
.B1(n_134),
.B2(n_136),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_65),
.B(n_78),
.C(n_92),
.Y(n_164)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_35),
.B1(n_23),
.B2(n_30),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_30),
.B1(n_33),
.B2(n_25),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_0),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_47),
.B1(n_54),
.B2(n_10),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_54),
.C(n_47),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_90),
.B(n_72),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_143),
.A2(n_162),
.B(n_165),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_99),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_103),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_162),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_103),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_157),
.Y(n_191)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_158),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_14),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_163),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_65),
.B1(n_68),
.B2(n_90),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_68),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_101),
.B1(n_86),
.B2(n_92),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_169),
.B1(n_137),
.B2(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_113),
.A2(n_101),
.B1(n_92),
.B2(n_67),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_108),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_173),
.B(n_8),
.Y(n_207)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_185),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_189),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_130),
.B1(n_121),
.B2(n_131),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_178),
.A2(n_168),
.B1(n_152),
.B2(n_165),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_143),
.A2(n_104),
.B(n_107),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_208),
.B(n_176),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_104),
.C(n_107),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_171),
.C(n_166),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_147),
.A2(n_161),
.B1(n_142),
.B2(n_144),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_196),
.B1(n_169),
.B2(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_137),
.B1(n_124),
.B2(n_114),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_67),
.B1(n_10),
.B2(n_15),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_140),
.B(n_9),
.CI(n_15),
.CON(n_199),
.SN(n_199)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_200),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_69),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_208),
.B(n_0),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_145),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_157),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_220),
.B1(n_190),
.B2(n_186),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_3),
.B(n_4),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_213),
.B(n_236),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_139),
.C(n_166),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_202),
.C(n_175),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_223),
.B1(n_209),
.B2(n_193),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_168),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_152),
.B1(n_138),
.B2(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_235),
.B1(n_1),
.B2(n_2),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_0),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_176),
.B(n_202),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_14),
.B(n_8),
.Y(n_260)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_180),
.B(n_182),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_246),
.C(n_216),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_251),
.B1(n_214),
.B2(n_215),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_199),
.B1(n_194),
.B2(n_203),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_253),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_199),
.B1(n_203),
.B2(n_198),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_243),
.A2(n_250),
.B1(n_220),
.B2(n_234),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_186),
.C(n_206),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_198),
.B1(n_193),
.B2(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_209),
.B1(n_191),
.B2(n_3),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_191),
.B1(n_10),
.B2(n_3),
.Y(n_253)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_8),
.B(n_11),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_224),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_233),
.Y(n_275)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_221),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_270),
.C(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_244),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_248),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_262),
.B1(n_240),
.B2(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_219),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_271),
.B(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_237),
.C(n_232),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_253),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_226),
.C(n_210),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_235),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_222),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_283),
.B(n_286),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_290),
.C(n_292),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_272),
.B1(n_250),
.B2(n_264),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_287),
.B(n_249),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_257),
.B(n_242),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_241),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_301),
.Y(n_309)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_307),
.Y(n_313)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_277),
.B1(n_248),
.B2(n_275),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_290),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_314),
.B1(n_284),
.B2(n_297),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_281),
.B(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_312),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_292),
.C(n_291),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_223),
.B1(n_247),
.B2(n_255),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_283),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_210),
.C(n_227),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_300),
.B1(n_301),
.B2(n_306),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_313),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_298),
.B1(n_259),
.B2(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_286),
.CI(n_297),
.CON(n_321),
.SN(n_321)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_322),
.B(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_308),
.C(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_320),
.B1(n_322),
.B2(n_321),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.C(n_326),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_314),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_315),
.B(n_229),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_231),
.C(n_217),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_214),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_13),
.Y(n_336)
);


endmodule