module real_jpeg_3820_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_0),
.A2(n_54),
.B1(n_223),
.B2(n_326),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_0),
.A2(n_54),
.B1(n_178),
.B2(n_179),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_0),
.A2(n_54),
.B1(n_345),
.B2(n_410),
.Y(n_409)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_1),
.Y(n_210)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_1),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_2),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_2),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_2),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_2),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_97),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_3),
.A2(n_97),
.B1(n_220),
.B2(n_394),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_4),
.A2(n_139),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_4),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_4),
.A2(n_152),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_4),
.A2(n_152),
.B1(n_374),
.B2(n_377),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_4),
.A2(n_152),
.B1(n_405),
.B2(n_408),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_5),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_60),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_6),
.A2(n_60),
.B1(n_237),
.B2(n_245),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_6),
.A2(n_60),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_7),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_7),
.A2(n_51),
.B1(n_91),
.B2(n_138),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_7),
.A2(n_91),
.B1(n_296),
.B2(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_7),
.A2(n_91),
.B1(n_377),
.B2(n_420),
.Y(n_419)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_8),
.Y(n_343)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_9),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_10),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_10),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_10),
.A2(n_184),
.B1(n_219),
.B2(n_223),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_10),
.A2(n_184),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_10),
.A2(n_184),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_11),
.Y(n_193)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_15),
.A2(n_199),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_15),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_15),
.A2(n_203),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_15),
.A2(n_203),
.B1(n_286),
.B2(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_15),
.A2(n_203),
.B1(n_413),
.B2(n_415),
.Y(n_412)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_17),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_17),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_17),
.B(n_193),
.C(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_17),
.B(n_72),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_17),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_17),
.B(n_187),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_17),
.B(n_281),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_18),
.A2(n_77),
.B1(n_178),
.B2(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_18),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_18),
.A2(n_229),
.B1(n_244),
.B2(n_249),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_18),
.A2(n_45),
.B1(n_229),
.B2(n_288),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_18),
.A2(n_31),
.B1(n_32),
.B2(n_229),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_510),
.B(n_513),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_167),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_165),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_143),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_23),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_131),
.B2(n_132),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_61),
.C(n_98),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_26),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_55),
.B1(n_57),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_27),
.A2(n_47),
.B1(n_55),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_27),
.A2(n_364),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_27),
.A2(n_38),
.B1(n_412),
.B2(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_28),
.A2(n_361),
.B(n_363),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_28),
.B(n_365),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_33),
.Y(n_340)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_38),
.B(n_180),
.Y(n_323)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_40),
.Y(n_278)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_41),
.Y(n_161)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_43),
.Y(n_407)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_50),
.Y(n_362)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_55),
.A2(n_433),
.B(n_455),
.Y(n_465)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_56),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_56),
.B(n_151),
.Y(n_454)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_98),
.B1(n_99),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_84),
.B1(n_92),
.B2(n_93),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_62),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_62),
.A2(n_84),
.B1(n_92),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_62),
.A2(n_92),
.B1(n_319),
.B2(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_62),
.A2(n_92),
.B1(n_404),
.B2(n_409),
.Y(n_403)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_72),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_63)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_64),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_71),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_71),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_71),
.Y(n_371)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g434 ( 
.A1(n_72),
.A2(n_134),
.B1(n_321),
.B2(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_72),
.A2(n_134),
.B1(n_160),
.B2(n_443),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_75),
.Y(n_306)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_77),
.B(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_77),
.Y(n_399)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_78),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_80),
.Y(n_376)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_80),
.Y(n_379)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_86),
.Y(n_287)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_90),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_92),
.B(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_92),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_94),
.Y(n_410)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_149),
.C(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_98),
.A2(n_99),
.B1(n_157),
.B2(n_158),
.Y(n_499)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_116),
.B(n_125),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_100),
.A2(n_177),
.B(n_181),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_100),
.A2(n_116),
.B1(n_228),
.B2(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_100),
.A2(n_181),
.B(n_271),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_100),
.A2(n_116),
.B1(n_373),
.B2(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_101),
.B(n_182),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_101),
.A2(n_187),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_101),
.A2(n_187),
.B1(n_398),
.B2(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_101),
.A2(n_187),
.B1(n_419),
.B2(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_109),
.B2(n_113),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx5_ASAP7_75t_SL g305 ( 
.A(n_113),
.Y(n_305)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_116),
.A2(n_228),
.B(n_230),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_116),
.A2(n_230),
.B(n_373),
.Y(n_372)
);

AOI22x1_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_119),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_120),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_120),
.Y(n_395)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_125),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_130),
.Y(n_420)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_134),
.A2(n_277),
.B(n_284),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_134),
.B(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_134),
.A2(n_284),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_139),
.B(n_180),
.Y(n_349)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_155),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_505)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_148),
.A2(n_149),
.B1(n_499),
.B2(n_500),
.Y(n_498)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_155),
.A2(n_156),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_494),
.B(n_507),
.Y(n_168)
);

OAI311xp33_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_382),
.A3(n_470),
.B1(n_488),
.C1(n_489),
.Y(n_169)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_332),
.B(n_381),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_310),
.B(n_331),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_265),
.B(n_309),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_233),
.B(n_264),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_196),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_175),
.B(n_196),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_188),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_176),
.A2(n_188),
.B1(n_189),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_207),
.B(n_214),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_180),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_SL g361 ( 
.A1(n_180),
.A2(n_349),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_225),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_197),
.B(n_226),
.C(n_232),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_207),
.B(n_214),
.Y(n_197)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_207),
.A2(n_216),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_207),
.A2(n_388),
.B1(n_391),
.B2(n_393),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_207),
.A2(n_216),
.B(n_393),
.Y(n_421)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_218),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_208),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_208),
.A2(n_294),
.B1(n_325),
.B2(n_328),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_208),
.A2(n_354),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_210),
.Y(n_329)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_213),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_243),
.B(n_252),
.Y(n_242)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_255),
.B(n_263),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_241),
.B(n_254),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_253),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_253),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_293),
.B(n_299),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_261),
.Y(n_263)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_267),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_291),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_275),
.C(n_291),
.Y(n_311)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_274),
.Y(n_401)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_303),
.A3(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_290),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_302),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

INVx4_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_311),
.B(n_312),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_317),
.B2(n_330),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_316),
.C(n_330),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_322),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_323),
.C(n_324),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_333),
.B(n_334),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_358),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_335)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_350),
.B2(n_351),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_338),
.B(n_350),
.Y(n_466)
);

OAI32xp33_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.A3(n_341),
.B1(n_344),
.B2(n_349),
.Y(n_338)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_355),
.B(n_357),
.C(n_358),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_368),
.B2(n_380),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_359),
.B(n_369),
.C(n_372),
.Y(n_479)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_456),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_383),
.A2(n_456),
.B(n_490),
.C(n_493),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_436),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_384),
.B(n_436),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_416),
.C(n_423),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_385),
.B(n_416),
.CI(n_423),
.CON(n_469),
.SN(n_469)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_402),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_403),
.C(n_411),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_396),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_387),
.B(n_396),
.Y(n_462)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_411),
.Y(n_402)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx6_ASAP7_75t_SL g406 ( 
.A(n_407),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_421),
.B2(n_422),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_421),
.Y(n_450)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_421),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_421),
.A2(n_422),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_421),
.A2(n_450),
.B(n_453),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_431),
.C(n_434),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_427),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_427),
.Y(n_478)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_431),
.A2(n_432),
.B1(n_434),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_434),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_437),
.B(n_440),
.C(n_448),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_448),
.B2(n_449),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_444),
.B(n_447),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_442),
.B(n_445),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g496 ( 
.A(n_447),
.B(n_497),
.CI(n_498),
.CON(n_496),
.SN(n_496)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_497),
.C(n_498),
.Y(n_506)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_469),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_469),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_462),
.C(n_463),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_458),
.A2(n_459),
.B1(n_462),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.C(n_467),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_466),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_467),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_469),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_483),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_472),
.A2(n_491),
.B(n_492),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_480),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_480),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.C(n_479),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_486),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_478),
.B1(n_479),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_479),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_484),
.B(n_485),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_502),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_501),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_501),
.Y(n_508)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_496),
.Y(n_517)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_499),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_502),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_506),
.Y(n_509)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx4f_ASAP7_75t_SL g510 ( 
.A(n_511),
.Y(n_510)
);

INVx13_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx6_ASAP7_75t_L g514 ( 
.A(n_512),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);


endmodule