module real_jpeg_6396_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_31;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B1(n_38),
.B2(n_39),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_29),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_7),
.C(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_35),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_11),
.C(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_17),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_19),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_18),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B(n_37),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B(n_36),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_33),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_43),
.C(n_44),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_41),
.C(n_45),
.Y(n_40)
);


endmodule