module fake_jpeg_20086_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_20),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_11),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_9),
.B(n_13),
.C(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_12),
.B1(n_11),
.B2(n_17),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_9),
.C(n_13),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_11),
.B1(n_8),
.B2(n_19),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_15),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_28),
.B(n_2),
.C(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_36),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_26),
.B1(n_28),
.B2(n_23),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_31),
.B(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_47),
.B(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_46),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_0),
.B(n_52),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_0),
.Y(n_57)
);


endmodule