module real_jpeg_17054_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_0),
.B(n_61),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_0),
.A2(n_84),
.A3(n_275),
.B1(n_276),
.B2(n_279),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_0),
.A2(n_30),
.B1(n_186),
.B2(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_0),
.B(n_100),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_0),
.A2(n_157),
.B1(n_172),
.B2(n_406),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_1),
.A2(n_26),
.B1(n_70),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_1),
.A2(n_70),
.B1(n_280),
.B2(n_309),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_1),
.A2(n_70),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_55),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_2),
.A2(n_55),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_2),
.A2(n_55),
.B1(n_407),
.B2(n_409),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_3),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_3),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_3),
.A2(n_116),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_3),
.A2(n_116),
.B1(n_287),
.B2(n_292),
.Y(n_286)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_5),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_5),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_6),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_147),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_7),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g417 ( 
.A(n_7),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_8),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_8),
.A2(n_167),
.B1(n_235),
.B2(n_240),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_9),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_9),
.Y(n_278)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_102),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_10),
.A2(n_107),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_10),
.A2(n_107),
.B1(n_361),
.B2(n_364),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_12),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_14),
.A2(n_174),
.B1(n_175),
.B2(n_180),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_14),
.Y(n_180)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_15),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_15),
.Y(n_254)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_262),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_261),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_212),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_21),
.B(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_155),
.C(n_189),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_22),
.B(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_23),
.B(n_63),
.C(n_114),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B1(n_54),
.B2(n_61),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_30),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_30),
.B(n_339),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_30),
.A2(n_338),
.B(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_30),
.B(n_402),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_30),
.B(n_154),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_31),
.A2(n_65),
.B1(n_182),
.B2(n_188),
.Y(n_181)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_34),
.A2(n_54),
.B1(n_61),
.B2(n_218),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B(n_44),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_37),
.Y(n_185)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_39),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_40),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_50),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_114),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_75),
.B1(n_100),
.B2(n_101),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_64),
.A2(n_75),
.B1(n_100),
.B2(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_65),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_67),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_76),
.A2(n_223),
.B1(n_224),
.B2(n_229),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_76),
.A2(n_192),
.B1(n_229),
.B2(n_315),
.Y(n_314)
);

AO21x2_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_89),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_82),
.Y(n_193)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_91),
.Y(n_239)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_91),
.Y(n_283)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_100),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_101),
.Y(n_223)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_113),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_124),
.B1(n_144),
.B2(n_153),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_115),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_119),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_119),
.Y(n_353)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_124),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_124),
.A2(n_153),
.B1(n_296),
.B2(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_124),
.A2(n_153),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_124),
.A2(n_153),
.B1(n_308),
.B2(n_352),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_136),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_128),
.B1(n_131),
.B2(n_134),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_137),
.B1(n_139),
.B2(n_142),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_129),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_131),
.Y(n_331)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_133),
.Y(n_291)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_133),
.Y(n_367)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_137),
.Y(n_297)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_141),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_145),
.A2(n_154),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_154),
.A2(n_233),
.B1(n_295),
.B2(n_301),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_155),
.B(n_189),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_181),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_181),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_164),
.B1(n_172),
.B2(n_173),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_157),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_157),
.A2(n_173),
.B1(n_244),
.B2(n_255),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_157),
.A2(n_360),
.B1(n_368),
.B2(n_371),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_157),
.A2(n_381),
.B1(n_406),
.B2(n_414),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_158),
.A2(n_201),
.B1(n_202),
.B2(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_158),
.A2(n_201),
.B1(n_380),
.B2(n_389),
.Y(n_379)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_163),
.Y(n_363)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_163),
.Y(n_388)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_165),
.A2(n_201),
.B1(n_202),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.C(n_211),
.Y(n_189)
);

XOR2x1_ASAP7_75t_L g269 ( 
.A(n_190),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_200),
.B(n_211),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_230),
.B2(n_260),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2x1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_259),
.Y(n_230)
);

XOR2x2_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_238),
.Y(n_329)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_239),
.Y(n_357)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_253),
.Y(n_400)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_253),
.Y(n_411)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_254),
.Y(n_346)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_256),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_257),
.Y(n_404)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_429),
.B(n_433),
.Y(n_264)
);

OAI21x1_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_322),
.B(n_428),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_304),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_267),
.B(n_304),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_268),
.B(n_294),
.C(n_302),
.Y(n_432)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_294),
.B1(n_302),
.B2(n_303),
.Y(n_272)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_284),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_284),
.B1(n_285),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_286),
.Y(n_371)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_290),
.Y(n_383)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_313),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_305),
.B(n_425),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_307),
.A2(n_313),
.B1(n_314),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_307),
.Y(n_426)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_422),
.B(n_427),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_377),
.B(n_421),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_358),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_325),
.B(n_358),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_347),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_327),
.A2(n_347),
.B1(n_348),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_330),
.A3(n_332),
.B1(n_338),
.B2(n_340),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_372),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_359),
.B(n_374),
.C(n_376),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.Y(n_372)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_373),
.Y(n_376)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

AOI21x1_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_392),
.B(n_420),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_390),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_390),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_412),
.B(n_419),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_405),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_401),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_399),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_418),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_418),
.Y(n_419)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_424),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_432),
.Y(n_433)
);


endmodule