module fake_jpeg_28513_n_90 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_16),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_12),
.A3(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_54),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_9),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_64),
.B1(n_42),
.B2(n_44),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_60),
.Y(n_69)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_26),
.A2(n_7),
.B1(n_8),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_76),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_70),
.C(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_27),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_62),
.C(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_45),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_73),
.B(n_68),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.C(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_81),
.B(n_69),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_65),
.B(n_67),
.C(n_63),
.D(n_52),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_73),
.B(n_69),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_8),
.B(n_40),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_64),
.B(n_41),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);


endmodule