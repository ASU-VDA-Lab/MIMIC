module fake_jpeg_12847_n_68 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_22;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_28;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_2),
.B(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_20),
.A2(n_4),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_39),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_32),
.Y(n_49)
);

OR2x4_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_52),
.C(n_24),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_50),
.C(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_49),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_47),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_34),
.C(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_22),
.B1(n_28),
.B2(n_26),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_36),
.C(n_46),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_30),
.B(n_38),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_33),
.B(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_46),
.C(n_45),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_66),
.C(n_43),
.Y(n_68)
);


endmodule