module fake_jpeg_16943_n_358 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_9),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_0),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_35),
.B(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_48),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_10),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_82),
.B1(n_101),
.B2(n_118),
.Y(n_126)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_87),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_19),
.B1(n_28),
.B2(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_42),
.B1(n_19),
.B2(n_24),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_16),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_66),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_40),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_102),
.C(n_103),
.Y(n_133)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_92),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_34),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_31),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_21),
.B1(n_36),
.B2(n_35),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_47),
.C(n_34),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_37),
.C(n_34),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_18),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_34),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_14),
.B1(n_16),
.B2(n_15),
.Y(n_145)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_1),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_1),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_112),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_89),
.B1(n_105),
.B2(n_114),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_118),
.B1(n_116),
.B2(n_119),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_134),
.B1(n_119),
.B2(n_94),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_128),
.B(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_53),
.B1(n_52),
.B2(n_45),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_53),
.C(n_52),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_102),
.C(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_34),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_97),
.B(n_37),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_89),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_79),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_161),
.Y(n_196)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_157),
.A2(n_168),
.B1(n_131),
.B2(n_95),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_164),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_80),
.B1(n_124),
.B2(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_92),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_164),
.B(n_176),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_171),
.C(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_100),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_109),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_116),
.B1(n_113),
.B2(n_104),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_147),
.B1(n_140),
.B2(n_131),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_173),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_93),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_106),
.C(n_115),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_85),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_108),
.C(n_45),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_130),
.C(n_136),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_178),
.Y(n_194)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_125),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_32),
.C(n_18),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_125),
.B(n_141),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_185),
.B(n_189),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_128),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_134),
.B1(n_135),
.B2(n_139),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_195),
.B1(n_205),
.B2(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_141),
.B1(n_139),
.B2(n_151),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_204),
.B(n_169),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_145),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_130),
.B(n_150),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_169),
.B(n_174),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_138),
.B(n_129),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_117),
.B1(n_136),
.B2(n_147),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_R g207 ( 
.A(n_163),
.B(n_124),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_169),
.B1(n_160),
.B2(n_162),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_55),
.B1(n_54),
.B2(n_41),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_83),
.B1(n_174),
.B2(n_23),
.Y(n_230)
);

OAI22x1_ASAP7_75t_L g262 ( 
.A1(n_211),
.A2(n_230),
.B1(n_232),
.B2(n_23),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_200),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_218),
.B(n_223),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_219),
.A2(n_222),
.B1(n_192),
.B2(n_26),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_194),
.A2(n_168),
.B1(n_157),
.B2(n_152),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_18),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_195),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_174),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_182),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_11),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_236),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_198),
.A2(n_23),
.B(n_26),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_181),
.A2(n_11),
.B(n_15),
.C(n_14),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_32),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_32),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_37),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_192),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_186),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_239),
.C(n_225),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_191),
.B1(n_189),
.B2(n_202),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_255),
.B1(n_262),
.B2(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_220),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_205),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_185),
.B1(n_204),
.B2(n_184),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_210),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_260),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_193),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_221),
.B1(n_220),
.B2(n_234),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_239),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_273),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_269),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_280),
.C(n_282),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_252),
.C(n_244),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_247),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_212),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_277),
.B1(n_262),
.B2(n_247),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_215),
.B1(n_238),
.B2(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_197),
.C(n_212),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_263),
.B1(n_245),
.B2(n_233),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_254),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_215),
.C(n_229),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_285),
.C(n_241),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_226),
.C(n_224),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_232),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_244),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_304),
.Y(n_317)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

BUFx4f_ASAP7_75t_SL g292 ( 
.A(n_272),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_241),
.CI(n_231),
.CON(n_294),
.SN(n_294)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_294),
.B(n_26),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_266),
.C(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_263),
.C(n_242),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_12),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_274),
.B(n_230),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_278),
.A2(n_270),
.B(n_277),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_1),
.B(n_3),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_245),
.B1(n_2),
.B2(n_3),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_267),
.B1(n_276),
.B2(n_5),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_285),
.C(n_275),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_321),
.C(n_306),
.Y(n_325)
);

BUFx12_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_10),
.C(n_13),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_1),
.B(n_3),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_331),
.C(n_332),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_308),
.B(n_288),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_330),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_295),
.B1(n_296),
.B2(n_299),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_327),
.B(n_307),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_297),
.C(n_302),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_302),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_316),
.B(n_311),
.Y(n_333)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

NOR2x1_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_311),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_336),
.Y(n_342)
);

INVx11_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_341),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_307),
.B(n_313),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_323),
.B1(n_310),
.B2(n_328),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_334),
.Y(n_346)
);

AOI322xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_340),
.A3(n_339),
.B1(n_321),
.B2(n_333),
.C1(n_309),
.C2(n_331),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_338),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_349),
.B(n_343),
.Y(n_351)
);

AOI221xp5_ASAP7_75t_L g353 ( 
.A1(n_351),
.A2(n_352),
.B1(n_342),
.B2(n_338),
.C(n_332),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_350),
.A2(n_347),
.B(n_341),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_290),
.C(n_317),
.Y(n_354)
);

NAND4xp25_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_290),
.C(n_289),
.D(n_304),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_3),
.Y(n_356)
);

A2O1A1O1Ixp25_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_5),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_357)
);

AOI221xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_6),
.B1(n_7),
.B2(n_37),
.C(n_334),
.Y(n_358)
);


endmodule