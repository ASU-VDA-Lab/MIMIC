module fake_jpeg_13735_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_42),
.B1(n_43),
.B2(n_41),
.Y(n_60)
);

NAND2xp67_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_44),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_56),
.B1(n_38),
.B2(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_44),
.B1(n_45),
.B2(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_15),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_49),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_49),
.B(n_22),
.C(n_23),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_14),
.B(n_29),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_85),
.B1(n_8),
.B2(n_13),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_86),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_87),
.Y(n_91)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_92),
.Y(n_98)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_81),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

NAND4xp25_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_96),
.C(n_98),
.D(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_94),
.Y(n_107)
);


endmodule