module real_jpeg_22952_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_0),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_0),
.B(n_33),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_0),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_0),
.B(n_103),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_0),
.B(n_75),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_0),
.B(n_57),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_103),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_2),
.B(n_75),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_33),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_2),
.B(n_29),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_3),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_75),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_57),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_33),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_3),
.B(n_29),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_3),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_3),
.B(n_36),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_103),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_75),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_5),
.B(n_29),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_5),
.B(n_25),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_10),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_10),
.B(n_17),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_10),
.B(n_57),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_10),
.B(n_33),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_29),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_10),
.B(n_25),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_10),
.B(n_54),
.Y(n_270)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_12),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_12),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_12),
.B(n_75),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_12),
.B(n_57),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_12),
.B(n_33),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_12),
.B(n_29),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_12),
.B(n_54),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_14),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_14),
.B(n_173),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_14),
.B(n_75),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_14),
.B(n_57),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_14),
.B(n_33),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_15),
.B(n_57),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_15),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_29),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_15),
.B(n_25),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_16),
.B(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_16),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_16),
.B(n_57),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_33),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_29),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_16),
.B(n_25),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_16),
.B(n_36),
.Y(n_253)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.C(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_52),
.C(n_55),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_49),
.B1(n_55),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_33),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_43),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_43),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_44),
.B(n_124),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_44),
.B(n_250),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_51),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_53),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_72),
.C(n_74),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_55),
.A2(n_74),
.B1(n_79),
.B2(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_56),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_56),
.B(n_73),
.Y(n_261)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.C(n_81),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_60),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.C(n_77),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_61),
.B(n_372),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_62),
.B(n_81),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.CI(n_65),
.CON(n_62),
.SN(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.C(n_69),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_66),
.B(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_71),
.B(n_77),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_72),
.B(n_353),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_74),
.A2(n_299),
.B1(n_300),
.B2(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_74),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_SL g357 ( 
.A(n_74),
.B(n_299),
.C(n_326),
.Y(n_357)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_376),
.C(n_377),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_367),
.C(n_368),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_345),
.C(n_346),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_321),
.C(n_322),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_289),
.C(n_290),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_255),
.C(n_256),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_220),
.C(n_221),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_188),
.C(n_189),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_167),
.C(n_168),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_147),
.C(n_148),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_125),
.C(n_126),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.C(n_115),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_106),
.B2(n_107),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_108),
.C(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_103),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.C(n_120),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_124),
.B(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.C(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_146),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_151),
.C(n_156),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_166),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_182),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_183),
.C(n_187),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_177),
.C(n_178),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_176),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_178),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.CI(n_181),
.CON(n_178),
.SN(n_178)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.CI(n_186),
.CON(n_183),
.SN(n_183)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_204),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_193),
.C(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_200),
.C(n_203),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_195),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.CI(n_198),
.CON(n_195),
.SN(n_195)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_211),
.C(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_211),
.B1(n_218),
.B2(n_219),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_210),
.B(n_245),
.C(n_246),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_216),
.C(n_217),
.Y(n_240)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_241),
.B2(n_254),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_242),
.C(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_226),
.C(n_234),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_230),
.C(n_233),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_232),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_238),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_253),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_251),
.C(n_253),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_287),
.B2(n_288),
.Y(n_256)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_278),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_278),
.C(n_287),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_268),
.C(n_269),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_277),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_270),
.Y(n_277)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_274),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_273),
.B(n_296),
.C(n_299),
.Y(n_343)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_281),
.C(n_282),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_293),
.C(n_320),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_307),
.B2(n_320),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_301),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_302),
.C(n_303),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_303),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.CI(n_306),
.CON(n_303),
.SN(n_303)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_305),
.C(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_310),
.C(n_311),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_319),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_314),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_315),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_316),
.A2(n_317),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_342),
.C(n_343),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_344),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_335),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_335),
.C(n_344),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_330),
.C(n_331),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_331),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.CI(n_334),
.CON(n_331),
.SN(n_331)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_333),
.C(n_334),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_338),
.C(n_339),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_341),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_349),
.C(n_359),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_358),
.B2(n_359),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_356),
.C(n_357),
.Y(n_370)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_362),
.C(n_365),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_368)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_369),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_371),
.C(n_375),
.Y(n_376)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);


endmodule