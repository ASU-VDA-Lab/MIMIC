module fake_jpeg_310_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_52),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_46),
.B(n_48),
.C(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_56),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_47),
.B1(n_41),
.B2(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_54),
.B1(n_53),
.B2(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_77),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_45),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_0),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_1),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_16),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_97),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_45),
.C(n_40),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_45),
.B1(n_43),
.B2(n_18),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_12),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_80),
.B(n_43),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_13),
.B(n_37),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_83),
.B1(n_14),
.B2(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_112),
.B1(n_8),
.B2(n_10),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_113),
.C(n_26),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_3),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_111),
.B(n_7),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_4),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_6),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_23),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_92),
.C(n_9),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_121),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_103),
.B(n_100),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_8),
.B(n_10),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_38),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_120),
.B1(n_123),
.B2(n_115),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_118),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_136)
);

OAI21x1_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_134),
.B(n_133),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_127),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_122),
.B1(n_21),
.B2(n_27),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_11),
.B(n_30),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_33),
.C(n_35),
.Y(n_145)
);


endmodule