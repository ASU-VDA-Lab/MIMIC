module fake_jpeg_8198_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_1),
.C(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_59),
.B1(n_20),
.B2(n_17),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_27),
.B(n_21),
.Y(n_76)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_62),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_42),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_63),
.B(n_90),
.C(n_25),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_42),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_89),
.Y(n_120)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_74),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_33),
.B1(n_17),
.B2(n_43),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_84),
.B1(n_25),
.B2(n_30),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_39),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_22),
.A3(n_16),
.B1(n_23),
.B2(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

OR2x4_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_43),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_23),
.B(n_18),
.C(n_26),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_33),
.B1(n_20),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_20),
.B1(n_37),
.B2(n_23),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_40),
.B1(n_34),
.B2(n_27),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_39),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_39),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_37),
.B1(n_33),
.B2(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_113),
.B1(n_30),
.B2(n_26),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_41),
.B1(n_80),
.B2(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_14),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_28),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_78),
.C(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_74),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_126),
.C(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_141),
.Y(n_155)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_71),
.B1(n_76),
.B2(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_134),
.B1(n_138),
.B2(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_85),
.B1(n_90),
.B2(n_64),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_95),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_62),
.C(n_75),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_61),
.B1(n_67),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_93),
.B1(n_61),
.B2(n_80),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_30),
.B1(n_18),
.B2(n_28),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_144),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_75),
.B(n_83),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_105),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_87),
.B1(n_69),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_88),
.B1(n_32),
.B2(n_19),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_154),
.Y(n_156)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_32),
.B1(n_19),
.B2(n_28),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_102),
.B1(n_116),
.B2(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_98),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_176),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_109),
.C(n_98),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_174),
.C(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_122),
.B1(n_114),
.B2(n_97),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_181),
.B1(n_187),
.B2(n_184),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_123),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_179),
.B1(n_141),
.B2(n_129),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_102),
.B1(n_116),
.B2(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_115),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_182),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_101),
.B1(n_115),
.B2(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_101),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_184),
.A2(n_153),
.B(n_145),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_127),
.C(n_154),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_10),
.C(n_13),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_88),
.B1(n_32),
.B2(n_19),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_188),
.A2(n_197),
.B1(n_200),
.B2(n_202),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_136),
.B(n_137),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_160),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_191),
.B(n_192),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_1),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_150),
.B(n_147),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_205),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_151),
.B1(n_143),
.B2(n_32),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_29),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_199),
.C(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_200)
);

NAND2x1_ASAP7_75t_SL g201 ( 
.A(n_164),
.B(n_29),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_201),
.B(n_155),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_29),
.B(n_3),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_29),
.B1(n_4),
.B2(n_5),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_207),
.B1(n_187),
.B2(n_158),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_9),
.B(n_14),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_156),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_163),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_5),
.C(n_6),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_214),
.C(n_217),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_10),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_10),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_165),
.B1(n_168),
.B2(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_179),
.B1(n_178),
.B2(n_161),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_221),
.A2(n_202),
.B1(n_160),
.B2(n_201),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_167),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_234),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_206),
.B(n_158),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_240),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_162),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_195),
.C(n_215),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_244),
.B(n_220),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_190),
.B(n_193),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_195),
.C(n_198),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_226),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_217),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_214),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_194),
.B1(n_161),
.B2(n_173),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_260),
.B1(n_221),
.B2(n_219),
.Y(n_265)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_232),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_218),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_238),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_173),
.B1(n_159),
.B2(n_185),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_235),
.B1(n_227),
.B2(n_231),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_270),
.B1(n_258),
.B2(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_230),
.B1(n_222),
.B2(n_233),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_228),
.B1(n_219),
.B2(n_226),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_274),
.C(n_247),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_186),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_275),
.B(n_157),
.Y(n_281)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_253),
.B1(n_157),
.B2(n_213),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_290),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_287),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.C(n_289),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_245),
.C(n_241),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_264),
.B1(n_260),
.B2(n_270),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_249),
.B(n_244),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_277),
.B(n_280),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_251),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_267),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_286),
.C(n_11),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_282),
.B1(n_286),
.B2(n_289),
.C(n_12),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_272),
.B(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_209),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_171),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_263),
.C(n_248),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_263),
.C(n_6),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_9),
.Y(n_304)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_306),
.Y(n_311)
);

AOI21x1_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_15),
.B(n_6),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_13),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_292),
.B(n_301),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_303),
.B(n_310),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_302),
.A3(n_313),
.B1(n_315),
.B2(n_298),
.C(n_311),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_300),
.B1(n_7),
.B2(n_8),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_7),
.Y(n_321)
);


endmodule