module fake_jpeg_170_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_21),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_44),
.C(n_41),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_47),
.C(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_35),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_75),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_38),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_36),
.B1(n_49),
.B2(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_3),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_56),
.B1(n_62),
.B2(n_58),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_88),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_59),
.B1(n_54),
.B2(n_48),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_19),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_7),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_97),
.B1(n_84),
.B2(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_11),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_98),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_105),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_86),
.B(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_106),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_88),
.B(n_26),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_12),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_110),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_104),
.C(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_102),
.Y(n_117)
);

OAI21x1_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_118),
.B(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_97),
.B1(n_90),
.B2(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_113),
.B1(n_115),
.B2(n_111),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_120),
.A3(n_103),
.B1(n_17),
.B2(n_18),
.C1(n_20),
.C2(n_22),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_28),
.B(n_32),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_27),
.A3(n_31),
.B1(n_24),
.B2(n_25),
.C(n_33),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_29),
.Y(n_125)
);


endmodule