module fake_jpeg_6406_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_20),
.B1(n_32),
.B2(n_17),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_16),
.B1(n_17),
.B2(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_16),
.B1(n_17),
.B2(n_28),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_25),
.B1(n_33),
.B2(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_69),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_33),
.B1(n_30),
.B2(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_73),
.Y(n_120)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_42),
.B(n_38),
.C(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_96),
.Y(n_103)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_80),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_89),
.B1(n_99),
.B2(n_34),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_94),
.Y(n_122)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_93),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

OR2x4_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_43),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_60),
.B(n_59),
.C(n_39),
.Y(n_105)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_43),
.B1(n_64),
.B2(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_27),
.B1(n_34),
.B2(n_19),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_27),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_78),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_50),
.B1(n_54),
.B2(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_82),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_115),
.B(n_26),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_93),
.B(n_71),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_126),
.B(n_74),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_42),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_61),
.CI(n_68),
.CON(n_117),
.SN(n_117)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_77),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_50),
.B1(n_46),
.B2(n_45),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_85),
.B1(n_79),
.B2(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_105),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_36),
.B(n_19),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_129),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_131),
.A2(n_136),
.B(n_110),
.Y(n_176)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_133),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_137),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_70),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_157),
.C(n_121),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_46),
.B1(n_45),
.B2(n_41),
.Y(n_136)
);

AOI22x1_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_45),
.B1(n_46),
.B2(n_41),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_46),
.B1(n_92),
.B2(n_27),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_19),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_142),
.A2(n_150),
.B(n_22),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_65),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_149),
.B1(n_154),
.B2(n_113),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_65),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_92),
.B1(n_21),
.B2(n_90),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_26),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_21),
.B1(n_52),
.B2(n_26),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_155),
.B1(n_159),
.B2(n_102),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_65),
.Y(n_153)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_103),
.A2(n_52),
.B1(n_21),
.B2(n_23),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_122),
.B(n_115),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_52),
.C(n_26),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_23),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_158),
.Y(n_168)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_122),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_178),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_165),
.B(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_10),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_179),
.B1(n_181),
.B2(n_100),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_126),
.B(n_120),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_174),
.B(n_176),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_177),
.C(n_190),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_125),
.B(n_117),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_143),
.C(n_146),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_117),
.B(n_128),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_127),
.B1(n_102),
.B2(n_110),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_123),
.B1(n_111),
.B2(n_127),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_152),
.B1(n_134),
.B2(n_142),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_102),
.B1(n_111),
.B2(n_100),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_22),
.A3(n_23),
.B1(n_52),
.B2(n_3),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_0),
.B(n_1),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_193),
.B(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_144),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_116),
.C(n_100),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_116),
.C(n_23),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_149),
.B1(n_151),
.B2(n_155),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_161),
.B1(n_183),
.B2(n_193),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_216),
.B1(n_221),
.B2(n_182),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_207),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_2),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_218),
.B(n_219),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_215),
.B1(n_220),
.B2(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_173),
.C(n_188),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_116),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_180),
.B1(n_189),
.B2(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_164),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_228),
.C(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_160),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_6),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_186),
.C(n_178),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_220),
.C(n_194),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_167),
.B1(n_161),
.B2(n_186),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_170),
.C(n_187),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_239),
.C(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_216),
.C(n_214),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_184),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_15),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_8),
.C(n_9),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

AO22x1_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_210),
.B1(n_205),
.B2(n_197),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_248),
.A2(n_204),
.B1(n_209),
.B2(n_212),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_207),
.B(n_203),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_223),
.B(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_15),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_241),
.B1(n_246),
.B2(n_235),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_11),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_231),
.B1(n_248),
.B2(n_232),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_11),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_269),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_11),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_241),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_226),
.B(n_9),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_249),
.C(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_273),
.C(n_269),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_249),
.C(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_239),
.B1(n_238),
.B2(n_228),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_278),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_254),
.C(n_261),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_234),
.B(n_240),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_251),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_303)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_279),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_298),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_287),
.A2(n_266),
.B1(n_264),
.B2(n_251),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_296),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_268),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_253),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_301),
.C(n_302),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_243),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_284),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_264),
.C(n_250),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_6),
.C(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_300),
.A2(n_286),
.B1(n_281),
.B2(n_278),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_306),
.B(n_312),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_275),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_311),
.B(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_7),
.C(n_9),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_12),
.C(n_13),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_14),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_12),
.C(n_13),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_12),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_313),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_305),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_328),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_314),
.C(n_307),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_14),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_327),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_324),
.B(n_329),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_331),
.B(n_333),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_324),
.Y(n_338)
);


endmodule