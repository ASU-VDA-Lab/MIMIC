module real_aes_939_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_512, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_512;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g264 ( .A(n_0), .B(n_188), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_1), .A2(n_62), .B1(n_85), .B2(n_102), .Y(n_84) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_2), .A2(n_51), .B1(n_89), .B2(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g162 ( .A(n_3), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_4), .B(n_194), .Y(n_207) );
NAND2xp33_ASAP7_75t_SL g256 ( .A(n_5), .B(n_192), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_6), .A2(n_67), .B1(n_113), .B2(n_115), .Y(n_112) );
INVx1_ASAP7_75t_L g239 ( .A(n_7), .Y(n_239) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_8), .A2(n_19), .B1(n_89), .B2(n_90), .Y(n_88) );
AND2x2_ASAP7_75t_L g205 ( .A(n_9), .B(n_198), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_10), .A2(n_55), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx2_ASAP7_75t_L g199 ( .A(n_11), .Y(n_199) );
AOI221x1_ASAP7_75t_L g250 ( .A1(n_12), .A2(n_177), .B1(n_251), .B2(n_253), .C(n_255), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_13), .A2(n_144), .B1(n_145), .B2(n_148), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_13), .B(n_194), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_14), .A2(n_48), .B1(n_137), .B2(n_138), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_15), .A2(n_177), .B(n_209), .Y(n_208) );
AOI221xp5_ASAP7_75t_SL g219 ( .A1(n_16), .A2(n_29), .B1(n_177), .B2(n_194), .C(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g493 ( .A(n_16), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_17), .B(n_188), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_18), .A2(n_35), .B1(n_118), .B2(n_121), .Y(n_117) );
OAI221xp5_ASAP7_75t_L g154 ( .A1(n_19), .A2(n_51), .B1(n_53), .B2(n_155), .C(n_157), .Y(n_154) );
OR2x2_ASAP7_75t_L g200 ( .A(n_20), .B(n_65), .Y(n_200) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_20), .A2(n_65), .B(n_199), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_21), .B(n_184), .Y(n_231) );
INVxp67_ASAP7_75t_L g249 ( .A(n_22), .Y(n_249) );
AND2x2_ASAP7_75t_L g280 ( .A(n_23), .B(n_197), .Y(n_280) );
INVx3_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_25), .A2(n_177), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_26), .B(n_184), .Y(n_221) );
INVx1_ASAP7_75t_SL g100 ( .A(n_27), .Y(n_100) );
INVx1_ASAP7_75t_L g164 ( .A(n_28), .Y(n_164) );
AND2x2_ASAP7_75t_L g178 ( .A(n_28), .B(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g192 ( .A(n_28), .B(n_162), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_30), .A2(n_58), .B1(n_177), .B2(n_244), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_31), .B(n_188), .Y(n_278) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_32), .A2(n_53), .B1(n_89), .B2(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g267 ( .A(n_33), .B(n_197), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_34), .B(n_197), .Y(n_223) );
INVx1_ASAP7_75t_L g181 ( .A(n_36), .Y(n_181) );
INVx1_ASAP7_75t_L g190 ( .A(n_36), .Y(n_190) );
INVx1_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_38), .B(n_194), .Y(n_279) );
AND2x2_ASAP7_75t_L g201 ( .A(n_39), .B(n_197), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_40), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_41), .B(n_184), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_42), .B(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_43), .B(n_198), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_44), .A2(n_177), .B(n_276), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_45), .A2(n_68), .B1(n_146), .B2(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_45), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_46), .B(n_184), .Y(n_211) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_47), .B(n_232), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_49), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_49), .B(n_80), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_50), .A2(n_80), .B1(n_81), .B2(n_141), .Y(n_79) );
INVx1_ASAP7_75t_L g141 ( .A(n_50), .Y(n_141) );
INVxp33_ASAP7_75t_L g159 ( .A(n_51), .Y(n_159) );
INVx1_ASAP7_75t_L g179 ( .A(n_52), .Y(n_179) );
INVx1_ASAP7_75t_L g186 ( .A(n_52), .Y(n_186) );
INVxp67_ASAP7_75t_L g158 ( .A(n_53), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_54), .A2(n_63), .B1(n_129), .B2(n_130), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_56), .B(n_194), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_57), .A2(n_59), .B1(n_194), .B2(n_240), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_60), .B(n_188), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_61), .B(n_188), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_64), .A2(n_177), .B(n_182), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_66), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g147 ( .A(n_68), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_69), .A2(n_75), .B1(n_133), .B2(n_134), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_70), .A2(n_143), .B1(n_149), .B2(n_150), .Y(n_142) );
INVx1_ASAP7_75t_L g149 ( .A(n_70), .Y(n_149) );
INVxp67_ASAP7_75t_L g252 ( .A(n_71), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_72), .B(n_194), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_73), .B(n_184), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_74), .A2(n_177), .B(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_SL g156 ( .A(n_76), .Y(n_156) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_151), .B1(n_165), .B2(n_489), .C(n_490), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_142), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_80), .A2(n_81), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_81), .B(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp67_ASAP7_75t_L g82 ( .A(n_83), .B(n_122), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_107), .C(n_112), .D(n_117), .Y(n_83) );
AND2x6_ASAP7_75t_L g85 ( .A(n_86), .B(n_94), .Y(n_85) );
AND2x2_ASAP7_75t_L g113 ( .A(n_86), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g120 ( .A(n_86), .B(n_103), .Y(n_120) );
AND2x2_ASAP7_75t_L g126 ( .A(n_86), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g86 ( .A(n_87), .B(n_91), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g106 ( .A(n_88), .Y(n_106) );
AND2x2_ASAP7_75t_L g111 ( .A(n_88), .B(n_92), .Y(n_111) );
AND2x4_ASAP7_75t_L g116 ( .A(n_88), .B(n_91), .Y(n_116) );
INVx2_ASAP7_75t_L g90 ( .A(n_89), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_89), .Y(n_96) );
OAI22x1_ASAP7_75t_L g98 ( .A1(n_89), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
INVxp67_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g105 ( .A(n_92), .B(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g108 ( .A(n_94), .B(n_105), .Y(n_108) );
AND2x2_ASAP7_75t_L g133 ( .A(n_94), .B(n_116), .Y(n_133) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_97), .Y(n_94) );
INVx2_ASAP7_75t_L g104 ( .A(n_95), .Y(n_104) );
BUFx2_ASAP7_75t_L g110 ( .A(n_95), .Y(n_110) );
AND2x2_ASAP7_75t_L g127 ( .A(n_95), .B(n_98), .Y(n_127) );
AND2x4_ASAP7_75t_L g103 ( .A(n_97), .B(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g114 ( .A(n_98), .B(n_104), .Y(n_114) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
AND2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
AND2x2_ASAP7_75t_L g115 ( .A(n_103), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g121 ( .A(n_103), .B(n_111), .Y(n_121) );
AND2x4_ASAP7_75t_L g137 ( .A(n_105), .B(n_114), .Y(n_137) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_106), .Y(n_140) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_111), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g129 ( .A(n_114), .B(n_116), .Y(n_129) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx8_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND4xp25_ASAP7_75t_SL g122 ( .A(n_123), .B(n_128), .C(n_132), .D(n_136), .Y(n_122) );
INVx4_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx6_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g134 ( .A(n_127), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g138 ( .A(n_127), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_143), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_153), .Y(n_152) );
AND3x1_ASAP7_75t_SL g153 ( .A(n_154), .B(n_160), .C(n_163), .Y(n_153) );
INVxp67_ASAP7_75t_L g498 ( .A(n_154), .Y(n_498) );
CKINVDCx8_ASAP7_75t_R g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_160), .Y(n_496) );
AO21x1_ASAP7_75t_SL g508 ( .A1(n_160), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g241 ( .A(n_161), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_SL g505 ( .A(n_161), .B(n_163), .Y(n_505) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g180 ( .A(n_162), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_163), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2x1p5_ASAP7_75t_L g245 ( .A(n_164), .B(n_246), .Y(n_245) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_428), .Y(n_166) );
NOR3xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_321), .C(n_372), .Y(n_167) );
OAI211xp5_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_213), .B(n_268), .C(n_299), .Y(n_168) );
INVxp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_202), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_173), .B(n_273), .Y(n_436) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g281 ( .A(n_174), .B(n_204), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_174), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g298 ( .A(n_174), .B(n_288), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_174), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g335 ( .A(n_174), .B(n_311), .Y(n_335) );
INVx2_ASAP7_75t_L g361 ( .A(n_174), .Y(n_361) );
AND2x4_ASAP7_75t_L g370 ( .A(n_174), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g475 ( .A(n_174), .B(n_342), .Y(n_475) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_196), .B(n_201), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_193), .Y(n_175) );
AND2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
BUFx3_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
AND2x6_ASAP7_75t_L g188 ( .A(n_179), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g247 ( .A(n_179), .Y(n_247) );
AND2x4_ASAP7_75t_L g244 ( .A(n_180), .B(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g184 ( .A(n_181), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_187), .B(n_191), .Y(n_182) );
AND2x4_ASAP7_75t_L g195 ( .A(n_185), .B(n_189), .Y(n_195) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_191), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_191), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_191), .A2(n_264), .B(n_265), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_191), .A2(n_277), .B(n_278), .Y(n_276) );
INVx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x4_ASAP7_75t_L g194 ( .A(n_192), .B(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_194), .Y(n_489) );
INVx1_ASAP7_75t_L g257 ( .A(n_195), .Y(n_257) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_196), .A2(n_274), .B(n_280), .Y(n_273) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_196), .A2(n_274), .B(n_280), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_197), .Y(n_196) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_197), .A2(n_219), .B(n_223), .Y(n_218) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AND2x4_ASAP7_75t_L g212 ( .A(n_199), .B(n_200), .Y(n_212) );
AND2x2_ASAP7_75t_L g359 ( .A(n_202), .B(n_360), .Y(n_359) );
OAI32xp33_ASAP7_75t_L g442 ( .A1(n_202), .A2(n_364), .A3(n_368), .B1(n_375), .B2(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_202), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_297), .Y(n_296) );
NAND3xp33_ASAP7_75t_L g369 ( .A(n_203), .B(n_291), .C(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g395 ( .A(n_203), .B(n_298), .Y(n_395) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_204), .Y(n_285) );
INVx5_ASAP7_75t_L g320 ( .A(n_204), .Y(n_320) );
AND2x4_ASAP7_75t_L g376 ( .A(n_204), .B(n_288), .Y(n_376) );
OR2x2_ASAP7_75t_L g391 ( .A(n_204), .B(n_311), .Y(n_391) );
OR2x2_ASAP7_75t_L g417 ( .A(n_204), .B(n_273), .Y(n_417) );
AND2x2_ASAP7_75t_L g425 ( .A(n_204), .B(n_371), .Y(n_425) );
AND2x4_ASAP7_75t_SL g450 ( .A(n_204), .B(n_370), .Y(n_450) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_212), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_212), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_212), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_212), .B(n_252), .Y(n_251) );
NOR3xp33_ASAP7_75t_L g255 ( .A(n_212), .B(n_256), .C(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_214), .B(n_370), .Y(n_446) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_215), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x6_ASAP7_75t_SL g270 ( .A(n_216), .B(n_271), .Y(n_270) );
INVxp67_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g295 ( .A(n_217), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_217), .B(n_330), .Y(n_348) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_217), .Y(n_486) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
AND2x2_ASAP7_75t_L g328 ( .A(n_218), .B(n_259), .Y(n_328) );
INVx2_ASAP7_75t_L g356 ( .A(n_218), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_218), .B(n_225), .Y(n_397) );
BUFx3_ASAP7_75t_L g421 ( .A(n_218), .Y(n_421) );
OR2x2_ASAP7_75t_L g433 ( .A(n_218), .B(n_225), .Y(n_433) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_218), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_224), .A2(n_464), .B1(n_467), .B2(n_468), .Y(n_463) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
INVx1_ASAP7_75t_L g291 ( .A(n_225), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_225), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g309 ( .A(n_225), .Y(n_309) );
AND2x4_ASAP7_75t_SL g326 ( .A(n_225), .B(n_236), .Y(n_326) );
AND2x4_ASAP7_75t_L g331 ( .A(n_225), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g340 ( .A(n_225), .Y(n_340) );
OR2x2_ASAP7_75t_L g346 ( .A(n_225), .B(n_236), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_225), .B(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_225), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_225), .B(n_328), .Y(n_462) );
OR2x2_ASAP7_75t_L g478 ( .A(n_225), .B(n_381), .Y(n_478) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_234), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_232), .Y(n_226) );
INVx2_ASAP7_75t_SL g313 ( .A(n_232), .Y(n_313) );
BUFx4f_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_235), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g304 ( .A(n_235), .Y(n_304) );
AND2x2_ASAP7_75t_SL g411 ( .A(n_235), .B(n_295), .Y(n_411) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_258), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_236), .B(n_259), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_236), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_236), .B(n_303), .Y(n_307) );
INVx3_ASAP7_75t_L g332 ( .A(n_236), .Y(n_332) );
INVx1_ASAP7_75t_L g365 ( .A(n_236), .Y(n_365) );
AND2x2_ASAP7_75t_L g445 ( .A(n_236), .B(n_309), .Y(n_445) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B1(n_244), .B2(n_248), .Y(n_237) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_242), .Y(n_510) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_245), .Y(n_509) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx4_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AOI21x1_ASAP7_75t_L g260 ( .A1(n_254), .A2(n_261), .B(n_267), .Y(n_260) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_259), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g330 ( .A(n_259), .Y(n_330) );
AND2x2_ASAP7_75t_L g355 ( .A(n_259), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g381 ( .A(n_259), .B(n_303), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_259), .B(n_332), .Y(n_398) );
INVx1_ASAP7_75t_L g404 ( .A(n_259), .Y(n_404) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_266), .Y(n_261) );
AOI222xp33_ASAP7_75t_SL g268 ( .A1(n_269), .A2(n_272), .B1(n_282), .B2(n_289), .C1(n_292), .C2(n_296), .Y(n_268) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_281), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_273), .B(n_342), .Y(n_393) );
AND2x4_ASAP7_75t_L g409 ( .A(n_273), .B(n_320), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_279), .Y(n_274) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g334 ( .A(n_285), .B(n_335), .Y(n_334) );
AOI222xp33_ASAP7_75t_L g299 ( .A1(n_286), .A2(n_300), .B1(n_305), .B2(n_310), .C1(n_318), .C2(n_512), .Y(n_299) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g438 ( .A(n_287), .B(n_342), .Y(n_438) );
OR2x2_ASAP7_75t_L g481 ( .A(n_287), .B(n_387), .Y(n_481) );
AND2x2_ASAP7_75t_L g310 ( .A(n_288), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g371 ( .A(n_288), .Y(n_371) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_288), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_289), .A2(n_400), .B(n_405), .C(n_406), .Y(n_399) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g427 ( .A(n_291), .Y(n_427) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
AND2x2_ASAP7_75t_L g341 ( .A(n_297), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g350 ( .A(n_297), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI31xp33_ASAP7_75t_L g392 ( .A1(n_300), .A2(n_318), .A3(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g394 ( .A1(n_301), .A2(n_351), .B(n_395), .C(n_396), .Y(n_394) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
OR2x2_ASAP7_75t_L g383 ( .A(n_302), .B(n_332), .Y(n_383) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
BUFx2_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
AND2x2_ASAP7_75t_L g360 ( .A(n_311), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
AOI21x1_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_317), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_320), .B(n_377), .Y(n_469) );
OAI211xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_333), .B(n_336), .C(n_358), .Y(n_321) );
INVxp33_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_324), .B(n_329), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g362 ( .A(n_326), .B(n_355), .Y(n_362) );
OR2x2_ASAP7_75t_L g338 ( .A(n_327), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g368 ( .A(n_327), .B(n_342), .Y(n_368) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g444 ( .A(n_328), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g467 ( .A(n_329), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_331), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_331), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g479 ( .A(n_331), .B(n_355), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_331), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g422 ( .A(n_332), .B(n_404), .Y(n_422) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AOI322xp5_ASAP7_75t_L g476 ( .A1(n_335), .A2(n_355), .A3(n_409), .B1(n_434), .B2(n_477), .C1(n_479), .C2(n_480), .Y(n_476) );
AOI211xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_341), .B(n_343), .C(n_352), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_339), .B(n_367), .Y(n_389) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g354 ( .A(n_340), .B(n_355), .Y(n_354) );
NOR2x1p5_ASAP7_75t_L g420 ( .A(n_340), .B(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_340), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_341), .A2(n_359), .B(n_362), .C(n_363), .Y(n_358) );
AND2x4_ASAP7_75t_L g377 ( .A(n_342), .B(n_361), .Y(n_377) );
INVx2_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_342), .B(n_376), .Y(n_407) );
AND2x2_ASAP7_75t_L g449 ( .A(n_342), .B(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_342), .B(n_466), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_342), .B(n_370), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_349), .Y(n_343) );
AND2x2_ASAP7_75t_L g439 ( .A(n_345), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g367 ( .A(n_348), .Y(n_367) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_357), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_360), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g454 ( .A(n_360), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_366), .B(n_368), .C(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_367), .Y(n_451) );
INVx3_ASAP7_75t_SL g466 ( .A(n_370), .Y(n_466) );
NAND5xp2_ASAP7_75t_L g372 ( .A(n_373), .B(n_392), .C(n_399), .D(n_412), .E(n_423), .Y(n_372) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_382), .B2(n_384), .C1(n_388), .C2(n_390), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_375), .A2(n_456), .B1(n_460), .B2(n_461), .Y(n_455) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g405 ( .A(n_376), .B(n_377), .Y(n_405) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_386), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_387), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g424 ( .A(n_387), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g435 ( .A(n_387), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g465 ( .A(n_391), .B(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_410), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_409), .A2(n_413), .B1(n_414), .B2(n_418), .Y(n_412) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_409), .Y(n_460) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g426 ( .A(n_411), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g431 ( .A(n_413), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_SL g459 ( .A(n_422), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_447), .C(n_470), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_430), .B(n_446), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B1(n_437), .B2(n_439), .C(n_442), .Y(n_430) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_459), .Y(n_471) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
OAI321xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .A3(n_452), .B1(n_454), .B2(n_455), .C(n_463), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_461), .A2(n_483), .B1(n_487), .B2(n_488), .Y(n_482) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_472), .B(n_476), .C(n_482), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_493), .B1(n_494), .B2(n_499), .C1(n_503), .C2(n_506), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
endmodule