module fake_jpeg_19060_n_343 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_19),
.B1(n_35),
.B2(n_22),
.Y(n_71)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_36),
.B1(n_19),
.B2(n_35),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_69),
.B1(n_47),
.B2(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_39),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_36),
.B1(n_27),
.B2(n_28),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_71),
.B1(n_22),
.B2(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_36),
.B1(n_19),
.B2(n_35),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_29),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_43),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_39),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_94),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_90),
.B1(n_47),
.B2(n_44),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_49),
.B1(n_28),
.B2(n_38),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_91),
.B1(n_51),
.B2(n_41),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_49),
.B1(n_28),
.B2(n_38),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_100),
.B1(n_59),
.B2(n_44),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_43),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_39),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_81),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_117),
.B1(n_127),
.B2(n_134),
.Y(n_136)
);

NOR4xp25_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_96),
.C(n_90),
.D(n_102),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_86),
.B1(n_100),
.B2(n_97),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_47),
.B1(n_44),
.B2(n_49),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_24),
.B(n_22),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_133),
.B1(n_20),
.B2(n_26),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_125),
.B1(n_92),
.B2(n_34),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_34),
.B1(n_27),
.B2(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_41),
.B1(n_51),
.B2(n_18),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_41),
.B1(n_51),
.B2(n_42),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_143),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_87),
.C(n_75),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_156),
.C(n_131),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_145),
.B(n_153),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_74),
.B1(n_73),
.B2(n_86),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_151),
.B1(n_160),
.B2(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_152),
.B1(n_134),
.B2(n_111),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_42),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_120),
.B1(n_105),
.B2(n_117),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_97),
.B1(n_42),
.B2(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_39),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_81),
.C(n_29),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_29),
.Y(n_168)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_89),
.B1(n_20),
.B2(n_32),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_166),
.B1(n_136),
.B2(n_139),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_125),
.B(n_128),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_140),
.B(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_173),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_172),
.B1(n_148),
.B2(n_152),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_111),
.B1(n_119),
.B2(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_188),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_132),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_122),
.C(n_132),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_177),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_136),
.B1(n_151),
.B2(n_135),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_25),
.C(n_26),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_180),
.B(n_38),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_186),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_114),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_25),
.C(n_9),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_107),
.B(n_114),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_182),
.B(n_141),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_138),
.A2(n_106),
.B(n_31),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_187),
.C(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_130),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_189),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_200),
.B1(n_211),
.B2(n_217),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_214),
.C(n_29),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_195),
.Y(n_227)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_155),
.B(n_143),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_165),
.B1(n_167),
.B2(n_161),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_209),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_184),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_150),
.B(n_154),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_182),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_172),
.A2(n_130),
.B1(n_118),
.B2(n_131),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_167),
.B(n_131),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_118),
.C(n_29),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_215),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_163),
.A2(n_33),
.B(n_31),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_0),
.B(n_1),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_185),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_222),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_190),
.B1(n_215),
.B2(n_211),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_187),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_171),
.Y(n_224)
);

OAI322xp33_ASAP7_75t_L g267 ( 
.A1(n_224),
.A2(n_217),
.A3(n_194),
.B1(n_21),
.B2(n_33),
.C1(n_30),
.C2(n_8),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_178),
.B(n_183),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_228),
.C(n_240),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_205),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_203),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_21),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_243),
.C(n_202),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_21),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_209),
.B(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_256),
.B1(n_257),
.B2(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_213),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_263),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_208),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_225),
.B(n_199),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_216),
.B(n_219),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_204),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_230),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

OAI22x1_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_241),
.B1(n_234),
.B2(n_221),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_271),
.A2(n_254),
.B1(n_252),
.B2(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_228),
.C(n_226),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_280),
.C(n_257),
.Y(n_294)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_220),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_279),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_224),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_222),
.C(n_243),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_240),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_246),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_290),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_259),
.C(n_258),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_248),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_262),
.B1(n_261),
.B2(n_260),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_298),
.B1(n_2),
.B2(n_17),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_256),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_253),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_236),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_11),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_229),
.B1(n_232),
.B2(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_300),
.B1(n_278),
.B2(n_273),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_284),
.B(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_312),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_281),
.B1(n_3),
.B2(n_4),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_306),
.A2(n_314),
.B1(n_10),
.B2(n_7),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_11),
.CI(n_3),
.CON(n_307),
.SN(n_307)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_14),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_12),
.C(n_5),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_287),
.C(n_7),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_294),
.A2(n_13),
.B1(n_7),
.B2(n_8),
.Y(n_314)
);

NAND2x1p5_ASAP7_75t_R g315 ( 
.A(n_310),
.B(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_293),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_320),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_14),
.B(n_8),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_314),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_302),
.C(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_329),
.Y(n_334)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_302),
.C(n_303),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_326),
.B1(n_316),
.B2(n_315),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_331),
.B(n_333),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_303),
.B(n_307),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_327),
.C(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_332),
.Y(n_337)
);

OAI311xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_336),
.A3(n_9),
.B1(n_10),
.C1(n_15),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_17),
.B(n_10),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_15),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_16),
.B(n_2),
.Y(n_343)
);


endmodule