module fake_jpeg_12363_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_51),
.B(n_68),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g152 ( 
.A(n_52),
.Y(n_152)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_45),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_12),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_18),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_48),
.B1(n_27),
.B2(n_44),
.Y(n_111)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_12),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_80),
.B(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_9),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_9),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_111),
.A2(n_22),
.B1(n_40),
.B2(n_18),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_52),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_113),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_48),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_119),
.B(n_123),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_30),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_27),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_44),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_36),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_52),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_60),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_46),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_58),
.B(n_36),
.Y(n_151)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_49),
.Y(n_154)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_174),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_33),
.B1(n_19),
.B2(n_39),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_98),
.B1(n_74),
.B2(n_56),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_162),
.A2(n_172),
.B1(n_173),
.B2(n_71),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_40),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_163),
.B(n_175),
.Y(n_229)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

INVx5_ASAP7_75t_SL g165 ( 
.A(n_155),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_165),
.Y(n_212)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_101),
.A2(n_75),
.B1(n_89),
.B2(n_55),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_38),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_32),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_190),
.C(n_199),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_116),
.A2(n_61),
.B1(n_59),
.B2(n_70),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_121),
.B1(n_153),
.B2(n_144),
.Y(n_223)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_33),
.B1(n_39),
.B2(n_62),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_65),
.B1(n_76),
.B2(n_83),
.Y(n_214)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_34),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_131),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_195),
.Y(n_213)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_32),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_131),
.B(n_34),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_194),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_34),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_134),
.B1(n_132),
.B2(n_106),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_117),
.B(n_38),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_22),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_146),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_179),
.C(n_199),
.Y(n_240)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_206),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_214),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_158),
.B(n_117),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_224),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_201),
.B1(n_200),
.B2(n_202),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_159),
.A2(n_132),
.B1(n_134),
.B2(n_106),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_155),
.B1(n_188),
.B2(n_104),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_127),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_213),
.Y(n_274)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_169),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_248),
.B(n_264),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_165),
.B(n_190),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_249),
.A2(n_261),
.B(n_237),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_266),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_174),
.B1(n_104),
.B2(n_146),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_158),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_169),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_253),
.B(n_254),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_163),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_205),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_259),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_189),
.B1(n_191),
.B2(n_187),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_262),
.A2(n_279),
.B1(n_221),
.B2(n_217),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_240),
.B(n_171),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_263),
.B(n_267),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_232),
.B(n_170),
.Y(n_264)
);

AO21x1_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_223),
.B(n_196),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_226),
.B(n_237),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_177),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_186),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_270),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_213),
.B(n_178),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_213),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_276),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_221),
.B1(n_217),
.B2(n_222),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_197),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_273),
.B(n_238),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_230),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_212),
.B1(n_206),
.B2(n_230),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_231),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_212),
.B1(n_243),
.B2(n_164),
.Y(n_284)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_129),
.B1(n_116),
.B2(n_144),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_224),
.B(n_215),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_280),
.A2(n_314),
.B(n_277),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_283),
.A2(n_290),
.B(n_294),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_289),
.B1(n_291),
.B2(n_261),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_298),
.C(n_299),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_212),
.B1(n_237),
.B2(n_230),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_274),
.B(n_181),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_307),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_222),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_252),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_305),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_262),
.A2(n_129),
.B1(n_125),
.B2(n_127),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_245),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_250),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_193),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_313),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_258),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_245),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_278),
.Y(n_328)
);

XOR2x2_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_96),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_260),
.A2(n_234),
.B(n_241),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_317),
.B(n_319),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_246),
.C(n_272),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_333),
.C(n_310),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_312),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_324),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_264),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_303),
.B(n_248),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_331),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_265),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_238),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_334),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_272),
.C(n_275),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_247),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_336),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_285),
.Y(n_336)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_279),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_339),
.Y(n_367)
);

AO22x1_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_276),
.B1(n_257),
.B2(n_256),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_283),
.A2(n_288),
.B1(n_282),
.B2(n_291),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_341),
.A2(n_288),
.B1(n_314),
.B2(n_290),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_298),
.B(n_247),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_342),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_304),
.A2(n_276),
.B1(n_235),
.B2(n_269),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_345),
.B1(n_301),
.B2(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_346),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_288),
.A2(n_235),
.B1(n_269),
.B2(n_210),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_168),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_348),
.Y(n_366)
);

NOR4xp25_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_296),
.C(n_297),
.D(n_287),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_355),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_351),
.A2(n_339),
.B1(n_333),
.B2(n_337),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_352),
.A2(n_379),
.B1(n_204),
.B2(n_203),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_335),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_334),
.A2(n_302),
.B1(n_293),
.B2(n_286),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_360),
.A2(n_362),
.B1(n_373),
.B2(n_380),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_307),
.C(n_293),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_365),
.C(n_372),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_286),
.B1(n_300),
.B2(n_209),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_300),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_370),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_216),
.C(n_219),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_183),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_219),
.C(n_216),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_348),
.A2(n_210),
.B1(n_176),
.B2(n_125),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_160),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_332),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_315),
.A2(n_122),
.B1(n_153),
.B2(n_193),
.Y(n_377)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_377),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_346),
.A2(n_122),
.B1(n_31),
.B2(n_228),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_234),
.B1(n_241),
.B2(n_228),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_328),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_338),
.B(n_330),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_386),
.A2(n_108),
.B(n_88),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_394),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_344),
.C(n_322),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_395),
.C(n_396),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_316),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_320),
.Y(n_391)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_391),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_363),
.B1(n_359),
.B2(n_379),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_375),
.B(n_327),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_338),
.C(n_318),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_339),
.C(n_343),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_345),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_402),
.Y(n_432)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_365),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_406),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_376),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_411),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_378),
.B(n_259),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_185),
.C(n_166),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_412),
.C(n_397),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_152),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_407),
.A2(n_351),
.B1(n_373),
.B2(n_380),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_152),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_106),
.Y(n_437)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_192),
.C(n_160),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

AOI211xp5_ASAP7_75t_L g417 ( 
.A1(n_386),
.A2(n_408),
.B(n_353),
.C(n_367),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_417),
.A2(n_418),
.B1(n_420),
.B2(n_406),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_407),
.A2(n_363),
.B1(n_353),
.B2(n_367),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_419),
.A2(n_433),
.B1(n_434),
.B2(n_422),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_391),
.A2(n_359),
.B1(n_360),
.B2(n_374),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_403),
.A2(n_362),
.B1(n_368),
.B2(n_354),
.Y(n_426)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_388),
.A2(n_368),
.B1(n_354),
.B2(n_383),
.Y(n_427)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_0),
.Y(n_428)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_428),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_385),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_430),
.A2(n_434),
.B(n_435),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_412),
.Y(n_431)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_410),
.A2(n_18),
.B1(n_43),
.B2(n_31),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_108),
.C(n_31),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_135),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_20),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_384),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_438),
.B(n_413),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_439),
.A2(n_418),
.B1(n_415),
.B2(n_432),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_441),
.B(n_447),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_423),
.B(n_395),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_444),
.B(n_455),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_400),
.C(n_385),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_448),
.Y(n_474)
);

XNOR2x2_ASAP7_75t_SL g446 ( 
.A(n_432),
.B(n_394),
.Y(n_446)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

A2O1A1O1Ixp25_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_413),
.B(n_396),
.C(n_402),
.D(n_392),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_387),
.C(n_409),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_423),
.C(n_421),
.Y(n_462)
);

BUFx12_ASAP7_75t_L g451 ( 
.A(n_420),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_452),
.A2(n_458),
.B1(n_38),
.B2(n_34),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_405),
.Y(n_454)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_454),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_436),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_43),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_459),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_428),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_462),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_452),
.A2(n_419),
.B(n_430),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_461),
.A2(n_470),
.B(n_0),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_429),
.C(n_421),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_468),
.B(n_469),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_465),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_437),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_433),
.C(n_135),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_448),
.A2(n_0),
.B(n_1),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_442),
.A2(n_38),
.B1(n_34),
.B2(n_46),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_477),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_476),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_443),
.A2(n_38),
.B1(n_20),
.B2(n_2),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_450),
.C(n_444),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_480),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_446),
.C(n_440),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_476),
.A2(n_440),
.B1(n_451),
.B2(n_449),
.Y(n_481)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

FAx1_ASAP7_75t_SL g482 ( 
.A(n_474),
.B(n_451),
.CI(n_458),
.CON(n_482),
.SN(n_482)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_488),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_462),
.C(n_468),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_483),
.A2(n_485),
.B(n_486),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_455),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_20),
.C(n_1),
.Y(n_486)
);

HAxp5_ASAP7_75t_SL g487 ( 
.A(n_463),
.B(n_20),
.CON(n_487),
.SN(n_487)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_470),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_0),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_489),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_467),
.B(n_8),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_1),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_477),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_478),
.A2(n_492),
.B(n_483),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_494),
.B(n_501),
.Y(n_509)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_495),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_498),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_461),
.C(n_472),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_493),
.A2(n_469),
.B(n_473),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_489),
.B1(n_486),
.B2(n_487),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_505),
.B(n_499),
.Y(n_506)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_506),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_503),
.A2(n_480),
.B(n_482),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_511),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_502),
.B(n_482),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_SL g514 ( 
.A1(n_508),
.A2(n_496),
.B(n_500),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_479),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_512),
.A2(n_500),
.B(n_472),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_515),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_497),
.C(n_479),
.Y(n_518)
);

AOI322xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_509),
.A3(n_513),
.B1(n_510),
.B2(n_6),
.C1(n_2),
.C2(n_8),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g522 ( 
.A1(n_519),
.A2(n_520),
.B(n_5),
.Y(n_522)
);

AOI321xp33_ASAP7_75t_L g520 ( 
.A1(n_516),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_521),
.C(n_517),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_523),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_5),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_7),
.B1(n_317),
.B2(n_434),
.Y(n_526)
);


endmodule