module fake_jpeg_15118_n_105 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_10),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_4),
.B(n_5),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_20),
.B(n_15),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_17),
.B(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_49),
.B1(n_8),
.B2(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_25),
.A2(n_19),
.B1(n_13),
.B2(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_21),
.B1(n_29),
.B2(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_26),
.A2(n_21),
.B1(n_12),
.B2(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_63),
.B1(n_44),
.B2(n_38),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_65),
.B(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_36),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_61),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_66),
.C(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_72),
.B1(n_56),
.B2(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_48),
.B1(n_42),
.B2(n_40),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_57),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_60),
.B1(n_38),
.B2(n_54),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_54),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_36),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_68),
.B1(n_67),
.B2(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_74),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_80),
.B1(n_86),
.B2(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_83),
.C(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_70),
.B1(n_58),
.B2(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_96),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_87),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_88),
.B(n_91),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_90),
.C(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_47),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_99),
.B(n_96),
.C(n_70),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);


endmodule