module fake_jpeg_7388_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_21),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_10),
.B1(n_16),
.B2(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_22),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_25),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_23),
.B1(n_22),
.B2(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_25),
.B(n_26),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_19),
.B(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_20),
.B1(n_24),
.B2(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_24),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_31),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_52),
.B(n_40),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_24),
.B1(n_35),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_18),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_43),
.C(n_37),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_57),
.B1(n_15),
.B2(n_8),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_40),
.B1(n_17),
.B2(n_9),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_15),
.B1(n_2),
.B2(n_4),
.Y(n_62)
);

AOI321xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_51),
.A3(n_50),
.B1(n_52),
.B2(n_47),
.C(n_18),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_54),
.B(n_53),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_17),
.A3(n_9),
.B1(n_12),
.B2(n_15),
.C1(n_13),
.C2(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_68),
.C(n_65),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_62),
.C(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_1),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_5),
.B(n_6),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_69),
.C(n_5),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_76),
.B1(n_74),
.B2(n_6),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_6),
.Y(n_79)
);


endmodule