module fake_jpeg_14922_n_121 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_1),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_29),
.A2(n_30),
.B1(n_23),
.B2(n_16),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_32),
.B(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_60),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_51),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_17),
.B(n_27),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_8),
.B(n_11),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_3),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_22),
.B1(n_24),
.B2(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_45),
.B1(n_64),
.B2(n_47),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_6),
.B(n_7),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_64),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_41),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_18),
.C(n_20),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_24),
.B1(n_35),
.B2(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_72),
.B1(n_79),
.B2(n_50),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_27),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_75),
.C(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_24),
.B1(n_35),
.B2(n_5),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_78),
.B1(n_53),
.B2(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_20),
.B1(n_9),
.B2(n_10),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_52),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_91),
.B(n_81),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_42),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_84),
.C(n_76),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_89),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_46),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_67),
.Y(n_96)
);

XNOR2x2_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_51),
.B1(n_76),
.B2(n_79),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.C(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_95),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_69),
.B(n_80),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_75),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_84),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_88),
.B1(n_97),
.B2(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_115),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_110),
.A3(n_108),
.B1(n_62),
.B2(n_66),
.C1(n_72),
.C2(n_54),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_118),
.A3(n_112),
.B1(n_54),
.B2(n_13),
.C1(n_8),
.C2(n_47),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_114),
.B1(n_115),
.B2(n_111),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_120),
.B(n_81),
.Y(n_121)
);


endmodule