module fake_netlist_6_4681_n_3120 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_3120);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_3120;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_835;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_462;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_595;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3037;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_432;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_1475;
wire n_884;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_600;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_444;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2502;
wire n_2131;
wire n_488;
wire n_2226;
wire n_2801;
wire n_497;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_1459;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_3109;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_906;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_501;
wire n_2276;
wire n_960;
wire n_956;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_3016;
wire n_1134;
wire n_3004;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_466;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_2050;
wire n_1472;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_2789;
wire n_3105;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_2670;
wire n_1332;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_2258;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_3075;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_799;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_706;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_911;
wire n_1737;
wire n_1464;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_3035;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1362;
wire n_1156;
wire n_2600;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_753;
wire n_1753;
wire n_3095;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_457;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_629;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_3054;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g420 ( 
.A(n_125),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_125),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_5),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_347),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_212),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_39),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_153),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_306),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_392),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_187),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_155),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_130),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_284),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_311),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_37),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_161),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_227),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_82),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_163),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_45),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_61),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_281),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_244),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_50),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_61),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_112),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_49),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_243),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_139),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_267),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_81),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_69),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_207),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_50),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_191),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_333),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_291),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_376),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_131),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_245),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_8),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_222),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_137),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_387),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_323),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_143),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_225),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_367),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_330),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_95),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_349),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_116),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_138),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_32),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_51),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_242),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_146),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_115),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_410),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_98),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_248),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_101),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_181),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_37),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_342),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_350),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_343),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_124),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_143),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_55),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_59),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_182),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_268),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_30),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_355),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_94),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_326),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_256),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_319),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_198),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_341),
.Y(n_503)
);

BUFx5_ASAP7_75t_L g504 ( 
.A(n_111),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_142),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_298),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_278),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_219),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_77),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_325),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_45),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_254),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_403),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_312),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_41),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_127),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_204),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_301),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_4),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_107),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_384),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_411),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_38),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_381),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_370),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_229),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_173),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_48),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_137),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_395),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_38),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_190),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_405),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_14),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_246),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_339),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_199),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_28),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_280),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_54),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_238),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_320),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_64),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_331),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_364),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_317),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_5),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_121),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_358),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_197),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_161),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_146),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_372),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_189),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_345),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_318),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_336),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_150),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_83),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_262),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_378),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_293),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_170),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_252),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_390),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_203),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_194),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_329),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_141),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_153),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_231),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_41),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_232),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_175),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_62),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_201),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_338),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_59),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_216),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_3),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_83),
.Y(n_582)
);

BUFx5_ASAP7_75t_L g583 ( 
.A(n_346),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_380),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_180),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_71),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_186),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_103),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_271),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_383),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_406),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_68),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_96),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_56),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_401),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_249),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_133),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_288),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_71),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_253),
.Y(n_600)
);

BUFx2_ASAP7_75t_SL g601 ( 
.A(n_260),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_78),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_213),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_53),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_186),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_223),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_133),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_351),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_101),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_130),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_53),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_261),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_10),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_374),
.Y(n_614)
);

CKINVDCx14_ASAP7_75t_R g615 ( 
.A(n_294),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_158),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_18),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_234),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_366),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_295),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_314),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_88),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_76),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_104),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_90),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_10),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_251),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_175),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_386),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_283),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_171),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_279),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_328),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_34),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_135),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_211),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_76),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_56),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_396),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_235),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_413),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_321),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_181),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_162),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_139),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_6),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_182),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_409),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_48),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_105),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_27),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_40),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_163),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_128),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_369),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_78),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_277),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_35),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_9),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_159),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_124),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_303),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_33),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_191),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_286),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_51),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_115),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_138),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_385),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_66),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_275),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_12),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_302),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_12),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_308),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_172),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_208),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_200),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_353),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_171),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_94),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_104),
.Y(n_682)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_118),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_230),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_75),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_379),
.Y(n_686)
);

CKINVDCx14_ASAP7_75t_R g687 ( 
.A(n_322),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_131),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_15),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_44),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_147),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_217),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_136),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_8),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_316),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_189),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_272),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_128),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_106),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_25),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_263),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_210),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_127),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_26),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_266),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_359),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_142),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_99),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_418),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_148),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_80),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_221),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_18),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_141),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_255),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_144),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_120),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_167),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_205),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_178),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_190),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_123),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_335),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_407),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_23),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_4),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_504),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_473),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_504),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_504),
.Y(n_730)
);

INVxp33_ASAP7_75t_L g731 ( 
.A(n_429),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_469),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_504),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_504),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_442),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_559),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_504),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_504),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_504),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_433),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_645),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_645),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_645),
.Y(n_743)
);

INVxp33_ASAP7_75t_SL g744 ( 
.A(n_699),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_497),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_645),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_574),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_645),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_645),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_645),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_645),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_611),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_585),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_512),
.Y(n_754)
);

INVxp33_ASAP7_75t_SL g755 ( 
.A(n_425),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_585),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_585),
.Y(n_757)
);

INVx4_ASAP7_75t_R g758 ( 
.A(n_641),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_564),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_585),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_585),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_695),
.B(n_0),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_680),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_680),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_680),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_439),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_680),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_644),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_641),
.Y(n_769)
);

CKINVDCx16_ASAP7_75t_R g770 ( 
.A(n_607),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_683),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_680),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_721),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_721),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_721),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_721),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_439),
.Y(n_777)
);

INVxp33_ASAP7_75t_L g778 ( 
.A(n_420),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_433),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_509),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_509),
.Y(n_781)
);

INVxp33_ASAP7_75t_SL g782 ( 
.A(n_425),
.Y(n_782)
);

INVxp33_ASAP7_75t_L g783 ( 
.A(n_437),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_631),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_631),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_660),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_660),
.Y(n_787)
);

INVxp33_ASAP7_75t_SL g788 ( 
.A(n_430),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_430),
.Y(n_789)
);

INVxp33_ASAP7_75t_SL g790 ( 
.A(n_431),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_721),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_583),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_671),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_688),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_688),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_583),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_718),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_505),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_505),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_718),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_479),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_446),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_449),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_454),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_461),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_444),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_476),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_671),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_480),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_484),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_491),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_431),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_615),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_583),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_540),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_493),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_517),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_496),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_511),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_515),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_547),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_529),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_530),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_544),
.Y(n_824)
);

CKINVDCx14_ASAP7_75t_R g825 ( 
.A(n_687),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_434),
.Y(n_826)
);

INVxp33_ASAP7_75t_SL g827 ( 
.A(n_434),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_583),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_568),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_570),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_505),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_573),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_582),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_588),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_592),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_583),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_427),
.B(n_0),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_563),
.Y(n_838)
);

INVxp33_ASAP7_75t_SL g839 ( 
.A(n_438),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_597),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_450),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_605),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_427),
.B(n_1),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_457),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_609),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_610),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_616),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_458),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_444),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_460),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_494),
.Y(n_851)
);

INVxp33_ASAP7_75t_SL g852 ( 
.A(n_438),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_494),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_482),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_433),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_628),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_547),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_638),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_647),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_649),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_651),
.Y(n_861)
);

XOR2xp5_ASAP7_75t_L g862 ( 
.A(n_426),
.B(n_1),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_485),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_652),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_583),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_486),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_735),
.B(n_572),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_740),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_808),
.B(n_572),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_791),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_791),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_740),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_744),
.A2(n_535),
.B1(n_477),
.B2(n_445),
.Y(n_873)
);

BUFx12f_ASAP7_75t_L g874 ( 
.A(n_728),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_776),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_769),
.B(n_549),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_744),
.A2(n_762),
.B1(n_782),
.B2(n_755),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_740),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_821),
.Y(n_880)
);

BUFx8_ASAP7_75t_SL g881 ( 
.A(n_752),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_769),
.Y(n_882)
);

AND2x6_ASAP7_75t_L g883 ( 
.A(n_740),
.B(n_433),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_776),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_776),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_793),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_753),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_753),
.Y(n_888)
);

OAI22x1_ASAP7_75t_R g889 ( 
.A1(n_831),
.A2(n_519),
.B1(n_520),
.B2(n_516),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_755),
.A2(n_603),
.B1(n_636),
.B2(n_565),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_756),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_779),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_779),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_732),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_779),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_727),
.A2(n_470),
.B(n_443),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_756),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_757),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_747),
.B(n_614),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_771),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_779),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_757),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_793),
.B(n_549),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_779),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_760),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_855),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_855),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_760),
.Y(n_908)
);

BUFx12f_ASAP7_75t_L g909 ( 
.A(n_728),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_855),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_855),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_841),
.B(n_614),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_761),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_844),
.B(n_848),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_782),
.A2(n_669),
.B1(n_722),
.B2(n_672),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_745),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_761),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_855),
.Y(n_918)
);

AOI22x1_ASAP7_75t_SL g919 ( 
.A1(n_754),
.A2(n_541),
.B1(n_587),
.B2(n_523),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_763),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_763),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_764),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_764),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_765),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_788),
.A2(n_790),
.B1(n_839),
.B2(n_827),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_759),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_850),
.B(n_443),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_825),
.B(n_815),
.Y(n_928)
);

AOI22x1_ASAP7_75t_SL g929 ( 
.A1(n_817),
.A2(n_623),
.B1(n_661),
.B2(n_622),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_813),
.B(n_766),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_765),
.B(n_470),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_749),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_759),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_771),
.Y(n_934)
);

AND2x2_ASAP7_75t_SL g935 ( 
.A(n_837),
.B(n_508),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_767),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_766),
.B(n_508),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_767),
.B(n_569),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_772),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_772),
.Y(n_940)
);

OA21x2_ASAP7_75t_L g941 ( 
.A1(n_733),
.A2(n_584),
.B(n_569),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_773),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_734),
.A2(n_702),
.B(n_584),
.Y(n_943)
);

OA22x2_ASAP7_75t_SL g944 ( 
.A1(n_862),
.A2(n_663),
.B1(n_664),
.B2(n_659),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_821),
.B(n_702),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_737),
.A2(n_474),
.B(n_464),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_773),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_774),
.B(n_487),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_774),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_775),
.B(n_501),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_775),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_777),
.B(n_617),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_729),
.B(n_526),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_780),
.B(n_781),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_738),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_729),
.B(n_433),
.Y(n_956)
);

AOI22x1_ASAP7_75t_SL g957 ( 
.A1(n_838),
.A2(n_725),
.B1(n_691),
.B2(n_445),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_801),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_784),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_792),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_785),
.B(n_617),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_736),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_796),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_788),
.A2(n_492),
.B1(n_498),
.B2(n_490),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_730),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_730),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_739),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_801),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_739),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_802),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_854),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_814),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_741),
.Y(n_973)
);

BUFx8_ASAP7_75t_L g974 ( 
.A(n_752),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_741),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_SL g976 ( 
.A1(n_862),
.A2(n_447),
.B1(n_451),
.B2(n_440),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_854),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_742),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_742),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_743),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_743),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_828),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_790),
.A2(n_532),
.B1(n_533),
.B2(n_528),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_746),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_746),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_748),
.A2(n_536),
.B(n_527),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_748),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_977),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_977),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_969),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_880),
.B(n_863),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_914),
.B(n_935),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_969),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_894),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_882),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_881),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_894),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_916),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_975),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_867),
.B(n_843),
.C(n_863),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_882),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_986),
.A2(n_751),
.B(n_750),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_916),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_975),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_868),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_986),
.A2(n_946),
.B(n_941),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_874),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_914),
.B(n_750),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_970),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_980),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_880),
.B(n_866),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_874),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_909),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_909),
.Y(n_1014)
);

AND2x6_ASAP7_75t_L g1015 ( 
.A(n_953),
.B(n_525),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_881),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_886),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_914),
.B(n_751),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_R g1019 ( 
.A(n_958),
.B(n_866),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_926),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_980),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_870),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_980),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_870),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_974),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_871),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_871),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_868),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_926),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_935),
.B(n_857),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_981),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_868),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_933),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_886),
.Y(n_1034)
);

OA21x2_ASAP7_75t_L g1035 ( 
.A1(n_946),
.A2(n_836),
.B(n_828),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_981),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_887),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_933),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_868),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_981),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_868),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_958),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_968),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_971),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_900),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_876),
.B(n_440),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_974),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_953),
.B(n_803),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_R g1049 ( 
.A(n_930),
.B(n_770),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_954),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_900),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_954),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_962),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_974),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_890),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_876),
.B(n_857),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_872),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_959),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_SL g1059 ( 
.A(n_903),
.B(n_447),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_919),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_959),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_967),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_953),
.B(n_804),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_967),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_919),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_872),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_979),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_979),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_984),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_929),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_887),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_948),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_879),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_984),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_879),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_SL g1076 ( 
.A(n_934),
.B(n_558),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_928),
.B(n_481),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_903),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_888),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_925),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_929),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_948),
.B(n_805),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_957),
.Y(n_1083)
);

AND2x6_ASAP7_75t_L g1084 ( 
.A(n_912),
.B(n_525),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_985),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_888),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_948),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_957),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_950),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_985),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_878),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_987),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_899),
.B(n_789),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_889),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_912),
.B(n_506),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_987),
.Y(n_1096)
);

XNOR2xp5_ASAP7_75t_L g1097 ( 
.A(n_915),
.B(n_827),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_945),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_976),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_955),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_869),
.B(n_839),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_897),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_897),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_952),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_955),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_964),
.Y(n_1106)
);

BUFx8_ASAP7_75t_L g1107 ( 
.A(n_952),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_983),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_955),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_891),
.A2(n_865),
.B(n_836),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_898),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_955),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_879),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_879),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_912),
.B(n_812),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_898),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_955),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_965),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_927),
.B(n_590),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

NAND2x1_ASAP7_75t_L g1121 ( 
.A(n_883),
.B(n_758),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_965),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_873),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_902),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_965),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_927),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_965),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_927),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_966),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_902),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_936),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_961),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_892),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_892),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_966),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_966),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_966),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_961),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_901),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_950),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_937),
.B(n_483),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_950),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_966),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_931),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_973),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_973),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_931),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_973),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_973),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_931),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_938),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1053),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1098),
.B(n_932),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_992),
.B(n_1126),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1006),
.A2(n_550),
.B(n_543),
.Y(n_1155)
);

NAND2xp33_ASAP7_75t_L g1156 ( 
.A(n_1084),
.B(n_583),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1144),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1056),
.B(n_826),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1045),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1110),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1008),
.B(n_1018),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1110),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1072),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1009),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1128),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1110),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_990),
.B(n_932),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1022),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_995),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1072),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_1051),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1022),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_993),
.B(n_932),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1024),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1087),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1087),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1030),
.B(n_768),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1101),
.B(n_852),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1089),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1126),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1089),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1050),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1052),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1058),
.Y(n_1184)
);

BUFx4f_ASAP7_75t_L g1185 ( 
.A(n_991),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1024),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1138),
.B(n_973),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1095),
.A2(n_731),
.B1(n_852),
.B2(n_422),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1026),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1061),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1091),
.A2(n_709),
.B1(n_547),
.B2(n_601),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_999),
.B(n_960),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1004),
.B(n_960),
.Y(n_1193)
);

OR2x6_ASAP7_75t_L g1194 ( 
.A(n_996),
.B(n_798),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1048),
.Y(n_1195)
);

AND3x1_ASAP7_75t_L g1196 ( 
.A(n_1076),
.B(n_944),
.C(n_787),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1048),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_SL g1198 ( 
.A(n_1138),
.B(n_1115),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1093),
.B(n_960),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1026),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1011),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1048),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1078),
.B(n_963),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1000),
.B(n_963),
.Y(n_1204)
);

XNOR2xp5_ASAP7_75t_L g1205 ( 
.A(n_994),
.B(n_423),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1027),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1063),
.Y(n_1207)
);

BUFx4f_ASAP7_75t_L g1208 ( 
.A(n_1063),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1027),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1037),
.Y(n_1210)
);

AND2x6_ASAP7_75t_L g1211 ( 
.A(n_1010),
.B(n_525),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1063),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1119),
.B(n_963),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1082),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_995),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1082),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_994),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1082),
.Y(n_1218)
);

AND2x6_ASAP7_75t_L g1219 ( 
.A(n_1021),
.B(n_525),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1046),
.B(n_799),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1037),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1023),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1031),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1140),
.B(n_978),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1071),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1036),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1040),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1071),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1147),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1104),
.B(n_778),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1140),
.A2(n_1142),
.B1(n_1150),
.B2(n_1147),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1132),
.B(n_972),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1084),
.B(n_972),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1079),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1150),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1142),
.B(n_1151),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1006),
.A2(n_556),
.B(n_554),
.Y(n_1237)
);

NAND2xp33_ASAP7_75t_SL g1238 ( 
.A(n_1106),
.B(n_525),
.Y(n_1238)
);

BUFx8_ASAP7_75t_SL g1239 ( 
.A(n_1016),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1084),
.B(n_972),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1084),
.B(n_982),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1151),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1062),
.B(n_1064),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1079),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1086),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1086),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1084),
.B(n_982),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1102),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1042),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1102),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1067),
.B(n_978),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1001),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1068),
.B(n_978),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_997),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1084),
.A2(n_941),
.B1(n_943),
.B2(n_896),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1103),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_998),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1017),
.B(n_786),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1015),
.A2(n_941),
.B1(n_943),
.B2(n_896),
.Y(n_1259)
);

INVxp33_ASAP7_75t_L g1260 ( 
.A(n_1049),
.Y(n_1260)
);

AO22x2_ASAP7_75t_L g1261 ( 
.A1(n_1091),
.A2(n_435),
.B1(n_471),
.B2(n_421),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1069),
.B(n_982),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1074),
.B(n_1085),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1015),
.A2(n_943),
.B1(n_896),
.B2(n_666),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1034),
.B(n_783),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1103),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1107),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1111),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1111),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1116),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1090),
.B(n_978),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1116),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1124),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1028),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1092),
.B(n_561),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1123),
.A2(n_674),
.B1(n_685),
.B2(n_668),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1124),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1043),
.B(n_829),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1130),
.Y(n_1279)
);

AND2x6_ASAP7_75t_L g1280 ( 
.A(n_1118),
.B(n_1143),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1096),
.B(n_978),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1130),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1120),
.B(n_938),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1044),
.B(n_794),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1122),
.B(n_938),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1131),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1131),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1002),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1002),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1100),
.B(n_567),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1107),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1035),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1035),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1035),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1005),
.Y(n_1295)
);

AND2x6_ASAP7_75t_L g1296 ( 
.A(n_1125),
.B(n_606),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1127),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1028),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1107),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1015),
.A2(n_698),
.B1(n_707),
.B2(n_703),
.Y(n_1300)
);

INVxp33_ASAP7_75t_L g1301 ( 
.A(n_1097),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1015),
.A2(n_720),
.B1(n_710),
.B2(n_700),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1005),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1077),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1003),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1005),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1007),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1121),
.B(n_795),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1129),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1015),
.A2(n_553),
.B1(n_642),
.B2(n_606),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1028),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1039),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1106),
.A2(n_489),
.B1(n_495),
.B2(n_488),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1028),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1039),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1135),
.B(n_905),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1136),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1054),
.B(n_797),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1032),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1137),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1145),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1039),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1032),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1146),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1046),
.B(n_800),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1057),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1148),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1057),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1057),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1105),
.B(n_580),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1066),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1032),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1108),
.B(n_423),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1149),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1059),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1109),
.B(n_606),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1112),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1117),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1108),
.B(n_424),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1012),
.B(n_846),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1032),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1059),
.B(n_807),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1015),
.A2(n_606),
.B1(n_719),
.B2(n_642),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1055),
.B(n_809),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1066),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1066),
.B(n_591),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1073),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1250),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1168),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1168),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1163),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1268),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1270),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1172),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1169),
.B(n_810),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1230),
.B(n_1080),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1152),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1163),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1169),
.B(n_632),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1199),
.B(n_1141),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1215),
.B(n_633),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1199),
.B(n_1139),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1265),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1278),
.B(n_1123),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1277),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1163),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1215),
.B(n_639),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1217),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1172),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1258),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1174),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1158),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1185),
.B(n_1041),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1163),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1252),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1170),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1161),
.B(n_1232),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1174),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1232),
.B(n_1139),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1344),
.B(n_988),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1186),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1195),
.B(n_811),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1287),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1153),
.B(n_1073),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1197),
.B(n_640),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1202),
.B(n_816),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1239),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1186),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1207),
.B(n_818),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1263),
.Y(n_1390)
);

NAND2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1208),
.B(n_1073),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1210),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1291),
.B(n_1012),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1210),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1178),
.A2(n_1099),
.B1(n_1094),
.B2(n_1060),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1239),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1189),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1221),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1221),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1178),
.B(n_1139),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1213),
.B(n_1075),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1225),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1189),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1254),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1200),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1225),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1234),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_1333),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1170),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1212),
.B(n_819),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1200),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1170),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1165),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1154),
.B(n_988),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1170),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1234),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1295),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1284),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1203),
.B(n_1204),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1177),
.B(n_989),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1311),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1214),
.B(n_820),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1209),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1311),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1244),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1217),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1238),
.A2(n_1204),
.B(n_1182),
.C(n_1183),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1209),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1244),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1246),
.Y(n_1430)
);

BUFx4f_ASAP7_75t_L g1431 ( 
.A(n_1235),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1246),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1248),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1216),
.B(n_665),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1248),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1218),
.B(n_822),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1256),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1159),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1256),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1201),
.B(n_989),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1154),
.B(n_1335),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1276),
.A2(n_1019),
.B1(n_1099),
.B2(n_452),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1266),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1311),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1266),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1269),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1185),
.B(n_1041),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1171),
.B(n_1033),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1269),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1272),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1272),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1311),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1273),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1175),
.B(n_1176),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1333),
.B(n_1013),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1273),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1279),
.Y(n_1457)
);

INVx8_ASAP7_75t_L g1458 ( 
.A(n_1258),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1314),
.Y(n_1459)
);

NOR2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1267),
.B(n_1013),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1314),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1295),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1276),
.A2(n_452),
.B1(n_455),
.B2(n_451),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1279),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1314),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1208),
.B(n_1041),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1249),
.B(n_1038),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1295),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1282),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1310),
.A2(n_583),
.B1(n_642),
.B2(n_606),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1198),
.A2(n_1113),
.B1(n_1114),
.B2(n_1075),
.Y(n_1471)
);

AND2x6_ASAP7_75t_L g1472 ( 
.A(n_1160),
.B(n_642),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1282),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1286),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1314),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1179),
.B(n_673),
.Y(n_1476)
);

AO22x2_ASAP7_75t_L g1477 ( 
.A1(n_1342),
.A2(n_686),
.B1(n_712),
.B2(n_675),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1286),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1164),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1292),
.B(n_1075),
.Y(n_1480)
);

BUFx4f_ASAP7_75t_L g1481 ( 
.A(n_1242),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1258),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1222),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1223),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1319),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1160),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1226),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1227),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1252),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1180),
.B(n_1014),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1319),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1292),
.B(n_1113),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1180),
.B(n_1014),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1187),
.B(n_1113),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1228),
.Y(n_1495)
);

NOR2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1267),
.B(n_1020),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1303),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1319),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1229),
.B(n_1020),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1358),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1377),
.B(n_1187),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1357),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1390),
.B(n_1304),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1419),
.B(n_1181),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1470),
.A2(n_1302),
.B1(n_1310),
.B2(n_1261),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1441),
.B(n_1339),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1441),
.B(n_1229),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1360),
.B(n_1198),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1486),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1427),
.B(n_1264),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1372),
.B(n_1418),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1427),
.A2(n_1220),
.B(n_1325),
.C(n_1236),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1400),
.B(n_1339),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_SL g1514 ( 
.A(n_1455),
.B(n_1254),
.C(n_1191),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1408),
.B(n_1358),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1408),
.B(n_1264),
.Y(n_1516)
);

OR2x2_ASAP7_75t_SL g1517 ( 
.A(n_1448),
.B(n_1094),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1470),
.A2(n_1302),
.B1(n_1261),
.B2(n_1238),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1479),
.B(n_1224),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1372),
.B(n_1418),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1358),
.B(n_1224),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1363),
.A2(n_1260),
.B1(n_1257),
.B2(n_1313),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1375),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1358),
.B(n_1231),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1483),
.B(n_1184),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1409),
.B(n_1196),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1368),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1356),
.B(n_1157),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1409),
.Y(n_1529)
);

NAND3xp33_ASAP7_75t_SL g1530 ( 
.A(n_1455),
.B(n_1029),
.C(n_1260),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1392),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1364),
.A2(n_1236),
.B1(n_1190),
.B2(n_1305),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1404),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1484),
.B(n_1188),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1487),
.B(n_1275),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1488),
.B(n_1363),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1362),
.B(n_1275),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1477),
.A2(n_1261),
.B1(n_1300),
.B2(n_1343),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1348),
.B(n_1275),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1394),
.Y(n_1540)
);

NOR3xp33_ASAP7_75t_L g1541 ( 
.A(n_1380),
.B(n_1029),
.C(n_1070),
.Y(n_1541)
);

NOR2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1387),
.B(n_1299),
.Y(n_1542)
);

NOR2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1387),
.B(n_1299),
.Y(n_1543)
);

AND2x6_ASAP7_75t_SL g1544 ( 
.A(n_1393),
.B(n_1194),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1352),
.B(n_1167),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1413),
.B(n_1301),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1490),
.B(n_1205),
.Y(n_1547)
);

INVx6_ASAP7_75t_L g1548 ( 
.A(n_1375),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1398),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1414),
.A2(n_1243),
.B1(n_1330),
.B2(n_1290),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1399),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1420),
.B(n_1438),
.Y(n_1552)
);

AND2x6_ASAP7_75t_L g1553 ( 
.A(n_1486),
.B(n_1293),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1353),
.B(n_1365),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1413),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1349),
.Y(n_1556)
);

BUFx4f_ASAP7_75t_L g1557 ( 
.A(n_1458),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1414),
.A2(n_1243),
.B1(n_1330),
.B2(n_1290),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1442),
.B(n_1301),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_L g1560 ( 
.A(n_1409),
.B(n_1280),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1402),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1383),
.B(n_1173),
.Y(n_1562)
);

NOR2x1p5_ASAP7_75t_L g1563 ( 
.A(n_1396),
.B(n_1307),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1480),
.A2(n_1298),
.B(n_1274),
.Y(n_1564)
);

AND2x6_ASAP7_75t_SL g1565 ( 
.A(n_1393),
.B(n_1194),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1406),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1379),
.B(n_1192),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1421),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1385),
.B(n_1193),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1395),
.A2(n_1025),
.B1(n_1047),
.B2(n_1060),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1385),
.B(n_1228),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1385),
.B(n_1228),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1489),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1489),
.B(n_1307),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1494),
.A2(n_1401),
.B(n_1492),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1493),
.B(n_1340),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1355),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1409),
.B(n_1255),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1454),
.B(n_1308),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1407),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1434),
.B(n_1245),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1416),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1404),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1477),
.A2(n_1300),
.B1(n_1343),
.B2(n_1330),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1417),
.B(n_1255),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1434),
.B(n_1245),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1425),
.Y(n_1587)
);

AO22x1_ASAP7_75t_L g1588 ( 
.A1(n_1506),
.A2(n_1499),
.B1(n_1070),
.B2(n_1440),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1559),
.A2(n_1355),
.B1(n_1361),
.B2(n_1359),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1553),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1502),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1533),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_R g1593 ( 
.A(n_1530),
.B(n_1426),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1555),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1509),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1568),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1509),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1568),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1548),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1568),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1512),
.B(n_1391),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1568),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1548),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1513),
.A2(n_1481),
.B1(n_1431),
.B2(n_1467),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1503),
.B(n_1546),
.Y(n_1606)
);

AO22x1_ASAP7_75t_L g1607 ( 
.A1(n_1559),
.A2(n_1088),
.B1(n_1083),
.B2(n_1359),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1548),
.Y(n_1608)
);

BUFx4f_ASAP7_75t_L g1609 ( 
.A(n_1579),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1553),
.Y(n_1610)
);

INVx5_ASAP7_75t_L g1611 ( 
.A(n_1553),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1554),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1546),
.B(n_1507),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1556),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1519),
.B(n_1477),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1552),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1511),
.B(n_1442),
.Y(n_1618)
);

BUFx8_ASAP7_75t_L g1619 ( 
.A(n_1527),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1583),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_SL g1621 ( 
.A(n_1514),
.B(n_1088),
.C(n_1083),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1528),
.B(n_1349),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1583),
.B(n_1426),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1556),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1511),
.B(n_1382),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_SL g1626 ( 
.A(n_1522),
.B(n_1463),
.C(n_1396),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1520),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1553),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_SL g1629 ( 
.A(n_1532),
.B(n_1047),
.C(n_1025),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1577),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1553),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1574),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1508),
.A2(n_1481),
.B(n_1431),
.C(n_1434),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1531),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1507),
.B(n_1536),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1574),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1557),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1540),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1547),
.B(n_1370),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1534),
.B(n_1382),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1595),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1631),
.A2(n_1575),
.B(n_1564),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1631),
.A2(n_1510),
.B(n_1521),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1590),
.A2(n_1510),
.B(n_1521),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1606),
.A2(n_1505),
.B1(n_1518),
.B2(n_1584),
.Y(n_1645)
);

AOI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1601),
.A2(n_1508),
.B(n_1567),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1637),
.B(n_1524),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1626),
.A2(n_1505),
.B(n_1518),
.C(n_1584),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1590),
.A2(n_1578),
.B(n_1515),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1590),
.A2(n_1578),
.B(n_1515),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1612),
.A2(n_1537),
.B(n_1585),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1368),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1601),
.A2(n_1585),
.B(n_1560),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1610),
.A2(n_1391),
.B(n_1289),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1640),
.A2(n_1569),
.B(n_1558),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1637),
.B(n_1524),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1601),
.A2(n_1516),
.B(n_1545),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1613),
.B(n_1576),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1601),
.A2(n_1516),
.B(n_1562),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1589),
.A2(n_1618),
.B1(n_1625),
.B2(n_1605),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1627),
.B(n_1463),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1611),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1633),
.B(n_1550),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1616),
.B(n_1549),
.Y(n_1664)
);

AOI21x1_ASAP7_75t_SL g1665 ( 
.A1(n_1616),
.A2(n_1635),
.B(n_1361),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1594),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1610),
.A2(n_1628),
.B(n_1615),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1617),
.B(n_1016),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1611),
.A2(n_1466),
.B(n_1447),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1610),
.A2(n_1289),
.B(n_1288),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1592),
.Y(n_1672)
);

INVx5_ASAP7_75t_L g1673 ( 
.A(n_1611),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1628),
.A2(n_1288),
.B(n_1466),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1603),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1622),
.B(n_1525),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1609),
.A2(n_1517),
.B1(n_1538),
.B2(n_1557),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1622),
.B(n_1535),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1611),
.A2(n_1447),
.B(n_1373),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1611),
.A2(n_1366),
.B(n_1351),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1593),
.B(n_1541),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1615),
.Y(n_1682)
);

AOI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1634),
.A2(n_1373),
.B(n_1526),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1638),
.A2(n_1384),
.B(n_1316),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1632),
.B(n_1579),
.Y(n_1685)
);

AOI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1638),
.A2(n_1526),
.B(n_1253),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1609),
.B(n_1539),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1595),
.B(n_1597),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1632),
.B(n_1386),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1597),
.A2(n_1281),
.B(n_1271),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1669),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1676),
.B(n_1591),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1672),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1675),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1641),
.Y(n_1695)
);

AND2x2_ASAP7_75t_SL g1696 ( 
.A(n_1647),
.B(n_1538),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1647),
.B(n_1636),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1641),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1664),
.B(n_1596),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1647),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1656),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1663),
.A2(n_1609),
.B(n_1572),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1666),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1666),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1655),
.B(n_1621),
.Y(n_1705)
);

BUFx12f_ASAP7_75t_L g1706 ( 
.A(n_1672),
.Y(n_1706)
);

BUFx12f_ASAP7_75t_L g1707 ( 
.A(n_1675),
.Y(n_1707)
);

CKINVDCx8_ASAP7_75t_R g1708 ( 
.A(n_1668),
.Y(n_1708)
);

INVxp67_ASAP7_75t_SL g1709 ( 
.A(n_1684),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1652),
.B(n_1592),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1657),
.A2(n_1581),
.B(n_1571),
.Y(n_1711)
);

INVx3_ASAP7_75t_SL g1712 ( 
.A(n_1681),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1664),
.B(n_1636),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1656),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1685),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1656),
.B(n_1608),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1678),
.B(n_1588),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1688),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1658),
.Y(n_1719)
);

OR2x6_ASAP7_75t_L g1720 ( 
.A(n_1653),
.B(n_1588),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1688),
.B(n_1596),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1677),
.Y(n_1722)
);

INVx2_ASAP7_75t_R g1723 ( 
.A(n_1673),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1662),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1682),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1661),
.Y(n_1727)
);

AND2x4_ASAP7_75t_SL g1728 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1643),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1673),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1673),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1643),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1660),
.B(n_1630),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1673),
.B(n_1608),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1689),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_SL g1737 ( 
.A1(n_1645),
.A2(n_1065),
.B1(n_1081),
.B2(n_1629),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1683),
.Y(n_1738)
);

O2A1O1Ixp5_ASAP7_75t_L g1739 ( 
.A1(n_1646),
.A2(n_1607),
.B(n_1639),
.C(n_1366),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1659),
.B(n_1623),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1680),
.A2(n_1586),
.B(n_1237),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1648),
.B(n_1607),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1673),
.B(n_1596),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1687),
.B(n_1624),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1651),
.B(n_1624),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1667),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1649),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1649),
.B(n_1599),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1644),
.B(n_1359),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1651),
.A2(n_1081),
.B1(n_1065),
.B2(n_1570),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1667),
.Y(n_1751)
);

INVx5_ASAP7_75t_L g1752 ( 
.A(n_1665),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1683),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1670),
.B(n_459),
.C(n_455),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1686),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_SL g1756 ( 
.A(n_1679),
.B(n_1620),
.C(n_463),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1686),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1684),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1651),
.A2(n_1563),
.B1(n_1620),
.B2(n_1318),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1651),
.A2(n_463),
.B1(n_467),
.B2(n_459),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_SL g1761 ( 
.A(n_1680),
.B(n_1351),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1650),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1650),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1644),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1684),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1684),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1654),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1654),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_SL g1769 ( 
.A1(n_1646),
.A2(n_1376),
.B(n_1374),
.C(n_1529),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1674),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1674),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1642),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1671),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1671),
.Y(n_1774)
);

OR2x6_ASAP7_75t_SL g1775 ( 
.A(n_1642),
.B(n_467),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1690),
.A2(n_1156),
.B(n_1476),
.C(n_723),
.Y(n_1776)
);

OAI211xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1737),
.A2(n_824),
.B(n_830),
.C(n_823),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1705),
.B(n_1740),
.C(n_1754),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1741),
.A2(n_1690),
.B(n_1471),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1705),
.A2(n_1482),
.B(n_858),
.C(n_859),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1694),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1711),
.A2(n_1561),
.B(n_1551),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1742),
.B(n_1544),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1713),
.B(n_1599),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1715),
.B(n_1476),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1693),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1750),
.A2(n_1393),
.B1(n_1318),
.B2(n_1340),
.Y(n_1787)
);

NAND2x1p5_ASAP7_75t_L g1788 ( 
.A(n_1731),
.B(n_1752),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1707),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1772),
.A2(n_1580),
.B(n_1566),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1722),
.A2(n_1156),
.B(n_678),
.C(n_448),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1692),
.B(n_1476),
.Y(n_1792)
);

CKINVDCx16_ASAP7_75t_R g1793 ( 
.A(n_1693),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1764),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1698),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1691),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1707),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1772),
.A2(n_1587),
.B(n_1582),
.Y(n_1798)
);

INVx4_ASAP7_75t_L g1799 ( 
.A(n_1735),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1722),
.A2(n_571),
.B1(n_575),
.B2(n_475),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1700),
.B(n_1604),
.Y(n_1801)
);

OAI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1755),
.A2(n_1376),
.B(n_1374),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1755),
.A2(n_1529),
.B(n_1285),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_SL g1804 ( 
.A1(n_1740),
.A2(n_1604),
.B(n_1523),
.C(n_1565),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1700),
.B(n_1155),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1756),
.A2(n_1367),
.B(n_1361),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1699),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1695),
.Y(n_1808)
);

AOI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1761),
.A2(n_1336),
.B(n_1290),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1698),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1706),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1726),
.Y(n_1812)
);

OA21x2_ASAP7_75t_L g1813 ( 
.A1(n_1709),
.A2(n_849),
.B(n_806),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1757),
.A2(n_1283),
.B(n_1497),
.Y(n_1814)
);

OAI21x1_ASAP7_75t_L g1815 ( 
.A1(n_1757),
.A2(n_1497),
.B(n_1338),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1696),
.A2(n_571),
.B1(n_676),
.B2(n_575),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1718),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1763),
.A2(n_1337),
.B(n_1429),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1724),
.Y(n_1819)
);

OAI21x1_ASAP7_75t_L g1820 ( 
.A1(n_1763),
.A2(n_1478),
.B(n_1474),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1701),
.B(n_1714),
.Y(n_1821)
);

OAI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1738),
.A2(n_1432),
.B(n_1430),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1701),
.B(n_1542),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1726),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1714),
.B(n_1598),
.Y(n_1825)
);

AO21x2_ASAP7_75t_L g1826 ( 
.A1(n_1769),
.A2(n_1155),
.B(n_1336),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1730),
.Y(n_1827)
);

AO21x2_ASAP7_75t_L g1828 ( 
.A1(n_1769),
.A2(n_1367),
.B(n_1435),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1719),
.A2(n_1318),
.B1(n_1340),
.B2(n_1194),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1735),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1706),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1729),
.Y(n_1832)
);

INVxp67_ASAP7_75t_SL g1833 ( 
.A(n_1745),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1760),
.B(n_833),
.C(n_832),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1717),
.B(n_1367),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1719),
.B(n_539),
.Y(n_1836)
);

OA21x2_ASAP7_75t_L g1837 ( 
.A1(n_1709),
.A2(n_1758),
.B(n_1765),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_L g1838 ( 
.A1(n_1753),
.A2(n_1443),
.B(n_1437),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1697),
.B(n_1598),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1712),
.A2(n_1543),
.B1(n_1458),
.B2(n_1619),
.Y(n_1840)
);

OAI21x1_ASAP7_75t_L g1841 ( 
.A1(n_1774),
.A2(n_1450),
.B(n_1446),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1774),
.A2(n_1457),
.B(n_1453),
.Y(n_1842)
);

A2O1A1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1760),
.A2(n_428),
.B(n_432),
.C(n_424),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1748),
.Y(n_1844)
);

BUFx12f_ASAP7_75t_L g1845 ( 
.A(n_1736),
.Y(n_1845)
);

AOI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1749),
.A2(n_835),
.B(n_834),
.Y(n_1846)
);

NAND2x1p5_ASAP7_75t_L g1847 ( 
.A(n_1731),
.B(n_1598),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1748),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1767),
.A2(n_1464),
.B(n_1309),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_R g1850 ( 
.A(n_1727),
.B(n_1619),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1696),
.A2(n_432),
.B(n_436),
.C(n_428),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1712),
.B(n_856),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1703),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1704),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1758),
.A2(n_849),
.B(n_806),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1734),
.B(n_851),
.Y(n_1856)
);

BUFx4f_ASAP7_75t_SL g1857 ( 
.A(n_1716),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1767),
.A2(n_1317),
.B(n_1297),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1733),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1727),
.B(n_851),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1736),
.B(n_548),
.Y(n_1861)
);

OA21x2_ASAP7_75t_L g1862 ( 
.A1(n_1766),
.A2(n_853),
.B(n_856),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1720),
.B(n_853),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1768),
.A2(n_1321),
.B(n_1320),
.Y(n_1864)
);

AO21x2_ASAP7_75t_L g1865 ( 
.A1(n_1759),
.A2(n_1346),
.B(n_1327),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1702),
.A2(n_681),
.B1(n_682),
.B2(n_676),
.C(n_475),
.Y(n_1866)
);

AOI21x1_ASAP7_75t_L g1867 ( 
.A1(n_1720),
.A2(n_842),
.B(n_840),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1768),
.A2(n_1334),
.B(n_1324),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1766),
.A2(n_1739),
.B(n_1746),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1776),
.A2(n_1240),
.B(n_1233),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1746),
.A2(n_1354),
.B(n_1350),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1751),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1751),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1762),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1720),
.A2(n_682),
.B1(n_689),
.B2(n_681),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1776),
.A2(n_1389),
.B(n_1386),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1697),
.B(n_552),
.Y(n_1877)
);

AO21x2_ASAP7_75t_L g1878 ( 
.A1(n_1744),
.A2(n_1346),
.B(n_1253),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1762),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1762),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1699),
.B(n_1598),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1710),
.A2(n_1708),
.B1(n_1752),
.B2(n_1775),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1747),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1752),
.A2(n_1496),
.B1(n_1460),
.B2(n_1458),
.Y(n_1884)
);

OA21x2_ASAP7_75t_L g1885 ( 
.A1(n_1771),
.A2(n_859),
.B(n_858),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1725),
.A2(n_1354),
.B(n_1350),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1752),
.A2(n_1410),
.B(n_1389),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1747),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1699),
.B(n_555),
.Y(n_1889)
);

BUFx8_ASAP7_75t_L g1890 ( 
.A(n_1716),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1721),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1721),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1732),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1721),
.B(n_1598),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1725),
.A2(n_1422),
.B(n_1410),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1771),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1732),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1723),
.A2(n_1371),
.B(n_1369),
.Y(n_1898)
);

O2A1O1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1773),
.A2(n_861),
.B(n_864),
.C(n_860),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1762),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_SL g1901 ( 
.A(n_1743),
.B(n_1619),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1732),
.B(n_1600),
.Y(n_1902)
);

OA21x2_ASAP7_75t_L g1903 ( 
.A1(n_1743),
.A2(n_861),
.B(n_860),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1728),
.Y(n_1904)
);

OA21x2_ASAP7_75t_L g1905 ( 
.A1(n_1743),
.A2(n_864),
.B(n_847),
.Y(n_1905)
);

OA21x2_ASAP7_75t_L g1906 ( 
.A1(n_1723),
.A2(n_845),
.B(n_1251),
.Y(n_1906)
);

OAI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1731),
.A2(n_1436),
.B(n_1422),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1731),
.A2(n_1371),
.B(n_1369),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_SL g1909 ( 
.A(n_1730),
.B(n_1600),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1770),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1770),
.Y(n_1911)
);

OAI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1730),
.A2(n_1381),
.B(n_1378),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1730),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1728),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1715),
.B(n_560),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1707),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1741),
.A2(n_1381),
.B(n_1378),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1691),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1705),
.B(n_689),
.Y(n_1919)
);

CKINVDCx6p67_ASAP7_75t_R g1920 ( 
.A(n_1693),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1698),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1700),
.B(n_1600),
.Y(n_1922)
);

BUFx3_ASAP7_75t_L g1923 ( 
.A(n_1707),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1700),
.B(n_1436),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1691),
.Y(n_1925)
);

OAI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1705),
.A2(n_1454),
.B(n_1346),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1705),
.A2(n_1495),
.B(n_1251),
.C(n_1397),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1700),
.B(n_1600),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1807),
.B(n_1600),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1923),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1796),
.Y(n_1931)
);

NAND2x1_ASAP7_75t_L g1932 ( 
.A(n_1885),
.B(n_1602),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1918),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1778),
.A2(n_1415),
.B(n_1412),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1891),
.B(n_1602),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1919),
.A2(n_709),
.B1(n_719),
.B2(n_642),
.Y(n_1936)
);

BUFx10_ASAP7_75t_L g1937 ( 
.A(n_1852),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1851),
.A2(n_1415),
.B(n_1412),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1919),
.A2(n_709),
.B1(n_719),
.B2(n_693),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1925),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1816),
.A2(n_719),
.B1(n_693),
.B2(n_694),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1816),
.A2(n_719),
.B1(n_694),
.B2(n_696),
.Y(n_1942)
);

OA21x2_ASAP7_75t_L g1943 ( 
.A1(n_1869),
.A2(n_696),
.B(n_690),
.Y(n_1943)
);

OAI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1851),
.A2(n_708),
.B1(n_711),
.B2(n_704),
.C(n_690),
.Y(n_1944)
);

INVx5_ASAP7_75t_SL g1945 ( 
.A(n_1920),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1808),
.Y(n_1946)
);

NAND2xp33_ASAP7_75t_L g1947 ( 
.A(n_1843),
.B(n_704),
.Y(n_1947)
);

OAI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1787),
.A2(n_711),
.B1(n_713),
.B2(n_708),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1892),
.B(n_1781),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1783),
.A2(n_714),
.B1(n_716),
.B2(n_713),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1783),
.A2(n_716),
.B1(n_717),
.B2(n_714),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1833),
.B(n_1844),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1848),
.B(n_1602),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1786),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1923),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1810),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1843),
.A2(n_726),
.B1(n_717),
.B2(n_579),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1860),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1795),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1866),
.A2(n_726),
.B1(n_581),
.B2(n_586),
.Y(n_1960)
);

OAI21xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1866),
.A2(n_1500),
.B(n_2),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1795),
.Y(n_1962)
);

OAI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1834),
.A2(n_1602),
.B1(n_593),
.B2(n_594),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1781),
.B(n_576),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1921),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1875),
.A2(n_602),
.B1(n_604),
.B2(n_599),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1800),
.A2(n_624),
.B1(n_625),
.B2(n_613),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1921),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1927),
.A2(n_1247),
.B(n_1241),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1819),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1812),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1817),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1854),
.B(n_626),
.Y(n_1973)
);

O2A1O1Ixp33_ASAP7_75t_SL g1974 ( 
.A1(n_1875),
.A2(n_6),
.B(n_2),
.C(n_3),
.Y(n_1974)
);

CKINVDCx11_ASAP7_75t_R g1975 ( 
.A(n_1793),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1800),
.A2(n_635),
.B1(n_637),
.B2(n_634),
.Y(n_1976)
);

AOI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1852),
.A2(n_650),
.B1(n_653),
.B2(n_646),
.C(n_643),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1791),
.A2(n_656),
.B1(n_658),
.B2(n_654),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1835),
.A2(n_670),
.B1(n_667),
.B2(n_1308),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1835),
.A2(n_1308),
.B1(n_441),
.B2(n_448),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1812),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1827),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1882),
.A2(n_441),
.B1(n_453),
.B2(n_436),
.Y(n_1983)
);

BUFx12f_ASAP7_75t_L g1984 ( 
.A(n_1786),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1926),
.A2(n_456),
.B1(n_462),
.B2(n_453),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1824),
.Y(n_1986)
);

OAI221xp5_ASAP7_75t_L g1987 ( 
.A1(n_1889),
.A2(n_465),
.B1(n_466),
.B2(n_462),
.C(n_456),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1833),
.B(n_865),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1824),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1791),
.A2(n_1602),
.B1(n_1500),
.B2(n_466),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1853),
.B(n_7),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1882),
.A2(n_468),
.B1(n_472),
.B2(n_465),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1883),
.B(n_7),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1821),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1777),
.A2(n_472),
.B1(n_478),
.B2(n_468),
.Y(n_1995)
);

OR2x6_ASAP7_75t_L g1996 ( 
.A(n_1788),
.B(n_1388),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1927),
.A2(n_1870),
.B(n_1804),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1831),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_1885),
.Y(n_1999)
);

NAND3xp33_ASAP7_75t_SL g2000 ( 
.A(n_1780),
.B(n_677),
.C(n_478),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1897),
.Y(n_2001)
);

BUFx2_ASAP7_75t_L g2002 ( 
.A(n_1897),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1870),
.A2(n_1262),
.B(n_1475),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1832),
.Y(n_2004)
);

INVx4_ASAP7_75t_L g2005 ( 
.A(n_1845),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1777),
.A2(n_678),
.B1(n_679),
.B2(n_677),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1832),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1859),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1845),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1896),
.B(n_9),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1901),
.A2(n_684),
.B1(n_692),
.B2(n_679),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1856),
.B(n_11),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1784),
.B(n_11),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1829),
.A2(n_692),
.B1(n_697),
.B2(n_684),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1888),
.B(n_905),
.Y(n_2015)
);

OAI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1887),
.A2(n_701),
.B1(n_705),
.B2(n_697),
.Y(n_2016)
);

AND2x6_ASAP7_75t_L g2017 ( 
.A(n_1827),
.B(n_1421),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1806),
.A2(n_705),
.B1(n_706),
.B2(n_701),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1859),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1893),
.B(n_13),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1827),
.Y(n_2021)
);

OR2x6_ASAP7_75t_L g2022 ( 
.A(n_1788),
.B(n_1388),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1867),
.A2(n_715),
.B(n_706),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1874),
.B(n_13),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_1830),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1794),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1804),
.A2(n_1475),
.B(n_1424),
.Y(n_2027)
);

OR2x6_ASAP7_75t_L g2028 ( 
.A(n_1885),
.B(n_1397),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1863),
.A2(n_724),
.B1(n_715),
.B2(n_500),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1865),
.A2(n_724),
.B1(n_502),
.B2(n_503),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1792),
.B(n_14),
.Y(n_2031)
);

AO32x2_ASAP7_75t_L g2032 ( 
.A1(n_1799),
.A2(n_17),
.A3(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1830),
.B(n_16),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1801),
.B(n_17),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1865),
.A2(n_507),
.B1(n_510),
.B2(n_499),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1881),
.B(n_19),
.Y(n_2036)
);

INVxp67_ASAP7_75t_SL g2037 ( 
.A(n_1794),
.Y(n_2037)
);

AOI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_1780),
.A2(n_1836),
.B1(n_1915),
.B2(n_1861),
.C(n_1877),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1797),
.B(n_20),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1840),
.A2(n_514),
.B1(n_518),
.B2(n_513),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1872),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1876),
.A2(n_1424),
.B(n_1421),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1873),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_SL g2044 ( 
.A1(n_1907),
.A2(n_522),
.B1(n_524),
.B2(n_521),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1873),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1837),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1823),
.A2(n_534),
.B1(n_537),
.B2(n_531),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1831),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1910),
.B(n_908),
.Y(n_2049)
);

AOI21xp33_ASAP7_75t_SL g2050 ( 
.A1(n_1811),
.A2(n_20),
.B(n_21),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1874),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1890),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_SL g2053 ( 
.A1(n_1890),
.A2(n_542),
.B1(n_545),
.B2(n_538),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1797),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1789),
.A2(n_551),
.B1(n_557),
.B2(n_546),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1837),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1913),
.B(n_1839),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1899),
.A2(n_1424),
.B(n_1421),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1879),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1823),
.A2(n_566),
.B1(n_577),
.B2(n_562),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1895),
.A2(n_1801),
.B1(n_1924),
.B2(n_1916),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1825),
.B(n_21),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1857),
.A2(n_1785),
.B1(n_1799),
.B2(n_1894),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_1827),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1857),
.A2(n_1884),
.B1(n_1904),
.B2(n_1914),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1899),
.A2(n_1444),
.B(n_1424),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1902),
.B(n_22),
.Y(n_2067)
);

CKINVDCx6p67_ASAP7_75t_R g2068 ( 
.A(n_1850),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1894),
.A2(n_589),
.B1(n_595),
.B2(n_578),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1879),
.B(n_22),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1922),
.A2(n_1928),
.B1(n_1878),
.B2(n_1911),
.Y(n_2071)
);

OR2x6_ASAP7_75t_L g2072 ( 
.A(n_1847),
.B(n_1403),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1880),
.B(n_908),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1922),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1928),
.B(n_23),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_SL g2076 ( 
.A1(n_1905),
.A2(n_598),
.B1(n_600),
.B2(n_596),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_1880),
.B(n_1900),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_R g2078 ( 
.A(n_1846),
.B(n_24),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1900),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1847),
.A2(n_612),
.B1(n_618),
.B2(n_608),
.Y(n_2080)
);

CKINVDCx16_ASAP7_75t_R g2081 ( 
.A(n_1805),
.Y(n_2081)
);

INVx4_ASAP7_75t_SL g2082 ( 
.A(n_1909),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1878),
.A2(n_620),
.B1(n_621),
.B2(n_619),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1782),
.A2(n_629),
.B1(n_630),
.B2(n_627),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1837),
.B(n_24),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1802),
.B(n_25),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1994),
.B(n_1862),
.Y(n_2087)
);

BUFx2_ASAP7_75t_L g2088 ( 
.A(n_2037),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2046),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2004),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2007),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2008),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2019),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2081),
.B(n_1803),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2026),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2043),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1975),
.Y(n_2097)
);

OA21x2_ASAP7_75t_L g2098 ( 
.A1(n_2056),
.A2(n_1779),
.B(n_1818),
.Y(n_2098)
);

AOI21x1_ASAP7_75t_L g2099 ( 
.A1(n_2085),
.A2(n_1905),
.B(n_1855),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1949),
.B(n_1952),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1946),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1932),
.A2(n_1820),
.B(n_1849),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1986),
.Y(n_2103)
);

INVx2_ASAP7_75t_SL g2104 ( 
.A(n_2077),
.Y(n_2104)
);

AO21x2_ASAP7_75t_L g2105 ( 
.A1(n_1997),
.A2(n_1828),
.B(n_1814),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1962),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_2077),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1965),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1931),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1940),
.B(n_1790),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1933),
.Y(n_2111)
);

CKINVDCx20_ASAP7_75t_R g2112 ( 
.A(n_1954),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2045),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1970),
.B(n_1798),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1956),
.Y(n_2115)
);

AO21x2_ASAP7_75t_L g2116 ( 
.A1(n_2042),
.A2(n_1828),
.B(n_1815),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1968),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_L g2118 ( 
.A1(n_2071),
.A2(n_1864),
.B(n_1858),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1972),
.Y(n_2119)
);

NAND2x1p5_ASAP7_75t_L g2120 ( 
.A(n_1999),
.B(n_1905),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2057),
.B(n_1862),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_2064),
.Y(n_2122)
);

OA21x2_ASAP7_75t_L g2123 ( 
.A1(n_1999),
.A2(n_1868),
.B(n_1908),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1959),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2041),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_2025),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_1984),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1971),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2079),
.B(n_1862),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_2051),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1981),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1989),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2059),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2079),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1988),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1929),
.B(n_1903),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2001),
.B(n_1903),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_1958),
.B(n_1813),
.Y(n_2138)
);

INVxp67_ASAP7_75t_L g2139 ( 
.A(n_1937),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_2082),
.B(n_1841),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_L g2141 ( 
.A(n_2078),
.B(n_648),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1937),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2015),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2049),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2002),
.B(n_1903),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2028),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2028),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2028),
.B(n_1813),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_2082),
.B(n_1982),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2073),
.Y(n_2150)
);

INVx1_ASAP7_75t_SL g2151 ( 
.A(n_1998),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_L g2152 ( 
.A1(n_2058),
.A2(n_1842),
.B(n_1838),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_2009),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_1982),
.B(n_1813),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1953),
.B(n_1822),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1943),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1935),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2074),
.B(n_1855),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2074),
.B(n_1855),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2074),
.B(n_1906),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1953),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2021),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_2064),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_2084),
.A2(n_1871),
.B(n_1826),
.Y(n_2164)
);

HB1xp67_ASAP7_75t_L g2165 ( 
.A(n_2021),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_2052),
.Y(n_2166)
);

AO21x2_ASAP7_75t_L g2167 ( 
.A1(n_2084),
.A2(n_1826),
.B(n_1917),
.Y(n_2167)
);

BUFx2_ASAP7_75t_L g2168 ( 
.A(n_2021),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_1964),
.Y(n_2169)
);

AO21x2_ASAP7_75t_L g2170 ( 
.A1(n_2066),
.A2(n_1809),
.B(n_1898),
.Y(n_2170)
);

INVx2_ASAP7_75t_SL g2171 ( 
.A(n_1930),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1943),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2086),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_2065),
.A2(n_1906),
.B(n_1886),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2086),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2024),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2024),
.Y(n_2177)
);

AO21x2_ASAP7_75t_L g2178 ( 
.A1(n_2023),
.A2(n_1912),
.B(n_1906),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1955),
.B(n_26),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2013),
.B(n_27),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2062),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2005),
.B(n_28),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1996),
.Y(n_2183)
);

INVxp67_ASAP7_75t_L g2184 ( 
.A(n_1973),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2063),
.B(n_29),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2034),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2010),
.B(n_29),
.Y(n_2187)
);

BUFx2_ASAP7_75t_L g2188 ( 
.A(n_1996),
.Y(n_2188)
);

AO21x2_ASAP7_75t_L g2189 ( 
.A1(n_2023),
.A2(n_917),
.B(n_913),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2070),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_R g2191 ( 
.A(n_2005),
.B(n_655),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2031),
.B(n_30),
.Y(n_2192)
);

INVxp67_ASAP7_75t_L g2193 ( 
.A(n_2012),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2032),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1993),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2070),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2061),
.B(n_31),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2054),
.B(n_31),
.Y(n_2198)
);

OAI21x1_ASAP7_75t_L g2199 ( 
.A1(n_2027),
.A2(n_1405),
.B(n_1403),
.Y(n_2199)
);

OAI21x1_ASAP7_75t_L g2200 ( 
.A1(n_2035),
.A2(n_1411),
.B(n_1405),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1996),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_1991),
.Y(n_2202)
);

OAI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_1983),
.A2(n_662),
.B(n_657),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2022),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1993),
.Y(n_2205)
);

AO21x2_ASAP7_75t_L g2206 ( 
.A1(n_1983),
.A2(n_917),
.B(n_913),
.Y(n_2206)
);

HB1xp67_ASAP7_75t_L g2207 ( 
.A(n_2022),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2022),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2032),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2032),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2033),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2072),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2067),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_2072),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2072),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2039),
.B(n_32),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2036),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_2048),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2075),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2020),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2017),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_2017),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_1945),
.B(n_33),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2017),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2017),
.Y(n_2225)
);

AO31x2_ASAP7_75t_L g2226 ( 
.A1(n_1990),
.A2(n_939),
.A3(n_942),
.B(n_922),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1961),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1961),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1945),
.B(n_34),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2038),
.Y(n_2230)
);

OA21x2_ASAP7_75t_L g2231 ( 
.A1(n_2083),
.A2(n_939),
.B(n_922),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1974),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2050),
.Y(n_2233)
);

BUFx8_ASAP7_75t_SL g2234 ( 
.A(n_2068),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_2080),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2050),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2003),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_2014),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2060),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2060),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2030),
.B(n_35),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_1934),
.A2(n_1423),
.B(n_1411),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_2076),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1948),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_1992),
.B(n_36),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_1950),
.B(n_1951),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_2053),
.Y(n_2247)
);

BUFx4f_ASAP7_75t_SL g2248 ( 
.A(n_2112),
.Y(n_2248)
);

INVx4_ASAP7_75t_L g2249 ( 
.A(n_2234),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2143),
.B(n_1936),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2090),
.Y(n_2251)
);

AOI22xp33_ASAP7_75t_L g2252 ( 
.A1(n_2230),
.A2(n_1947),
.B1(n_1944),
.B2(n_2000),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2243),
.A2(n_1939),
.B1(n_1942),
.B2(n_1941),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2107),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_2243),
.A2(n_1957),
.B1(n_2018),
.B2(n_1987),
.Y(n_2255)
);

BUFx8_ASAP7_75t_SL g2256 ( 
.A(n_2234),
.Y(n_2256)
);

OAI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_2243),
.A2(n_2016),
.B1(n_1978),
.B2(n_1963),
.Y(n_2257)
);

AOI22xp33_ASAP7_75t_SL g2258 ( 
.A1(n_2141),
.A2(n_1967),
.B1(n_1976),
.B2(n_2040),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2090),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2232),
.A2(n_1985),
.B1(n_1980),
.B2(n_1979),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2141),
.A2(n_2011),
.B(n_1938),
.Y(n_2261)
);

INVx2_ASAP7_75t_SL g2262 ( 
.A(n_2097),
.Y(n_2262)
);

AOI222xp33_ASAP7_75t_L g2263 ( 
.A1(n_2246),
.A2(n_1966),
.B1(n_1960),
.B2(n_1977),
.C1(n_2006),
.C2(n_1995),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_L g2264 ( 
.A1(n_2246),
.A2(n_2044),
.B1(n_2029),
.B2(n_2069),
.Y(n_2264)
);

NAND3xp33_ASAP7_75t_L g2265 ( 
.A(n_2172),
.B(n_2047),
.C(n_2055),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_SL g2266 ( 
.A1(n_2209),
.A2(n_1969),
.B(n_36),
.Y(n_2266)
);

AOI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2239),
.A2(n_942),
.B1(n_947),
.B2(n_1472),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2107),
.Y(n_2268)
);

AOI221xp5_ASAP7_75t_L g2269 ( 
.A1(n_2233),
.A2(n_947),
.B1(n_42),
.B2(n_39),
.C(n_40),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2126),
.Y(n_2270)
);

INVx8_ASAP7_75t_L g2271 ( 
.A(n_2223),
.Y(n_2271)
);

OAI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2239),
.A2(n_1423),
.B1(n_1433),
.B2(n_1428),
.Y(n_2272)
);

OAI211xp5_ASAP7_75t_L g2273 ( 
.A1(n_2233),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2240),
.A2(n_1472),
.B1(n_949),
.B2(n_936),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2240),
.A2(n_1433),
.B1(n_1439),
.B2(n_1428),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2143),
.B(n_43),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2149),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2107),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2089),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2134),
.Y(n_2280)
);

OAI211xp5_ASAP7_75t_L g2281 ( 
.A1(n_2236),
.A2(n_49),
.B(n_46),
.C(n_47),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_SL g2282 ( 
.A1(n_2209),
.A2(n_46),
.B(n_47),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2096),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2236),
.A2(n_1445),
.B1(n_1449),
.B2(n_1439),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2173),
.B(n_52),
.Y(n_2285)
);

INVx4_ASAP7_75t_L g2286 ( 
.A(n_2097),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_SL g2287 ( 
.A1(n_2194),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2134),
.Y(n_2288)
);

AOI21xp33_ASAP7_75t_L g2289 ( 
.A1(n_2227),
.A2(n_57),
.B(n_58),
.Y(n_2289)
);

AOI221xp5_ASAP7_75t_L g2290 ( 
.A1(n_2238),
.A2(n_60),
.B1(n_57),
.B2(n_58),
.C(n_62),
.Y(n_2290)
);

AO31x2_ASAP7_75t_L g2291 ( 
.A1(n_2156),
.A2(n_949),
.A3(n_64),
.B(n_60),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_2189),
.A2(n_1449),
.B(n_1445),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_2112),
.Y(n_2293)
);

AOI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_2228),
.A2(n_921),
.B1(n_923),
.B2(n_920),
.Y(n_2294)
);

AOI21xp33_ASAP7_75t_SL g2295 ( 
.A1(n_2247),
.A2(n_63),
.B(n_65),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_2149),
.Y(n_2296)
);

AOI21xp33_ASAP7_75t_L g2297 ( 
.A1(n_2235),
.A2(n_63),
.B(n_65),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2175),
.B(n_66),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2149),
.B(n_67),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2244),
.A2(n_1472),
.B1(n_69),
.B2(n_67),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2104),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2155),
.B(n_2142),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2126),
.B(n_68),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2182),
.A2(n_884),
.B(n_875),
.Y(n_2304)
);

AOI221xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2194),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.C(n_74),
.Y(n_2305)
);

OAI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2247),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2096),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2104),
.B(n_74),
.Y(n_2308)
);

OAI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2210),
.A2(n_79),
.B1(n_75),
.B2(n_77),
.Y(n_2309)
);

AOI211xp5_ASAP7_75t_L g2310 ( 
.A1(n_2197),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2103),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2168),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_2100),
.B(n_82),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2150),
.B(n_84),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2150),
.B(n_84),
.Y(n_2315)
);

OAI21x1_ASAP7_75t_L g2316 ( 
.A1(n_2089),
.A2(n_1456),
.B(n_1451),
.Y(n_2316)
);

INVx5_ASAP7_75t_SL g2317 ( 
.A(n_2142),
.Y(n_2317)
);

AOI22xp33_ASAP7_75t_L g2318 ( 
.A1(n_2235),
.A2(n_921),
.B1(n_923),
.B2(n_920),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2244),
.A2(n_921),
.B1(n_923),
.B2(n_920),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_SL g2320 ( 
.A1(n_2197),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2189),
.A2(n_921),
.B1(n_923),
.B2(n_920),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2088),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2144),
.B(n_85),
.Y(n_2323)
);

AOI22xp33_ASAP7_75t_L g2324 ( 
.A1(n_2189),
.A2(n_921),
.B1(n_923),
.B2(n_920),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2144),
.B(n_86),
.Y(n_2325)
);

AOI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2139),
.A2(n_1472),
.B1(n_1451),
.B2(n_1469),
.Y(n_2326)
);

INVxp67_ASAP7_75t_L g2327 ( 
.A(n_2088),
.Y(n_2327)
);

AOI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2203),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_2142),
.Y(n_2329)
);

AOI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2241),
.A2(n_1472),
.B1(n_91),
.B2(n_89),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_2117),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2193),
.A2(n_1456),
.B1(n_1473),
.B2(n_1469),
.Y(n_2332)
);

OAI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2245),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_2333)
);

INVx4_ASAP7_75t_L g2334 ( 
.A(n_2166),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2168),
.Y(n_2335)
);

AOI22xp33_ASAP7_75t_L g2336 ( 
.A1(n_2241),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2181),
.A2(n_940),
.B1(n_924),
.B2(n_884),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_L g2338 ( 
.A1(n_2186),
.A2(n_940),
.B1(n_924),
.B2(n_885),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2133),
.Y(n_2339)
);

AOI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_2245),
.A2(n_97),
.B1(n_93),
.B2(n_96),
.Y(n_2340)
);

AOI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2206),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2157),
.B(n_100),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2161),
.B(n_100),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2133),
.Y(n_2344)
);

AOI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2142),
.A2(n_940),
.B1(n_924),
.B2(n_885),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2142),
.A2(n_924),
.B1(n_940),
.B2(n_875),
.Y(n_2346)
);

OAI21x1_ASAP7_75t_L g2347 ( 
.A1(n_2120),
.A2(n_1473),
.B(n_1294),
.Y(n_2347)
);

NOR2x1_ASAP7_75t_SL g2348 ( 
.A(n_2137),
.B(n_1498),
.Y(n_2348)
);

INVx11_ASAP7_75t_L g2349 ( 
.A(n_2218),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2165),
.B(n_102),
.Y(n_2350)
);

OAI22xp33_ASAP7_75t_L g2351 ( 
.A1(n_2195),
.A2(n_2205),
.B1(n_2177),
.B2(n_2190),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_2206),
.A2(n_940),
.B1(n_924),
.B2(n_1211),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2206),
.A2(n_1306),
.B(n_1303),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2176),
.A2(n_1462),
.B1(n_1468),
.B2(n_1417),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_2169),
.A2(n_1211),
.B1(n_1219),
.B2(n_1245),
.Y(n_2355)
);

OAI221xp5_ASAP7_75t_L g2356 ( 
.A1(n_2184),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.C(n_106),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2135),
.B(n_107),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_L g2358 ( 
.A1(n_2185),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2117),
.Y(n_2359)
);

HB1xp67_ASAP7_75t_L g2360 ( 
.A(n_2138),
.Y(n_2360)
);

AOI22xp33_ASAP7_75t_SL g2361 ( 
.A1(n_2185),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2103),
.Y(n_2362)
);

AOI21x1_ASAP7_75t_L g2363 ( 
.A1(n_2162),
.A2(n_1347),
.B(n_1345),
.Y(n_2363)
);

AOI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2237),
.A2(n_1312),
.B(n_1306),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2113),
.Y(n_2365)
);

OAI21x1_ASAP7_75t_L g2366 ( 
.A1(n_2120),
.A2(n_1468),
.B(n_1462),
.Y(n_2366)
);

AOI22xp33_ASAP7_75t_L g2367 ( 
.A1(n_2176),
.A2(n_1211),
.B1(n_1219),
.B2(n_1296),
.Y(n_2367)
);

OAI21x1_ASAP7_75t_L g2368 ( 
.A1(n_2120),
.A2(n_1166),
.B(n_1162),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_2192),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2369)
);

AOI22xp33_ASAP7_75t_L g2370 ( 
.A1(n_2177),
.A2(n_2190),
.B1(n_2196),
.B2(n_2219),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2113),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2135),
.B(n_113),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2196),
.A2(n_2202),
.B1(n_2153),
.B2(n_2188),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2251),
.Y(n_2374)
);

INVx3_ASAP7_75t_L g2375 ( 
.A(n_2277),
.Y(n_2375)
);

HB1xp67_ASAP7_75t_L g2376 ( 
.A(n_2322),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2276),
.B(n_2101),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2283),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2259),
.Y(n_2379)
);

OR2x2_ASAP7_75t_L g2380 ( 
.A(n_2327),
.B(n_2138),
.Y(n_2380)
);

INVxp67_ASAP7_75t_L g2381 ( 
.A(n_2270),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2279),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2307),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2277),
.B(n_2122),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2279),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2322),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2296),
.B(n_2122),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2359),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2311),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2323),
.B(n_2109),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2331),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2296),
.B(n_2122),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2362),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2327),
.B(n_2156),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_2329),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2360),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2302),
.B(n_2312),
.Y(n_2397)
);

INVx4_ASAP7_75t_L g2398 ( 
.A(n_2249),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2331),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2302),
.B(n_2140),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2286),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2325),
.B(n_2111),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2335),
.B(n_2163),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_2360),
.B(n_2339),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2280),
.Y(n_2405)
);

BUFx2_ASAP7_75t_L g2406 ( 
.A(n_2286),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2373),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2254),
.B(n_2163),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2268),
.B(n_2163),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2288),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2344),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2250),
.B(n_2119),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2348),
.B(n_2140),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2278),
.B(n_2171),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2365),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2371),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2314),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2315),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2303),
.B(n_2211),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2334),
.Y(n_2420)
);

BUFx3_ASAP7_75t_L g2421 ( 
.A(n_2256),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_2249),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2301),
.B(n_2171),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2317),
.B(n_2121),
.Y(n_2424)
);

INVx4_ASAP7_75t_L g2425 ( 
.A(n_2299),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2257),
.A2(n_2237),
.B1(n_2153),
.B2(n_2231),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2317),
.B(n_2121),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2357),
.B(n_2213),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2317),
.B(n_2136),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2291),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2370),
.B(n_2136),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2291),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2262),
.B(n_2222),
.Y(n_2433)
);

AND2x4_ASAP7_75t_SL g2434 ( 
.A(n_2334),
.B(n_2183),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2313),
.B(n_2137),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2342),
.B(n_2145),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2308),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2372),
.B(n_2217),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2351),
.B(n_2091),
.Y(n_2439)
);

OAI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2255),
.A2(n_2188),
.B1(n_2183),
.B2(n_2094),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2291),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2350),
.B(n_2343),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2299),
.B(n_2145),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2291),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2271),
.Y(n_2445)
);

BUFx2_ASAP7_75t_L g2446 ( 
.A(n_2271),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2351),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2271),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2285),
.Y(n_2449)
);

OR2x2_ASAP7_75t_L g2450 ( 
.A(n_2366),
.B(n_2092),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2298),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2248),
.B(n_2127),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_SL g2453 ( 
.A1(n_2260),
.A2(n_2229),
.B1(n_2223),
.B2(n_2198),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2293),
.B(n_2130),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2266),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2363),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2305),
.B(n_2115),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2347),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2282),
.Y(n_2459)
);

INVx2_ASAP7_75t_SL g2460 ( 
.A(n_2349),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_2316),
.B(n_2140),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2368),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2332),
.Y(n_2463)
);

NAND2x1p5_ASAP7_75t_SL g2464 ( 
.A(n_2310),
.B(n_2229),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2284),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2354),
.Y(n_2466)
);

HB1xp67_ASAP7_75t_L g2467 ( 
.A(n_2272),
.Y(n_2467)
);

BUFx12f_ASAP7_75t_L g2468 ( 
.A(n_2248),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2309),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2265),
.B(n_2093),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2309),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2275),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2257),
.B(n_2125),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2304),
.B(n_2146),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2364),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2356),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_2261),
.B(n_2146),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2333),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2326),
.Y(n_2479)
);

CKINVDCx20_ASAP7_75t_R g2480 ( 
.A(n_2297),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2255),
.A2(n_2231),
.B1(n_2220),
.B2(n_2167),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2287),
.B(n_2147),
.Y(n_2482)
);

OR2x2_ASAP7_75t_L g2483 ( 
.A(n_2337),
.B(n_2095),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2295),
.Y(n_2484)
);

OAI21xp5_ASAP7_75t_SL g2485 ( 
.A1(n_2252),
.A2(n_2198),
.B(n_2187),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2287),
.B(n_2147),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2481),
.A2(n_2426),
.B(n_2440),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2484),
.B(n_2216),
.Y(n_2488)
);

HB1xp67_ASAP7_75t_L g2489 ( 
.A(n_2396),
.Y(n_2489)
);

INVxp67_ASAP7_75t_SL g2490 ( 
.A(n_2376),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2484),
.B(n_2216),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2378),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2386),
.Y(n_2493)
);

NAND4xp25_ASAP7_75t_SL g2494 ( 
.A(n_2453),
.B(n_2253),
.C(n_2328),
.D(n_2290),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2375),
.Y(n_2495)
);

OAI221xp5_ASAP7_75t_L g2496 ( 
.A1(n_2485),
.A2(n_2476),
.B1(n_2407),
.B2(n_2470),
.C(n_2473),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2378),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2375),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2406),
.B(n_2127),
.Y(n_2499)
);

NOR2x1_ASAP7_75t_SL g2500 ( 
.A(n_2443),
.B(n_2273),
.Y(n_2500)
);

OAI31xp33_ASAP7_75t_L g2501 ( 
.A1(n_2469),
.A2(n_2306),
.A3(n_2333),
.B(n_2281),
.Y(n_2501)
);

NAND4xp25_ASAP7_75t_SL g2502 ( 
.A(n_2471),
.B(n_2253),
.C(n_2252),
.D(n_2269),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2389),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2375),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2389),
.Y(n_2505)
);

BUFx3_ASAP7_75t_L g2506 ( 
.A(n_2421),
.Y(n_2506)
);

OAI31xp33_ASAP7_75t_L g2507 ( 
.A1(n_2478),
.A2(n_2306),
.A3(n_2289),
.B(n_2358),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2401),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2374),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2401),
.Y(n_2510)
);

AND2x4_ASAP7_75t_L g2511 ( 
.A(n_2406),
.B(n_2166),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2401),
.Y(n_2512)
);

NOR4xp25_ASAP7_75t_SL g2513 ( 
.A(n_2395),
.B(n_2224),
.C(n_2108),
.D(n_2106),
.Y(n_2513)
);

OAI33xp33_ASAP7_75t_L g2514 ( 
.A1(n_2457),
.A2(n_2180),
.A3(n_2320),
.B1(n_2361),
.B2(n_2114),
.B3(n_2340),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2459),
.B(n_2216),
.Y(n_2515)
);

OAI31xp33_ASAP7_75t_L g2516 ( 
.A1(n_2476),
.A2(n_2358),
.A3(n_2340),
.B(n_2336),
.Y(n_2516)
);

INVxp67_ASAP7_75t_SL g2517 ( 
.A(n_2381),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_R g2518 ( 
.A(n_2420),
.B(n_2231),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2459),
.B(n_2179),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2468),
.Y(n_2520)
);

CKINVDCx20_ASAP7_75t_R g2521 ( 
.A(n_2421),
.Y(n_2521)
);

AOI211xp5_ASAP7_75t_L g2522 ( 
.A1(n_2470),
.A2(n_2191),
.B(n_2180),
.C(n_2179),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2425),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2443),
.B(n_2218),
.Y(n_2524)
);

AOI221xp5_ASAP7_75t_L g2525 ( 
.A1(n_2464),
.A2(n_2336),
.B1(n_2369),
.B2(n_2320),
.C(n_2361),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2446),
.B(n_2207),
.Y(n_2526)
);

OAI33xp33_ASAP7_75t_L g2527 ( 
.A1(n_2430),
.A2(n_2106),
.A3(n_2108),
.B1(n_2110),
.B2(n_2369),
.B3(n_2154),
.Y(n_2527)
);

OAI211xp5_ASAP7_75t_L g2528 ( 
.A1(n_2480),
.A2(n_2264),
.B(n_2263),
.C(n_2258),
.Y(n_2528)
);

BUFx2_ASAP7_75t_L g2529 ( 
.A(n_2420),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_L g2530 ( 
.A1(n_2480),
.A2(n_2264),
.B1(n_2258),
.B2(n_2330),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_SL g2531 ( 
.A1(n_2482),
.A2(n_2105),
.B1(n_2178),
.B2(n_2151),
.Y(n_2531)
);

NAND3xp33_ASAP7_75t_L g2532 ( 
.A(n_2475),
.B(n_2341),
.C(n_2330),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2455),
.B(n_2318),
.Y(n_2533)
);

OAI321xp33_ASAP7_75t_L g2534 ( 
.A1(n_2447),
.A2(n_2341),
.A3(n_2300),
.B1(n_2319),
.B2(n_2294),
.C(n_2148),
.Y(n_2534)
);

OAI22xp5_ASAP7_75t_L g2535 ( 
.A1(n_2446),
.A2(n_2300),
.B1(n_2183),
.B2(n_2148),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2398),
.B(n_2131),
.Y(n_2536)
);

OA21x2_ASAP7_75t_L g2537 ( 
.A1(n_2395),
.A2(n_2118),
.B(n_2102),
.Y(n_2537)
);

BUFx2_ASAP7_75t_L g2538 ( 
.A(n_2425),
.Y(n_2538)
);

AOI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2477),
.A2(n_2167),
.B(n_2105),
.Y(n_2539)
);

AO21x2_ASAP7_75t_L g2540 ( 
.A1(n_2382),
.A2(n_2353),
.B(n_2292),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2379),
.Y(n_2541)
);

NAND2xp33_ASAP7_75t_R g2542 ( 
.A(n_2477),
.B(n_114),
.Y(n_2542)
);

OAI21xp5_ASAP7_75t_SL g2543 ( 
.A1(n_2482),
.A2(n_2324),
.B(n_2321),
.Y(n_2543)
);

AOI21xp5_ASAP7_75t_L g2544 ( 
.A1(n_2477),
.A2(n_2486),
.B(n_2467),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2417),
.B(n_2132),
.Y(n_2545)
);

AOI22xp33_ASAP7_75t_L g2546 ( 
.A1(n_2486),
.A2(n_2167),
.B1(n_2105),
.B2(n_2164),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_2468),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2383),
.Y(n_2548)
);

NAND4xp25_ASAP7_75t_L g2549 ( 
.A(n_2398),
.B(n_2338),
.C(n_2346),
.D(n_2345),
.Y(n_2549)
);

NAND2xp33_ASAP7_75t_R g2550 ( 
.A(n_2452),
.B(n_114),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_R g2551 ( 
.A(n_2422),
.B(n_116),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2412),
.B(n_2124),
.Y(n_2552)
);

OAI221xp5_ASAP7_75t_L g2553 ( 
.A1(n_2398),
.A2(n_2204),
.B1(n_2201),
.B2(n_2208),
.C(n_2214),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_R g2554 ( 
.A(n_2422),
.B(n_117),
.Y(n_2554)
);

AOI221xp5_ASAP7_75t_SL g2555 ( 
.A1(n_2397),
.A2(n_2221),
.B1(n_2225),
.B2(n_2208),
.C(n_2201),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2433),
.B(n_2204),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2393),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2430),
.A2(n_2178),
.B(n_2164),
.Y(n_2558)
);

AO21x2_ASAP7_75t_L g2559 ( 
.A1(n_2382),
.A2(n_2225),
.B(n_2221),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2433),
.B(n_2155),
.Y(n_2560)
);

AOI221xp5_ASAP7_75t_L g2561 ( 
.A1(n_2464),
.A2(n_2087),
.B1(n_2124),
.B2(n_2128),
.C(n_2155),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2425),
.Y(n_2562)
);

AOI221xp5_ASAP7_75t_L g2563 ( 
.A1(n_2466),
.A2(n_2087),
.B1(n_2128),
.B2(n_2159),
.C(n_2352),
.Y(n_2563)
);

AOI211xp5_ASAP7_75t_L g2564 ( 
.A1(n_2422),
.A2(n_2212),
.B(n_2215),
.C(n_2160),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2384),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2397),
.B(n_2212),
.Y(n_2566)
);

AO21x2_ASAP7_75t_L g2567 ( 
.A1(n_2385),
.A2(n_2399),
.B(n_2391),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2418),
.B(n_2159),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2436),
.B(n_2448),
.Y(n_2569)
);

OA21x2_ASAP7_75t_L g2570 ( 
.A1(n_2448),
.A2(n_2118),
.B(n_2102),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2385),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2437),
.B(n_2160),
.Y(n_2572)
);

NAND2xp33_ASAP7_75t_R g2573 ( 
.A(n_2439),
.B(n_117),
.Y(n_2573)
);

AOI33xp33_ASAP7_75t_L g2574 ( 
.A1(n_2472),
.A2(n_2215),
.A3(n_2129),
.B1(n_2267),
.B2(n_2274),
.B3(n_2355),
.Y(n_2574)
);

AOI211xp5_ASAP7_75t_L g2575 ( 
.A1(n_2528),
.A2(n_2422),
.B(n_2445),
.C(n_2439),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2489),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2511),
.B(n_2524),
.Y(n_2577)
);

NAND3xp33_ASAP7_75t_L g2578 ( 
.A(n_2573),
.B(n_2422),
.C(n_2432),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2511),
.B(n_2445),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2529),
.Y(n_2580)
);

AO21x2_ASAP7_75t_L g2581 ( 
.A1(n_2544),
.A2(n_2399),
.B(n_2391),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2517),
.B(n_2449),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2489),
.Y(n_2583)
);

NOR2x1_ASAP7_75t_L g2584 ( 
.A(n_2528),
.B(n_2454),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2517),
.B(n_2437),
.Y(n_2585)
);

NOR2x1_ASAP7_75t_L g2586 ( 
.A(n_2494),
.B(n_2454),
.Y(n_2586)
);

NAND3xp33_ASAP7_75t_L g2587 ( 
.A(n_2573),
.B(n_2444),
.C(n_2441),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2500),
.B(n_2530),
.Y(n_2588)
);

NAND4xp75_ASAP7_75t_L g2589 ( 
.A(n_2487),
.B(n_2460),
.C(n_2429),
.D(n_2427),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2506),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2493),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2499),
.B(n_2435),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2499),
.B(n_2435),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2547),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2493),
.Y(n_2595)
);

NAND3xp33_ASAP7_75t_L g2596 ( 
.A(n_2525),
.B(n_2456),
.C(n_2483),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2530),
.B(n_2479),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2521),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2569),
.B(n_2566),
.Y(n_2599)
);

AO21x1_ASAP7_75t_SL g2600 ( 
.A1(n_2515),
.A2(n_2463),
.B(n_2442),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2538),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2526),
.B(n_2436),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2501),
.B(n_2507),
.Y(n_2603)
);

OA211x2_ASAP7_75t_L g2604 ( 
.A1(n_2502),
.A2(n_2377),
.B(n_2402),
.C(n_2390),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2556),
.B(n_2434),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2544),
.B(n_2479),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2568),
.B(n_2465),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2565),
.B(n_2434),
.Y(n_2608)
);

NAND4xp75_ASAP7_75t_L g2609 ( 
.A(n_2516),
.B(n_2460),
.C(n_2429),
.D(n_2427),
.Y(n_2609)
);

BUFx6f_ASAP7_75t_L g2610 ( 
.A(n_2520),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_2533),
.B(n_2419),
.Y(n_2611)
);

NOR3xp33_ASAP7_75t_L g2612 ( 
.A(n_2496),
.B(n_2438),
.C(n_2428),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2514),
.B(n_2451),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2523),
.B(n_2400),
.Y(n_2614)
);

AND2x4_ASAP7_75t_L g2615 ( 
.A(n_2562),
.B(n_2400),
.Y(n_2615)
);

OAI221xp5_ASAP7_75t_SL g2616 ( 
.A1(n_2543),
.A2(n_2431),
.B1(n_2380),
.B2(n_2483),
.C(n_2474),
.Y(n_2616)
);

NOR3xp33_ASAP7_75t_L g2617 ( 
.A(n_2514),
.B(n_2534),
.C(n_2532),
.Y(n_2617)
);

NAND4xp25_ASAP7_75t_L g2618 ( 
.A(n_2550),
.B(n_2431),
.C(n_2380),
.D(n_2394),
.Y(n_2618)
);

AOI221xp5_ASAP7_75t_L g2619 ( 
.A1(n_2527),
.A2(n_2474),
.B1(n_2415),
.B2(n_2411),
.C(n_2416),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2572),
.B(n_2394),
.Y(n_2620)
);

NAND3xp33_ASAP7_75t_SL g2621 ( 
.A(n_2531),
.B(n_2522),
.C(n_2513),
.Y(n_2621)
);

NAND3xp33_ASAP7_75t_L g2622 ( 
.A(n_2542),
.B(n_2404),
.C(n_2267),
.Y(n_2622)
);

NAND3xp33_ASAP7_75t_L g2623 ( 
.A(n_2542),
.B(n_2404),
.C(n_2411),
.Y(n_2623)
);

AOI211x1_ASAP7_75t_L g2624 ( 
.A1(n_2535),
.A2(n_2384),
.B(n_2392),
.C(n_2387),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2490),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2490),
.B(n_2400),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2560),
.B(n_2424),
.Y(n_2627)
);

NAND3xp33_ASAP7_75t_L g2628 ( 
.A(n_2531),
.B(n_2415),
.C(n_2416),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2488),
.B(n_2388),
.Y(n_2629)
);

OA211x2_ASAP7_75t_L g2630 ( 
.A1(n_2561),
.A2(n_2387),
.B(n_2392),
.C(n_2274),
.Y(n_2630)
);

OAI211xp5_ASAP7_75t_L g2631 ( 
.A1(n_2551),
.A2(n_2424),
.B(n_2458),
.C(n_2403),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2567),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2546),
.A2(n_2413),
.B1(n_2423),
.B2(n_2458),
.Y(n_2633)
);

AOI21xp33_ASAP7_75t_L g2634 ( 
.A1(n_2518),
.A2(n_2450),
.B(n_2462),
.Y(n_2634)
);

NAND3xp33_ASAP7_75t_L g2635 ( 
.A(n_2546),
.B(n_2388),
.C(n_2405),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2527),
.A2(n_2555),
.B1(n_2536),
.B2(n_2491),
.Y(n_2636)
);

NOR3xp33_ASAP7_75t_L g2637 ( 
.A(n_2549),
.B(n_2403),
.C(n_2462),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2508),
.B(n_2423),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2519),
.B(n_2414),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2492),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2510),
.B(n_2512),
.Y(n_2641)
);

OA211x2_ASAP7_75t_L g2642 ( 
.A1(n_2536),
.A2(n_2413),
.B(n_2408),
.C(n_2409),
.Y(n_2642)
);

NAND4xp75_ASAP7_75t_L g2643 ( 
.A(n_2539),
.B(n_2409),
.C(n_2408),
.D(n_2414),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2564),
.B(n_2413),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2574),
.B(n_2405),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2495),
.B(n_2498),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2504),
.B(n_2410),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_SL g2648 ( 
.A1(n_2554),
.A2(n_2540),
.B1(n_2553),
.B2(n_2567),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2563),
.A2(n_2461),
.B1(n_2410),
.B2(n_2450),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2571),
.B(n_2461),
.Y(n_2650)
);

NAND3xp33_ASAP7_75t_L g2651 ( 
.A(n_2518),
.B(n_2461),
.C(n_2367),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2497),
.Y(n_2652)
);

OAI211xp5_ASAP7_75t_SL g2653 ( 
.A1(n_2558),
.A2(n_2158),
.B(n_2154),
.C(n_120),
.Y(n_2653)
);

NAND4xp25_ASAP7_75t_L g2654 ( 
.A(n_2509),
.B(n_2158),
.C(n_2129),
.D(n_121),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2503),
.Y(n_2655)
);

NAND3xp33_ASAP7_75t_L g2656 ( 
.A(n_2558),
.B(n_2098),
.C(n_118),
.Y(n_2656)
);

NAND3xp33_ASAP7_75t_L g2657 ( 
.A(n_2617),
.B(n_2548),
.C(n_2541),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2583),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2581),
.Y(n_2659)
);

HB1xp67_ASAP7_75t_L g2660 ( 
.A(n_2580),
.Y(n_2660)
);

BUFx2_ASAP7_75t_L g2661 ( 
.A(n_2581),
.Y(n_2661)
);

NAND3xp33_ASAP7_75t_L g2662 ( 
.A(n_2578),
.B(n_2557),
.C(n_2505),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2602),
.B(n_2559),
.Y(n_2663)
);

AOI33xp33_ASAP7_75t_L g2664 ( 
.A1(n_2575),
.A2(n_2539),
.A3(n_2540),
.B1(n_2537),
.B2(n_2559),
.B3(n_2545),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2626),
.Y(n_2665)
);

OAI31xp33_ASAP7_75t_L g2666 ( 
.A1(n_2578),
.A2(n_2552),
.A3(n_2537),
.B(n_2570),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2610),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2584),
.B(n_2570),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2626),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2632),
.Y(n_2670)
);

NOR3xp33_ASAP7_75t_L g2671 ( 
.A(n_2603),
.B(n_2200),
.C(n_2174),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2575),
.B(n_2164),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2598),
.Y(n_2673)
);

AND2x4_ASAP7_75t_L g2674 ( 
.A(n_2623),
.B(n_2174),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2615),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2615),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2586),
.B(n_2226),
.Y(n_2677)
);

OAI221xp5_ASAP7_75t_L g2678 ( 
.A1(n_2588),
.A2(n_2098),
.B1(n_2099),
.B2(n_2123),
.C(n_2226),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2577),
.B(n_2098),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2601),
.B(n_2226),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2625),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2610),
.B(n_119),
.Y(n_2682)
);

OAI211xp5_ASAP7_75t_L g2683 ( 
.A1(n_2621),
.A2(n_2099),
.B(n_2123),
.C(n_2199),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2576),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2594),
.B(n_2644),
.Y(n_2685)
);

AOI221xp5_ASAP7_75t_L g2686 ( 
.A1(n_2596),
.A2(n_2178),
.B1(n_2116),
.B2(n_2170),
.C(n_126),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2591),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2595),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2605),
.B(n_2226),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2590),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2587),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2613),
.B(n_2618),
.Y(n_2692)
);

AOI33xp33_ASAP7_75t_L g2693 ( 
.A1(n_2648),
.A2(n_119),
.A3(n_122),
.B1(n_123),
.B2(n_126),
.B3(n_129),
.Y(n_2693)
);

HB1xp67_ASAP7_75t_L g2694 ( 
.A(n_2582),
.Y(n_2694)
);

OR2x2_ASAP7_75t_L g2695 ( 
.A(n_2623),
.B(n_2226),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2618),
.B(n_122),
.Y(n_2696)
);

NAND4xp25_ASAP7_75t_L g2697 ( 
.A(n_2604),
.B(n_134),
.C(n_129),
.D(n_132),
.Y(n_2697)
);

AOI33xp33_ASAP7_75t_L g2698 ( 
.A1(n_2649),
.A2(n_132),
.A3(n_134),
.B1(n_135),
.B2(n_136),
.B3(n_140),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2592),
.Y(n_2699)
);

OAI33xp33_ASAP7_75t_L g2700 ( 
.A1(n_2587),
.A2(n_140),
.A3(n_144),
.B1(n_145),
.B2(n_147),
.B3(n_148),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2585),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2593),
.Y(n_2702)
);

OAI221xp5_ASAP7_75t_L g2703 ( 
.A1(n_2596),
.A2(n_2616),
.B1(n_2636),
.B2(n_2612),
.C(n_2597),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2640),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2606),
.B(n_145),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2620),
.B(n_2116),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2610),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2645),
.B(n_2116),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2599),
.B(n_2123),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2627),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2609),
.B(n_149),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2652),
.Y(n_2712)
);

OAI21x1_ASAP7_75t_L g2713 ( 
.A1(n_2628),
.A2(n_2199),
.B(n_2152),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2579),
.B(n_2170),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2614),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2608),
.B(n_2170),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2655),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2641),
.B(n_149),
.Y(n_2718)
);

INVx2_ASAP7_75t_SL g2719 ( 
.A(n_2667),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2661),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2692),
.A2(n_2628),
.B(n_2656),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2661),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_L g2723 ( 
.A1(n_2703),
.A2(n_2630),
.B1(n_2656),
.B2(n_2642),
.Y(n_2723)
);

AOI21x1_ASAP7_75t_L g2724 ( 
.A1(n_2659),
.A2(n_2631),
.B(n_2633),
.Y(n_2724)
);

OR2x2_ASAP7_75t_SL g2725 ( 
.A(n_2660),
.B(n_2665),
.Y(n_2725)
);

HB1xp67_ASAP7_75t_L g2726 ( 
.A(n_2659),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2673),
.B(n_2611),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2707),
.B(n_2589),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2707),
.B(n_2600),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2707),
.B(n_2638),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2691),
.B(n_2622),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2697),
.A2(n_2653),
.B1(n_2637),
.B2(n_2622),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2658),
.Y(n_2733)
);

OAI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2668),
.A2(n_2654),
.B1(n_2651),
.B2(n_2635),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2658),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2670),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2665),
.B(n_2646),
.Y(n_2737)
);

INVxp67_ASAP7_75t_L g2738 ( 
.A(n_2691),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2667),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2670),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2681),
.Y(n_2741)
);

AOI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2686),
.A2(n_2643),
.B1(n_2639),
.B2(n_2651),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2685),
.B(n_2607),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2681),
.Y(n_2744)
);

AOI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2711),
.A2(n_2650),
.B1(n_2635),
.B2(n_2619),
.Y(n_2745)
);

INVx1_ASAP7_75t_SL g2746 ( 
.A(n_2685),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2696),
.A2(n_2647),
.B1(n_2629),
.B2(n_2634),
.Y(n_2747)
);

OAI22xp33_ASAP7_75t_L g2748 ( 
.A1(n_2677),
.A2(n_2624),
.B1(n_151),
.B2(n_152),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2684),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_SL g2750 ( 
.A(n_2700),
.B(n_150),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2669),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2684),
.Y(n_2752)
);

OAI322xp33_ASAP7_75t_L g2753 ( 
.A1(n_2657),
.A2(n_2695),
.A3(n_2672),
.B1(n_2708),
.B2(n_2662),
.C1(n_2701),
.C2(n_2688),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2687),
.Y(n_2754)
);

NAND2x1_ASAP7_75t_SL g2755 ( 
.A(n_2663),
.B(n_151),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2687),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2673),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2710),
.B(n_152),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2669),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2675),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2693),
.B(n_154),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2710),
.B(n_2699),
.Y(n_2762)
);

NOR2xp33_ASAP7_75t_L g2763 ( 
.A(n_2690),
.B(n_154),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2675),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2676),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2746),
.B(n_2676),
.Y(n_2766)
);

INVxp67_ASAP7_75t_L g2767 ( 
.A(n_2728),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2746),
.B(n_2699),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2726),
.Y(n_2769)
);

OR2x2_ASAP7_75t_L g2770 ( 
.A(n_2725),
.B(n_2690),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2719),
.B(n_2702),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_2721),
.B(n_2664),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2743),
.B(n_2702),
.Y(n_2773)
);

NAND2xp33_ASAP7_75t_L g2774 ( 
.A(n_2731),
.B(n_2705),
.Y(n_2774)
);

INVx1_ASAP7_75t_SL g2775 ( 
.A(n_2755),
.Y(n_2775)
);

AOI21xp33_ASAP7_75t_L g2776 ( 
.A1(n_2731),
.A2(n_2694),
.B(n_2708),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2726),
.Y(n_2777)
);

NAND4xp25_ASAP7_75t_L g2778 ( 
.A(n_2723),
.B(n_2715),
.C(n_2701),
.D(n_2698),
.Y(n_2778)
);

INVx1_ASAP7_75t_SL g2779 ( 
.A(n_2729),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2721),
.B(n_2715),
.Y(n_2780)
);

OR2x2_ASAP7_75t_L g2781 ( 
.A(n_2727),
.B(n_2751),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2737),
.B(n_2718),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2737),
.B(n_2682),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2730),
.B(n_2663),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2760),
.B(n_2704),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2739),
.B(n_2704),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2762),
.B(n_2689),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2759),
.B(n_2712),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2732),
.B(n_2712),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2758),
.B(n_2689),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2764),
.B(n_2717),
.Y(n_2791)
);

NAND2xp33_ASAP7_75t_SL g2792 ( 
.A(n_2761),
.B(n_2695),
.Y(n_2792)
);

OR2x2_ASAP7_75t_L g2793 ( 
.A(n_2765),
.B(n_2717),
.Y(n_2793)
);

BUFx2_ASAP7_75t_L g2794 ( 
.A(n_2757),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2720),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2722),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2747),
.B(n_2716),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2736),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2740),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2733),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2745),
.B(n_2680),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2738),
.B(n_2714),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2738),
.Y(n_2803)
);

NOR2xp67_ASAP7_75t_L g2804 ( 
.A(n_2770),
.B(n_2735),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2773),
.B(n_2763),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2784),
.B(n_2734),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2772),
.B(n_2749),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2768),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2775),
.B(n_2742),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2768),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2779),
.B(n_2767),
.Y(n_2811)
);

AND4x1_ASAP7_75t_L g2812 ( 
.A(n_2780),
.B(n_2750),
.C(n_2761),
.D(n_2754),
.Y(n_2812)
);

NAND2x1p5_ASAP7_75t_L g2813 ( 
.A(n_2794),
.B(n_2752),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2803),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2790),
.B(n_2756),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2772),
.B(n_2741),
.Y(n_2816)
);

OR2x2_ASAP7_75t_L g2817 ( 
.A(n_2766),
.B(n_2748),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2780),
.B(n_2748),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2803),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2769),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2777),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2788),
.B(n_2744),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2787),
.B(n_2724),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2778),
.B(n_2750),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2771),
.B(n_2716),
.Y(n_2825)
);

NAND3xp33_ASAP7_75t_L g2826 ( 
.A(n_2774),
.B(n_2666),
.C(n_2683),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2788),
.B(n_2674),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2797),
.B(n_2714),
.Y(n_2828)
);

NAND4xp25_ASAP7_75t_L g2829 ( 
.A(n_2789),
.B(n_2753),
.C(n_2674),
.D(n_2671),
.Y(n_2829)
);

NOR2xp67_ASAP7_75t_SL g2830 ( 
.A(n_2781),
.B(n_2706),
.Y(n_2830)
);

AOI211xp5_ASAP7_75t_L g2831 ( 
.A1(n_2776),
.A2(n_2674),
.B(n_2678),
.C(n_2713),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2783),
.B(n_2679),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2791),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2782),
.B(n_2679),
.Y(n_2834)
);

OR2x2_ASAP7_75t_L g2835 ( 
.A(n_2786),
.B(n_2706),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_R g2836 ( 
.A1(n_2812),
.A2(n_2788),
.B(n_2792),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2813),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2813),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2826),
.A2(n_2801),
.B1(n_2785),
.B2(n_2793),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2808),
.B(n_2791),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2805),
.B(n_2802),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2810),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2827),
.Y(n_2843)
);

A2O1A1Ixp33_ASAP7_75t_L g2844 ( 
.A1(n_2824),
.A2(n_2792),
.B(n_2774),
.C(n_2796),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2814),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2827),
.Y(n_2846)
);

OAI22xp33_ASAP7_75t_L g2847 ( 
.A1(n_2829),
.A2(n_2817),
.B1(n_2816),
.B2(n_2807),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2819),
.Y(n_2848)
);

HB1xp67_ASAP7_75t_L g2849 ( 
.A(n_2804),
.Y(n_2849)
);

NOR4xp25_ASAP7_75t_L g2850 ( 
.A(n_2807),
.B(n_2795),
.C(n_2799),
.D(n_2798),
.Y(n_2850)
);

OR2x2_ASAP7_75t_L g2851 ( 
.A(n_2809),
.B(n_2800),
.Y(n_2851)
);

OAI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2829),
.A2(n_2802),
.B1(n_2709),
.B2(n_2713),
.Y(n_2852)
);

OAI221xp5_ASAP7_75t_L g2853 ( 
.A1(n_2818),
.A2(n_2709),
.B1(n_156),
.B2(n_157),
.C(n_158),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2833),
.Y(n_2854)
);

OR2x2_ASAP7_75t_L g2855 ( 
.A(n_2806),
.B(n_155),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2816),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2815),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2831),
.A2(n_2200),
.B(n_2242),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_SL g2859 ( 
.A1(n_2822),
.A2(n_160),
.B(n_162),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2822),
.Y(n_2860)
);

XOR2xp5_ASAP7_75t_L g2861 ( 
.A(n_2839),
.B(n_2851),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2849),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2841),
.Y(n_2863)
);

INVxp67_ASAP7_75t_SL g2864 ( 
.A(n_2840),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2857),
.B(n_2811),
.Y(n_2865)
);

BUFx3_ASAP7_75t_L g2866 ( 
.A(n_2837),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2840),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2855),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2838),
.Y(n_2869)
);

AOI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2847),
.A2(n_2823),
.B1(n_2832),
.B2(n_2834),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2844),
.A2(n_2839),
.B(n_2859),
.Y(n_2871)
);

NOR4xp25_ASAP7_75t_L g2872 ( 
.A(n_2860),
.B(n_2820),
.C(n_2821),
.D(n_2825),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2845),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2848),
.B(n_2842),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2854),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2843),
.B(n_2835),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2846),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2836),
.B(n_2828),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2850),
.B(n_2830),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2866),
.Y(n_2880)
);

NAND2xp33_ASAP7_75t_SL g2881 ( 
.A(n_2879),
.B(n_2856),
.Y(n_2881)
);

AOI21xp33_ASAP7_75t_SL g2882 ( 
.A1(n_2863),
.A2(n_2853),
.B(n_2852),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2862),
.Y(n_2883)
);

OAI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2871),
.A2(n_2853),
.B(n_2856),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2865),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2861),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2876),
.Y(n_2887)
);

OAI32xp33_ASAP7_75t_L g2888 ( 
.A1(n_2869),
.A2(n_2858),
.A3(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2864),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2876),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2878),
.B(n_160),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2878),
.B(n_164),
.Y(n_2892)
);

NOR2x1_ASAP7_75t_L g2893 ( 
.A(n_2890),
.B(n_2887),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2891),
.Y(n_2894)
);

NOR2x1_ASAP7_75t_L g2895 ( 
.A(n_2880),
.B(n_2868),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2892),
.B(n_2870),
.Y(n_2896)
);

OAI211xp5_ASAP7_75t_SL g2897 ( 
.A1(n_2884),
.A2(n_2870),
.B(n_2867),
.C(n_2877),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2880),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2882),
.B(n_2872),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2885),
.B(n_2872),
.Y(n_2900)
);

OAI21xp5_ASAP7_75t_SL g2901 ( 
.A1(n_2884),
.A2(n_2874),
.B(n_2873),
.Y(n_2901)
);

OAI21xp33_ASAP7_75t_L g2902 ( 
.A1(n_2886),
.A2(n_2875),
.B(n_2242),
.Y(n_2902)
);

AOI211xp5_ASAP7_75t_L g2903 ( 
.A1(n_2888),
.A2(n_165),
.B(n_166),
.C(n_167),
.Y(n_2903)
);

NOR3xp33_ASAP7_75t_L g2904 ( 
.A(n_2881),
.B(n_168),
.C(n_169),
.Y(n_2904)
);

OR2x2_ASAP7_75t_L g2905 ( 
.A(n_2883),
.B(n_168),
.Y(n_2905)
);

AOI22xp33_ASAP7_75t_L g2906 ( 
.A1(n_2899),
.A2(n_2881),
.B1(n_2889),
.B2(n_2152),
.Y(n_2906)
);

BUFx3_ASAP7_75t_L g2907 ( 
.A(n_2894),
.Y(n_2907)
);

NAND2xp33_ASAP7_75t_SL g2908 ( 
.A(n_2896),
.B(n_169),
.Y(n_2908)
);

OR2x2_ASAP7_75t_L g2909 ( 
.A(n_2900),
.B(n_2898),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2893),
.B(n_170),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2905),
.Y(n_2911)
);

OAI21xp5_ASAP7_75t_SL g2912 ( 
.A1(n_2897),
.A2(n_172),
.B(n_173),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2904),
.B(n_174),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2895),
.Y(n_2914)
);

AOI221xp5_ASAP7_75t_SL g2915 ( 
.A1(n_2903),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.C(n_178),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2901),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2902),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2899),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_2897),
.B(n_179),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2893),
.B(n_180),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2893),
.B(n_183),
.Y(n_2921)
);

OAI211xp5_ASAP7_75t_L g2922 ( 
.A1(n_2899),
.A2(n_183),
.B(n_184),
.C(n_185),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2921),
.Y(n_2923)
);

AOI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2916),
.A2(n_1498),
.B1(n_1491),
.B2(n_1485),
.Y(n_2924)
);

AOI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2919),
.A2(n_1498),
.B1(n_1491),
.B2(n_1485),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2910),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2920),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_SL g2928 ( 
.A1(n_2914),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_2928)
);

NOR2x1_ASAP7_75t_L g2929 ( 
.A(n_2912),
.B(n_188),
.Y(n_2929)
);

OAI22xp33_ASAP7_75t_L g2930 ( 
.A1(n_2909),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2907),
.Y(n_2931)
);

NOR2xp67_ASAP7_75t_L g2932 ( 
.A(n_2922),
.B(n_192),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2913),
.Y(n_2933)
);

NOR2xp33_ASAP7_75t_SL g2934 ( 
.A(n_2912),
.B(n_193),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2918),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2911),
.Y(n_2936)
);

AOI221xp5_ASAP7_75t_L g2937 ( 
.A1(n_2908),
.A2(n_194),
.B1(n_1498),
.B2(n_1491),
.C(n_1485),
.Y(n_2937)
);

AOI211xp5_ASAP7_75t_L g2938 ( 
.A1(n_2932),
.A2(n_2915),
.B(n_2917),
.C(n_2906),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_R g2939 ( 
.A(n_2934),
.B(n_195),
.Y(n_2939)
);

AND3x1_ASAP7_75t_L g2940 ( 
.A(n_2929),
.B(n_951),
.C(n_196),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2928),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2931),
.Y(n_2942)
);

AOI221xp5_ASAP7_75t_L g2943 ( 
.A1(n_2936),
.A2(n_1491),
.B1(n_1485),
.B2(n_1465),
.C(n_1461),
.Y(n_2943)
);

OAI22xp33_ASAP7_75t_L g2944 ( 
.A1(n_2923),
.A2(n_1465),
.B1(n_1461),
.B2(n_1459),
.Y(n_2944)
);

AO22x2_ASAP7_75t_L g2945 ( 
.A1(n_2935),
.A2(n_202),
.B1(n_206),
.B2(n_209),
.Y(n_2945)
);

AOI322xp5_ASAP7_75t_L g2946 ( 
.A1(n_2926),
.A2(n_214),
.A3(n_215),
.B1(n_218),
.B2(n_220),
.C1(n_224),
.C2(n_226),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2930),
.B(n_228),
.Y(n_2947)
);

AOI311xp33_ASAP7_75t_L g2948 ( 
.A1(n_2927),
.A2(n_2933),
.A3(n_2937),
.B(n_2925),
.C(n_2924),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2929),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2949),
.B(n_233),
.Y(n_2950)
);

NOR2x1_ASAP7_75t_L g2951 ( 
.A(n_2941),
.B(n_1274),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2942),
.B(n_236),
.Y(n_2952)
);

OAI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2938),
.A2(n_2947),
.B(n_2940),
.Y(n_2953)
);

XNOR2x1_ASAP7_75t_L g2954 ( 
.A(n_2945),
.B(n_237),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2939),
.Y(n_2955)
);

INVxp67_ASAP7_75t_L g2956 ( 
.A(n_2945),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2948),
.B(n_239),
.Y(n_2957)
);

AOI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2943),
.A2(n_1465),
.B1(n_1461),
.B2(n_1459),
.Y(n_2958)
);

OR2x2_ASAP7_75t_L g2959 ( 
.A(n_2944),
.B(n_240),
.Y(n_2959)
);

INVxp67_ASAP7_75t_L g2960 ( 
.A(n_2946),
.Y(n_2960)
);

NAND4xp25_ASAP7_75t_L g2961 ( 
.A(n_2953),
.B(n_1259),
.C(n_951),
.D(n_250),
.Y(n_2961)
);

A2O1A1Ixp33_ASAP7_75t_L g2962 ( 
.A1(n_2956),
.A2(n_1465),
.B(n_1461),
.C(n_1459),
.Y(n_2962)
);

OAI211xp5_ASAP7_75t_L g2963 ( 
.A1(n_2960),
.A2(n_1259),
.B(n_1452),
.C(n_1444),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2957),
.A2(n_1459),
.B1(n_1452),
.B2(n_1444),
.Y(n_2964)
);

OAI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_2954),
.A2(n_1280),
.B(n_1296),
.Y(n_2965)
);

OAI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2950),
.A2(n_1452),
.B1(n_1444),
.B2(n_951),
.Y(n_2966)
);

AOI221x1_ASAP7_75t_L g2967 ( 
.A1(n_2955),
.A2(n_2952),
.B1(n_2951),
.B2(n_2959),
.C(n_2958),
.Y(n_2967)
);

OAI22xp5_ASAP7_75t_SL g2968 ( 
.A1(n_2956),
.A2(n_1452),
.B1(n_1332),
.B2(n_1341),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2954),
.Y(n_2969)
);

OAI221xp5_ASAP7_75t_L g2970 ( 
.A1(n_2956),
.A2(n_241),
.B1(n_247),
.B2(n_257),
.C(n_258),
.Y(n_2970)
);

OAI22x1_ASAP7_75t_L g2971 ( 
.A1(n_2956),
.A2(n_259),
.B1(n_264),
.B2(n_265),
.Y(n_2971)
);

NAND5xp2_ASAP7_75t_L g2972 ( 
.A(n_2953),
.B(n_269),
.C(n_270),
.D(n_273),
.E(n_274),
.Y(n_2972)
);

OAI222xp33_ASAP7_75t_L g2973 ( 
.A1(n_2956),
.A2(n_276),
.B1(n_282),
.B2(n_285),
.C1(n_287),
.C2(n_289),
.Y(n_2973)
);

AND4x1_ASAP7_75t_L g2974 ( 
.A(n_2957),
.B(n_290),
.C(n_292),
.D(n_296),
.Y(n_2974)
);

OAI21xp33_ASAP7_75t_L g2975 ( 
.A1(n_2957),
.A2(n_1206),
.B(n_1312),
.Y(n_2975)
);

AOI211xp5_ASAP7_75t_L g2976 ( 
.A1(n_2975),
.A2(n_297),
.B(n_299),
.C(n_300),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2974),
.B(n_304),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2964),
.Y(n_2978)
);

AND3x1_ASAP7_75t_L g2979 ( 
.A(n_2969),
.B(n_305),
.C(n_307),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2965),
.B(n_309),
.Y(n_2980)
);

NOR2x1_ASAP7_75t_L g2981 ( 
.A(n_2972),
.B(n_1274),
.Y(n_2981)
);

HB1xp67_ASAP7_75t_L g2982 ( 
.A(n_2971),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2967),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2962),
.B(n_310),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2977),
.Y(n_2985)
);

HB1xp67_ASAP7_75t_L g2986 ( 
.A(n_2979),
.Y(n_2986)
);

INVx1_ASAP7_75t_SL g2987 ( 
.A(n_2982),
.Y(n_2987)
);

CKINVDCx20_ASAP7_75t_R g2988 ( 
.A(n_2983),
.Y(n_2988)
);

OAI221xp5_ASAP7_75t_L g2989 ( 
.A1(n_2981),
.A2(n_2961),
.B1(n_2963),
.B2(n_2968),
.C(n_2970),
.Y(n_2989)
);

HB1xp67_ASAP7_75t_L g2990 ( 
.A(n_2984),
.Y(n_2990)
);

NAND2x1p5_ASAP7_75t_L g2991 ( 
.A(n_2978),
.B(n_2973),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2980),
.Y(n_2992)
);

CKINVDCx5p33_ASAP7_75t_R g2993 ( 
.A(n_2976),
.Y(n_2993)
);

CKINVDCx20_ASAP7_75t_R g2994 ( 
.A(n_2982),
.Y(n_2994)
);

OAI21xp33_ASAP7_75t_SL g2995 ( 
.A1(n_2983),
.A2(n_2966),
.B(n_1341),
.Y(n_2995)
);

INVxp67_ASAP7_75t_L g2996 ( 
.A(n_2979),
.Y(n_2996)
);

BUFx2_ASAP7_75t_L g2997 ( 
.A(n_2979),
.Y(n_2997)
);

HB1xp67_ASAP7_75t_L g2998 ( 
.A(n_2979),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2977),
.Y(n_2999)
);

OR2x6_ASAP7_75t_L g3000 ( 
.A(n_2983),
.B(n_313),
.Y(n_3000)
);

INVx3_ASAP7_75t_SL g3001 ( 
.A(n_2983),
.Y(n_3001)
);

CKINVDCx5p33_ASAP7_75t_R g3002 ( 
.A(n_2983),
.Y(n_3002)
);

INVxp67_ASAP7_75t_SL g3003 ( 
.A(n_2977),
.Y(n_3003)
);

NAND3xp33_ASAP7_75t_L g3004 ( 
.A(n_2983),
.B(n_1319),
.C(n_907),
.Y(n_3004)
);

AOI211x1_ASAP7_75t_L g3005 ( 
.A1(n_2983),
.A2(n_315),
.B(n_324),
.C(n_327),
.Y(n_3005)
);

OR2x2_ASAP7_75t_L g3006 ( 
.A(n_2977),
.B(n_332),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2977),
.Y(n_3007)
);

OAI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2987),
.A2(n_1211),
.B(n_1219),
.Y(n_3008)
);

OAI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2996),
.A2(n_1211),
.B(n_1219),
.Y(n_3009)
);

AOI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_2994),
.A2(n_2988),
.B1(n_3002),
.B2(n_3001),
.Y(n_3010)
);

INVxp67_ASAP7_75t_L g3011 ( 
.A(n_3000),
.Y(n_3011)
);

HB1xp67_ASAP7_75t_L g3012 ( 
.A(n_3000),
.Y(n_3012)
);

AO21x2_ASAP7_75t_L g3013 ( 
.A1(n_2985),
.A2(n_334),
.B(n_337),
.Y(n_3013)
);

HB1xp67_ASAP7_75t_L g3014 ( 
.A(n_2986),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_3006),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2997),
.B(n_340),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2998),
.Y(n_3017)
);

INVxp67_ASAP7_75t_L g3018 ( 
.A(n_2990),
.Y(n_3018)
);

INVxp67_ASAP7_75t_L g3019 ( 
.A(n_2991),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_3003),
.Y(n_3020)
);

OAI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2989),
.A2(n_1332),
.B1(n_1341),
.B2(n_1323),
.Y(n_3021)
);

OA22x2_ASAP7_75t_L g3022 ( 
.A1(n_2993),
.A2(n_3007),
.B1(n_2999),
.B2(n_2992),
.Y(n_3022)
);

AO22x2_ASAP7_75t_L g3023 ( 
.A1(n_3004),
.A2(n_344),
.B1(n_348),
.B2(n_352),
.Y(n_3023)
);

AND2x4_ASAP7_75t_L g3024 ( 
.A(n_3005),
.B(n_354),
.Y(n_3024)
);

HB1xp67_ASAP7_75t_L g3025 ( 
.A(n_2995),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_3000),
.Y(n_3026)
);

AOI31xp33_ASAP7_75t_L g3027 ( 
.A1(n_2991),
.A2(n_356),
.A3(n_357),
.B(n_361),
.Y(n_3027)
);

INVxp67_ASAP7_75t_L g3028 ( 
.A(n_3000),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_3001),
.B(n_362),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_3006),
.Y(n_3030)
);

XOR2xp5_ASAP7_75t_L g3031 ( 
.A(n_2994),
.B(n_363),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_3000),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_3006),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_3006),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_3001),
.B(n_365),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_2994),
.A2(n_1332),
.B1(n_877),
.B2(n_1329),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_3006),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_3006),
.Y(n_3038)
);

AOI221x1_ASAP7_75t_SL g3039 ( 
.A1(n_2985),
.A2(n_368),
.B1(n_371),
.B2(n_373),
.C(n_375),
.Y(n_3039)
);

NOR4xp75_ASAP7_75t_L g3040 ( 
.A(n_3029),
.B(n_377),
.C(n_382),
.D(n_388),
.Y(n_3040)
);

OAI222xp33_ASAP7_75t_L g3041 ( 
.A1(n_3010),
.A2(n_389),
.B1(n_391),
.B2(n_393),
.C1(n_394),
.C2(n_397),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_3019),
.A2(n_1296),
.B1(n_1219),
.B2(n_1280),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_3016),
.Y(n_3043)
);

OAI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_3018),
.A2(n_877),
.B1(n_1329),
.B2(n_1328),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_3013),
.Y(n_3045)
);

XOR2xp5_ASAP7_75t_L g3046 ( 
.A(n_3014),
.B(n_398),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_3017),
.A2(n_895),
.B(n_904),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_3035),
.Y(n_3048)
);

NAND4xp25_ASAP7_75t_L g3049 ( 
.A(n_3020),
.B(n_399),
.C(n_400),
.D(n_402),
.Y(n_3049)
);

AND3x1_ASAP7_75t_L g3050 ( 
.A(n_3032),
.B(n_414),
.C(n_415),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_3012),
.Y(n_3051)
);

NAND3xp33_ASAP7_75t_L g3052 ( 
.A(n_3011),
.B(n_904),
.C(n_918),
.Y(n_3052)
);

NAND4xp25_ASAP7_75t_L g3053 ( 
.A(n_3026),
.B(n_416),
.C(n_417),
.D(n_419),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_3028),
.A2(n_3024),
.B1(n_3038),
.B2(n_3037),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3023),
.Y(n_3055)
);

NOR3xp33_ASAP7_75t_L g3056 ( 
.A(n_3030),
.B(n_3033),
.C(n_3034),
.Y(n_3056)
);

XNOR2xp5_ASAP7_75t_L g3057 ( 
.A(n_3031),
.B(n_1331),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_3024),
.B(n_883),
.Y(n_3058)
);

INVx2_ASAP7_75t_SL g3059 ( 
.A(n_3015),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_3027),
.B(n_877),
.Y(n_3060)
);

XNOR2xp5_ASAP7_75t_L g3061 ( 
.A(n_3022),
.B(n_1331),
.Y(n_3061)
);

OAI222xp33_ASAP7_75t_L g3062 ( 
.A1(n_3025),
.A2(n_1298),
.B1(n_1323),
.B2(n_1328),
.C1(n_1326),
.C2(n_1322),
.Y(n_3062)
);

OAI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_3023),
.A2(n_877),
.B1(n_1326),
.B2(n_1315),
.Y(n_3063)
);

AND2x2_ASAP7_75t_SL g3064 ( 
.A(n_3039),
.B(n_895),
.Y(n_3064)
);

OA22x2_ASAP7_75t_L g3065 ( 
.A1(n_3036),
.A2(n_1322),
.B1(n_1315),
.B2(n_1323),
.Y(n_3065)
);

AOI22xp5_ASAP7_75t_L g3066 ( 
.A1(n_3051),
.A2(n_3021),
.B1(n_3008),
.B2(n_3009),
.Y(n_3066)
);

OAI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_3059),
.A2(n_1296),
.B(n_883),
.Y(n_3067)
);

AOI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_3056),
.A2(n_1296),
.B1(n_1280),
.B2(n_883),
.Y(n_3068)
);

INVx2_ASAP7_75t_SL g3069 ( 
.A(n_3045),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3057),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_3058),
.A2(n_895),
.B(n_906),
.Y(n_3071)
);

AND3x2_ASAP7_75t_L g3072 ( 
.A(n_3060),
.B(n_883),
.C(n_956),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3064),
.Y(n_3073)
);

OAI22xp33_ASAP7_75t_SL g3074 ( 
.A1(n_3043),
.A2(n_1298),
.B1(n_1206),
.B2(n_1114),
.Y(n_3074)
);

OAI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_3054),
.A2(n_1206),
.B1(n_907),
.B2(n_901),
.Y(n_3075)
);

AOI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_3050),
.A2(n_1280),
.B1(n_883),
.B2(n_956),
.Y(n_3076)
);

OA21x2_ASAP7_75t_L g3077 ( 
.A1(n_3055),
.A2(n_956),
.B(n_901),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_3046),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_3048),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_3061),
.A2(n_956),
.B1(n_901),
.B2(n_904),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3040),
.Y(n_3081)
);

AOI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_3063),
.A2(n_956),
.B1(n_901),
.B2(n_904),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3065),
.Y(n_3083)
);

INVxp67_ASAP7_75t_L g3084 ( 
.A(n_3069),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_3072),
.Y(n_3085)
);

NOR3xp33_ASAP7_75t_L g3086 ( 
.A(n_3079),
.B(n_3052),
.C(n_3047),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3081),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_3078),
.Y(n_3088)
);

XOR2xp5_ASAP7_75t_L g3089 ( 
.A(n_3070),
.B(n_3053),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_3073),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3083),
.Y(n_3091)
);

CKINVDCx20_ASAP7_75t_R g3092 ( 
.A(n_3066),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_3071),
.A2(n_3044),
.B(n_3062),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3076),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_3080),
.B(n_3049),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_3077),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_3082),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3074),
.Y(n_3098)
);

INVx1_ASAP7_75t_SL g3099 ( 
.A(n_3075),
.Y(n_3099)
);

AOI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_3084),
.A2(n_3041),
.B1(n_3067),
.B2(n_3068),
.Y(n_3100)
);

XNOR2xp5_ASAP7_75t_L g3101 ( 
.A(n_3089),
.B(n_3042),
.Y(n_3101)
);

OAI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_3092),
.A2(n_904),
.B1(n_906),
.B2(n_907),
.Y(n_3102)
);

OAI222xp33_ASAP7_75t_L g3103 ( 
.A1(n_3091),
.A2(n_1133),
.B1(n_1114),
.B2(n_1166),
.C1(n_1162),
.C2(n_893),
.Y(n_3103)
);

OAI21xp33_ASAP7_75t_L g3104 ( 
.A1(n_3087),
.A2(n_1133),
.B(n_906),
.Y(n_3104)
);

AOI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_3088),
.A2(n_956),
.B1(n_906),
.B2(n_907),
.Y(n_3105)
);

AOI221xp5_ASAP7_75t_L g3106 ( 
.A1(n_3090),
.A2(n_906),
.B1(n_907),
.B2(n_918),
.C(n_911),
.Y(n_3106)
);

OAI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_3095),
.A2(n_1133),
.B(n_910),
.Y(n_3107)
);

AOI221xp5_ASAP7_75t_L g3108 ( 
.A1(n_3086),
.A2(n_918),
.B1(n_911),
.B2(n_1134),
.C(n_1041),
.Y(n_3108)
);

OA21x2_ASAP7_75t_L g3109 ( 
.A1(n_3096),
.A2(n_918),
.B(n_911),
.Y(n_3109)
);

OAI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_3100),
.A2(n_3101),
.B(n_3094),
.Y(n_3110)
);

OAI321xp33_ASAP7_75t_L g3111 ( 
.A1(n_3104),
.A2(n_3085),
.A3(n_3098),
.B1(n_3097),
.B2(n_3093),
.C(n_3099),
.Y(n_3111)
);

NOR2xp67_ASAP7_75t_L g3112 ( 
.A(n_3107),
.B(n_911),
.Y(n_3112)
);

INVx4_ASAP7_75t_L g3113 ( 
.A(n_3109),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3102),
.Y(n_3114)
);

XOR2xp5_ASAP7_75t_L g3115 ( 
.A(n_3109),
.B(n_918),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_3111),
.B(n_3103),
.Y(n_3116)
);

AOI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_3116),
.A2(n_3110),
.B1(n_3114),
.B2(n_3112),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3117),
.Y(n_3118)
);

AO22x2_ASAP7_75t_L g3119 ( 
.A1(n_3118),
.A2(n_3113),
.B1(n_3115),
.B2(n_3106),
.Y(n_3119)
);

AOI211xp5_ASAP7_75t_L g3120 ( 
.A1(n_3119),
.A2(n_3108),
.B(n_3105),
.C(n_911),
.Y(n_3120)
);


endmodule