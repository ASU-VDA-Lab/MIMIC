module fake_jpeg_14244_n_559 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_559);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_559;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_58),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_30),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_51),
.B1(n_20),
.B2(n_25),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_11),
.Y(n_93)
);

NAND2x1_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_51),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_33),
.B(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_99),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_101),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_104),
.Y(n_160)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_37),
.Y(n_109)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_109),
.B(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_24),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_120),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_64),
.B(n_42),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_61),
.A2(n_35),
.B1(n_51),
.B2(n_29),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_150),
.B1(n_148),
.B2(n_129),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_24),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_26),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_101),
.A2(n_35),
.B1(n_19),
.B2(n_50),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_35),
.B1(n_27),
.B2(n_46),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g222 ( 
.A1(n_156),
.A2(n_27),
.B1(n_59),
.B2(n_50),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_64),
.B(n_46),
.Y(n_159)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_126),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_171),
.B(n_176),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_101),
.B1(n_88),
.B2(n_85),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_172),
.A2(n_184),
.B1(n_189),
.B2(n_207),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_60),
.B(n_29),
.C(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_182),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_94),
.B1(n_66),
.B2(n_67),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_177),
.Y(n_275)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_31),
.B(n_29),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_179),
.A2(n_136),
.B(n_50),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_114),
.Y(n_182)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_112),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_187),
.B(n_190),
.Y(n_262)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_102),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_122),
.B(n_42),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_201),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_20),
.C(n_31),
.Y(n_197)
);

AOI32xp33_ASAP7_75t_L g257 ( 
.A1(n_197),
.A2(n_11),
.A3(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_257)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_200),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_141),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_223),
.B1(n_227),
.B2(n_142),
.Y(n_238)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_156),
.A2(n_55),
.B1(n_69),
.B2(n_62),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_150),
.A2(n_113),
.B1(n_128),
.B2(n_145),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_208),
.A2(n_222),
.B1(n_225),
.B2(n_0),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_39),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_191),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_117),
.A2(n_97),
.B1(n_58),
.B2(n_76),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_216),
.B1(n_219),
.B2(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_130),
.B(n_39),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_164),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_125),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_147),
.B(n_26),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_162),
.A2(n_28),
.B1(n_19),
.B2(n_50),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_116),
.A2(n_102),
.B1(n_99),
.B2(n_82),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_105),
.A2(n_116),
.B1(n_127),
.B2(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_125),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_228),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_105),
.A2(n_99),
.B1(n_82),
.B2(n_50),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_232),
.A2(n_278),
.B(n_15),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_238),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_169),
.A2(n_136),
.B1(n_119),
.B2(n_158),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_246),
.B1(n_247),
.B2(n_251),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_244),
.A2(n_194),
.B1(n_8),
.B2(n_9),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_171),
.A2(n_158),
.B1(n_161),
.B2(n_110),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_182),
.A2(n_161),
.B1(n_110),
.B2(n_131),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_203),
.B1(n_207),
.B2(n_173),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_200),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_255),
.B(n_268),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_257),
.B(n_258),
.Y(n_330)
);

AOI32xp33_ASAP7_75t_L g258 ( 
.A1(n_191),
.A2(n_10),
.A3(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_189),
.A2(n_213),
.B1(n_210),
.B2(n_206),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_264),
.B1(n_265),
.B2(n_273),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_12),
.B1(n_2),
.B2(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_12),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_177),
.B(n_13),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_214),
.A2(n_10),
.B1(n_4),
.B2(n_7),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_209),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_277),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_211),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_280),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_214),
.A2(n_0),
.B1(n_7),
.B2(n_8),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_239),
.B1(n_246),
.B2(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_242),
.A2(n_179),
.B(n_205),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_284),
.A2(n_298),
.B(n_308),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_197),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_307),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_288),
.A2(n_297),
.B1(n_304),
.B2(n_305),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_198),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_299),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_225),
.B1(n_214),
.B2(n_229),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_205),
.B(n_227),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_199),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_233),
.B(n_170),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_302),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_235),
.A2(n_223),
.B1(n_221),
.B2(n_220),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_309),
.B1(n_313),
.B2(n_326),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_192),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_193),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_319),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_235),
.A2(n_188),
.B1(n_224),
.B2(n_228),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_238),
.A2(n_224),
.B1(n_204),
.B2(n_175),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_185),
.C(n_226),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_183),
.C(n_168),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_241),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_264),
.A2(n_195),
.B1(n_178),
.B2(n_212),
.Y(n_309)
);

BUFx12_ASAP7_75t_L g310 ( 
.A(n_236),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_312),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_280),
.A2(n_15),
.B1(n_8),
.B2(n_9),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_318),
.B1(n_237),
.B2(n_245),
.Y(n_359)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_236),
.A2(n_241),
.B(n_248),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_316),
.A2(n_323),
.B(n_237),
.Y(n_361)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_322),
.Y(n_333)
);

AO21x2_ASAP7_75t_L g318 ( 
.A1(n_236),
.A2(n_0),
.B(n_14),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_15),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_15),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_324),
.Y(n_365)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_230),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_260),
.B(n_267),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_327),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_258),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_236),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_328),
.Y(n_340)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_230),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_329),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_240),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_320),
.A2(n_257),
.B1(n_276),
.B2(n_272),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_350),
.B1(n_358),
.B2(n_313),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_341),
.A2(n_352),
.B(n_318),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_294),
.B(n_260),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_343),
.B(n_344),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_285),
.B(n_263),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_300),
.B(n_267),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_359),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_331),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_286),
.A2(n_276),
.B1(n_275),
.B2(n_269),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_303),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_353),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_284),
.A2(n_269),
.B(n_266),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_324),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_298),
.B(n_290),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_355),
.A2(n_363),
.B(n_366),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_252),
.B1(n_231),
.B2(n_275),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_356),
.A2(n_372),
.B1(n_305),
.B2(n_297),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_286),
.A2(n_231),
.B1(n_271),
.B2(n_237),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_316),
.A2(n_266),
.B(n_261),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_292),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_322),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_299),
.B(n_254),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_261),
.Y(n_367)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_367),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_271),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_368),
.B(n_374),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_271),
.B(n_279),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g398 ( 
.A1(n_370),
.A2(n_318),
.B(n_314),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_307),
.B(n_302),
.C(n_319),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_316),
.C(n_289),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_309),
.A2(n_240),
.B1(n_234),
.B2(n_279),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_283),
.B(n_234),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_378),
.C(n_380),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_377),
.A2(n_349),
.B1(n_350),
.B2(n_358),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_317),
.C(n_288),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_379),
.A2(n_398),
.B1(n_347),
.B2(n_351),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_304),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_293),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_392),
.C(n_394),
.Y(n_416)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_342),
.Y(n_428)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_389),
.Y(n_425)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_334),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_390),
.B(n_406),
.Y(n_417)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_402),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_329),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_341),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_354),
.B(n_312),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_403),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_310),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_397),
.C(n_405),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_332),
.B(n_310),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_401),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_327),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_332),
.B(n_245),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_340),
.B(n_245),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_409),
.Y(n_438)
);

OAI32xp33_ASAP7_75t_L g409 ( 
.A1(n_343),
.A2(n_325),
.A3(n_306),
.B1(n_318),
.B2(n_17),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_335),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_318),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_411),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_388),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_427),
.B1(n_441),
.B2(n_383),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_418),
.A2(n_432),
.B1(n_427),
.B2(n_421),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_376),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_419),
.B(n_424),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_434),
.B1(n_435),
.B2(n_440),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_408),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_371),
.C(n_353),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_393),
.C(n_397),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_408),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_430),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_342),
.Y(n_430)
);

XOR2x2_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_370),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_396),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_349),
.B1(n_339),
.B2(n_359),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_404),
.A2(n_361),
.B1(n_365),
.B2(n_340),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_433),
.A2(n_411),
.B(n_399),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_379),
.A2(n_347),
.B1(n_356),
.B2(n_366),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_366),
.B1(n_365),
.B2(n_372),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_392),
.B(n_354),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_443),
.Y(n_454)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_439),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_404),
.A2(n_367),
.B1(n_346),
.B2(n_335),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_401),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_375),
.B(n_373),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_373),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_393),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_445),
.B(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_447),
.B(n_455),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_378),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_458),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_450),
.A2(n_435),
.B1(n_434),
.B2(n_440),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_383),
.Y(n_451)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_451),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_409),
.Y(n_453)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_437),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_391),
.Y(n_459)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_461),
.A2(n_469),
.B(n_429),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_405),
.Y(n_462)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_422),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_470),
.Y(n_483)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

XNOR2x2_ASAP7_75t_SL g467 ( 
.A(n_433),
.B(n_399),
.Y(n_467)
);

NOR3xp33_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_438),
.C(n_431),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_400),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_471),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_429),
.A2(n_411),
.B(n_336),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_417),
.Y(n_470)
);

XNOR2x1_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_377),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_416),
.B(n_369),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_444),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_473),
.A2(n_462),
.B1(n_426),
.B2(n_467),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_486),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_461),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_478),
.B(n_479),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_448),
.B(n_412),
.C(n_443),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_423),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_489),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_430),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_492),
.B(n_493),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_428),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_336),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_495),
.B(n_459),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_483),
.A2(n_465),
.B1(n_457),
.B2(n_453),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_501),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_497),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_450),
.B1(n_485),
.B2(n_487),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_499),
.A2(n_505),
.B1(n_509),
.B2(n_481),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_457),
.B1(n_432),
.B2(n_418),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_512),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_490),
.A2(n_414),
.B1(n_463),
.B2(n_421),
.Y(n_505)
);

XNOR2x1_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_445),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_507),
.A2(n_474),
.B1(n_449),
.B2(n_454),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_479),
.B(n_458),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_475),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_490),
.A2(n_460),
.B1(n_472),
.B2(n_471),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_510),
.B(n_491),
.Y(n_516)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_481),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_513),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_454),
.C(n_449),
.Y(n_513)
);

OAI321xp33_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_491),
.A3(n_484),
.B1(n_494),
.B2(n_489),
.C(n_476),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_514),
.B(n_515),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_523),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_504),
.C(n_505),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_522),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_502),
.B(n_486),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_474),
.C(n_480),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_504),
.C(n_509),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_524),
.A2(n_498),
.B(n_338),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_480),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_525),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_527),
.Y(n_532)
);

NOR2x1_ASAP7_75t_SL g527 ( 
.A(n_506),
.B(n_436),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_531),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_499),
.C(n_511),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_533),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_524),
.A2(n_402),
.B(n_338),
.Y(n_535)
);

AOI21xp33_ASAP7_75t_L g541 ( 
.A1(n_535),
.A2(n_519),
.B(n_521),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_360),
.C(n_402),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_539),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_362),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_526),
.B(n_520),
.Y(n_540)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_540),
.Y(n_547)
);

NOR2x1_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_536),
.Y(n_549)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_534),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_545),
.C(n_536),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_538),
.A2(n_523),
.B1(n_525),
.B2(n_517),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_544),
.A2(n_532),
.B(n_530),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_548),
.A2(n_549),
.B(n_550),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_546),
.C(n_543),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_552),
.B(n_553),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_549),
.A2(n_530),
.B(n_540),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_551),
.A2(n_369),
.B(n_362),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_360),
.C(n_16),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_554),
.C(n_18),
.Y(n_557)
);

NAND3xp33_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_18),
.C(n_236),
.Y(n_558)
);

BUFx24_ASAP7_75t_SL g559 ( 
.A(n_558),
.Y(n_559)
);


endmodule