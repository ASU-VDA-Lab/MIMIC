module real_aes_10474_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_1893, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_1893;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_1883;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_1856;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1802;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_727;
wire n_1855;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1584;
wire n_466;
wire n_1277;
wire n_1049;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVxp67_ASAP7_75t_SL g1810 ( .A(n_0), .Y(n_1810) );
AOI22xp33_ASAP7_75t_L g1828 ( .A1(n_0), .A2(n_8), .B1(n_902), .B2(n_1829), .Y(n_1828) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_1), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_2), .A2(n_312), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g657 ( .A(n_2), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g1823 ( .A1(n_3), .A2(n_239), .B1(n_450), .B2(n_1017), .Y(n_1823) );
AOI22xp33_ASAP7_75t_L g1834 ( .A1(n_3), .A2(n_239), .B1(n_481), .B2(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1804 ( .A(n_4), .Y(n_1804) );
INVx1_ASAP7_75t_L g1248 ( .A(n_5), .Y(n_1248) );
CKINVDCx5p33_ASAP7_75t_R g1407 ( .A(n_6), .Y(n_1407) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_7), .Y(n_1426) );
INVx1_ASAP7_75t_L g1809 ( .A(n_8), .Y(n_1809) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_9), .A2(n_103), .B1(n_752), .B2(n_755), .Y(n_1446) );
INVx1_ASAP7_75t_L g1484 ( .A(n_9), .Y(n_1484) );
INVx1_ASAP7_75t_L g1508 ( .A(n_10), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g1534 ( .A1(n_10), .A2(n_149), .B1(n_1535), .B2(n_1536), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_11), .A2(n_210), .B1(n_432), .B2(n_436), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_11), .A2(n_210), .B1(n_472), .B2(n_474), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_12), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_13), .A2(n_200), .B1(n_633), .B2(n_711), .C(n_1065), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g1187 ( .A1(n_13), .A2(n_310), .B1(n_543), .B2(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1595 ( .A(n_14), .Y(n_1595) );
INVx1_ASAP7_75t_L g1059 ( .A(n_15), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_15), .A2(n_112), .B1(n_582), .B2(n_1076), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_16), .A2(n_35), .B1(n_1310), .B2(n_1311), .C(n_1313), .Y(n_1309) );
INVx1_ASAP7_75t_L g1372 ( .A(n_16), .Y(n_1372) );
OAI22xp33_ASAP7_75t_L g1873 ( .A1(n_17), .A2(n_102), .B1(n_613), .B2(n_642), .Y(n_1873) );
AOI221xp5_ASAP7_75t_L g1879 ( .A1(n_17), .A2(n_102), .B1(n_587), .B2(n_696), .C(n_1880), .Y(n_1879) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_18), .A2(n_270), .B1(n_769), .B2(n_1019), .C(n_1024), .Y(n_1228) );
OAI22xp33_ASAP7_75t_L g1234 ( .A1(n_18), .A2(n_110), .B1(n_866), .B2(n_869), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_19), .A2(n_121), .B1(n_704), .B2(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g1073 ( .A1(n_19), .A2(n_121), .B1(n_987), .B2(n_1006), .Y(n_1073) );
INVx1_ASAP7_75t_L g818 ( .A(n_20), .Y(n_818) );
OAI211xp5_ASAP7_75t_SL g848 ( .A1(n_20), .A2(n_613), .B(n_849), .C(n_859), .Y(n_848) );
INVx1_ASAP7_75t_L g1803 ( .A(n_21), .Y(n_1803) );
AOI22xp33_ASAP7_75t_L g1830 ( .A1(n_21), .A2(n_64), .B1(n_630), .B2(n_1019), .Y(n_1830) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_22), .Y(n_810) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_23), .A2(n_73), .B1(n_752), .B2(n_755), .Y(n_751) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_23), .A2(n_187), .B1(n_358), .B2(n_521), .Y(n_762) );
AO22x2_ASAP7_75t_L g370 ( .A1(n_24), .A2(n_371), .B1(n_523), .B2(n_524), .Y(n_370) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_24), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g1518 ( .A1(n_25), .A2(n_433), .B(n_1024), .Y(n_1518) );
INVx1_ASAP7_75t_L g1522 ( .A(n_25), .Y(n_1522) );
AOI22xp5_ASAP7_75t_L g1620 ( .A1(n_26), .A2(n_131), .B1(n_1581), .B2(n_1584), .Y(n_1620) );
AOI22xp33_ASAP7_75t_SL g1068 ( .A1(n_27), .A2(n_95), .B1(n_704), .B2(n_1069), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_27), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_28), .A2(n_341), .B1(n_486), .B2(n_787), .Y(n_1152) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_28), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_29), .A2(n_139), .B1(n_1296), .B2(n_1297), .Y(n_1295) );
INVx1_ASAP7_75t_L g1340 ( .A(n_29), .Y(n_1340) );
INVx1_ASAP7_75t_L g746 ( .A(n_30), .Y(n_746) );
OAI222xp33_ASAP7_75t_L g759 ( .A1(n_30), .A2(n_233), .B1(n_321), .B2(n_505), .C1(n_760), .C2(n_761), .Y(n_759) );
OAI222xp33_ASAP7_75t_L g939 ( .A1(n_31), .A2(n_71), .B1(n_151), .B2(n_684), .C1(n_940), .C2(n_943), .Y(n_939) );
INVx1_ASAP7_75t_L g960 ( .A(n_31), .Y(n_960) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_32), .Y(n_1029) );
CKINVDCx5p33_ASAP7_75t_R g1301 ( .A(n_33), .Y(n_1301) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_34), .A2(n_138), .B1(n_577), .B2(n_590), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_34), .A2(n_138), .B1(n_715), .B2(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g1368 ( .A(n_35), .Y(n_1368) );
INVx1_ASAP7_75t_L g680 ( .A(n_36), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_36), .A2(n_324), .B1(n_438), .B2(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g1390 ( .A(n_37), .Y(n_1390) );
AOI221xp5_ASAP7_75t_L g1415 ( .A1(n_37), .A2(n_161), .B1(n_1292), .B2(n_1293), .C(n_1416), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1445 ( .A(n_38), .B(n_750), .Y(n_1445) );
INVx1_ASAP7_75t_L g1482 ( .A(n_38), .Y(n_1482) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_39), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_40), .A2(n_160), .B1(n_591), .B2(n_724), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_40), .A2(n_160), .B1(n_450), .B2(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_41), .A2(n_259), .B1(n_443), .B2(n_448), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_41), .A2(n_259), .B1(n_478), .B2(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g349 ( .A(n_42), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g1615 ( .A1(n_43), .A2(n_124), .B1(n_1581), .B2(n_1584), .Y(n_1615) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_44), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_45), .A2(n_120), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_45), .A2(n_120), .B1(n_706), .B2(n_715), .Y(n_773) );
INVx1_ASAP7_75t_L g1251 ( .A(n_46), .Y(n_1251) );
OAI211xp5_ASAP7_75t_SL g1272 ( .A1(n_46), .A2(n_613), .B(n_1273), .C(n_1278), .Y(n_1272) );
AOI21xp33_ASAP7_75t_L g1505 ( .A1(n_47), .A2(n_769), .B(n_1020), .Y(n_1505) );
INVx1_ASAP7_75t_L g1532 ( .A(n_47), .Y(n_1532) );
INVx1_ASAP7_75t_L g1562 ( .A(n_48), .Y(n_1562) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_49), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_49), .A2(n_182), .B1(n_684), .B2(n_940), .Y(n_1084) );
INVx1_ASAP7_75t_L g1097 ( .A(n_50), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_50), .A2(n_219), .B1(n_711), .B2(n_770), .Y(n_1126) );
INVx1_ASAP7_75t_L g764 ( .A(n_51), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_51), .A2(n_232), .B1(n_486), .B2(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_52), .A2(n_152), .B1(n_630), .B2(n_770), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_52), .A2(n_152), .B1(n_694), .B2(n_696), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_53), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_54), .A2(n_247), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g649 ( .A(n_54), .Y(n_649) );
INVx1_ASAP7_75t_L g1397 ( .A(n_55), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_55), .A2(n_136), .B1(n_483), .B2(n_1079), .Y(n_1424) );
AOI22x1_ASAP7_75t_SL g737 ( .A1(n_56), .A2(n_738), .B1(n_788), .B2(n_789), .Y(n_737) );
INVx1_ASAP7_75t_L g788 ( .A(n_56), .Y(n_788) );
INVx1_ASAP7_75t_L g1284 ( .A(n_57), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1621 ( .A1(n_57), .A2(n_75), .B1(n_1552), .B2(n_1560), .Y(n_1621) );
XNOR2xp5_ASAP7_75t_L g792 ( .A(n_58), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g1206 ( .A(n_59), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1214 ( .A1(n_59), .A2(n_642), .B1(n_847), .B2(n_1215), .C(n_1219), .Y(n_1214) );
INVx1_ASAP7_75t_L g887 ( .A(n_60), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_60), .A2(n_613), .B1(n_908), .B2(n_916), .C(n_922), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g1258 ( .A1(n_61), .A2(n_245), .B1(n_536), .B2(n_543), .Y(n_1258) );
INVx1_ASAP7_75t_L g1276 ( .A(n_61), .Y(n_1276) );
INVx1_ASAP7_75t_L g1148 ( .A(n_62), .Y(n_1148) );
INVx1_ASAP7_75t_L g689 ( .A(n_63), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_63), .A2(n_185), .B1(n_704), .B2(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g1806 ( .A(n_64), .Y(n_1806) );
INVx1_ASAP7_75t_L g1813 ( .A(n_65), .Y(n_1813) );
AOI22xp33_ASAP7_75t_L g1837 ( .A1(n_65), .A2(n_264), .B1(n_582), .B2(n_596), .Y(n_1837) );
INVx1_ASAP7_75t_L g967 ( .A(n_66), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g984 ( .A1(n_66), .A2(n_119), .B1(n_696), .B2(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1858 ( .A(n_67), .Y(n_1858) );
AOI221xp5_ASAP7_75t_L g1875 ( .A1(n_67), .A2(n_255), .B1(n_696), .B2(n_1876), .C(n_1878), .Y(n_1875) );
AOI22xp33_ASAP7_75t_L g1599 ( .A1(n_68), .A2(n_209), .B1(n_1581), .B2(n_1584), .Y(n_1599) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_69), .Y(n_807) );
AO22x1_ASAP7_75t_SL g1608 ( .A1(n_70), .A2(n_133), .B1(n_1581), .B2(n_1584), .Y(n_1608) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_71), .A2(n_303), .B1(n_630), .B2(n_718), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_72), .A2(n_197), .B1(n_704), .B2(n_920), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_72), .A2(n_197), .B1(n_480), .B2(n_987), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_73), .A2(n_147), .B1(n_432), .B2(n_770), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_74), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_76), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_77), .A2(n_155), .B1(n_769), .B2(n_770), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_77), .A2(n_155), .B1(n_483), .B2(n_782), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_78), .Y(n_1320) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_79), .A2(n_336), .B1(n_828), .B2(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g861 ( .A(n_79), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g1600 ( .A1(n_80), .A2(n_229), .B1(n_1560), .B2(n_1587), .Y(n_1600) );
INVx1_ASAP7_75t_L g911 ( .A(n_81), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_81), .A2(n_175), .B1(n_536), .B2(n_543), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_82), .A2(n_250), .B1(n_1303), .B2(n_1306), .Y(n_1302) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_82), .A2(n_250), .B1(n_1352), .B2(n_1356), .C(n_1359), .Y(n_1351) );
INVx1_ASAP7_75t_L g1255 ( .A(n_83), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_83), .A2(n_231), .B1(n_835), .B2(n_836), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_84), .A2(n_337), .B1(n_583), .B2(n_587), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_84), .A2(n_642), .B1(n_644), .B2(n_656), .C(n_661), .Y(n_641) );
INVx1_ASAP7_75t_L g1098 ( .A(n_85), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_85), .A2(n_173), .B1(n_704), .B2(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1389 ( .A(n_86), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_86), .A2(n_226), .B1(n_478), .B2(n_1418), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_87), .A2(n_257), .B1(n_480), .B2(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g512 ( .A(n_87), .Y(n_512) );
XOR2xp5_ASAP7_75t_L g1849 ( .A(n_88), .B(n_1850), .Y(n_1849) );
INVx1_ASAP7_75t_L g402 ( .A(n_89), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_89), .A2(n_196), .B1(n_502), .B2(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g825 ( .A(n_90), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_90), .A2(n_294), .B1(n_835), .B2(n_836), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g1141 ( .A(n_91), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g1586 ( .A1(n_92), .A2(n_118), .B1(n_1560), .B2(n_1587), .Y(n_1586) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_93), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_93), .A2(n_261), .B1(n_987), .B2(n_1079), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1394 ( .A1(n_94), .A2(n_123), .B1(n_1352), .B2(n_1356), .C(n_1359), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_94), .A2(n_123), .B1(n_1303), .B2(n_1306), .Y(n_1420) );
INVxp33_ASAP7_75t_L g1089 ( .A(n_95), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g1867 ( .A(n_96), .Y(n_1867) );
BUFx2_ASAP7_75t_L g424 ( .A(n_97), .Y(n_424) );
INVx1_ASAP7_75t_L g461 ( .A(n_97), .Y(n_461) );
BUFx2_ASAP7_75t_L g489 ( .A(n_97), .Y(n_489) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_97), .B(n_609), .Y(n_1335) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_98), .A2(n_241), .B1(n_443), .B2(n_706), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_98), .A2(n_241), .B1(n_777), .B2(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g1499 ( .A(n_99), .Y(n_1499) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_99), .A2(n_141), .B1(n_487), .B2(n_779), .Y(n_1538) );
INVx1_ASAP7_75t_L g1569 ( .A(n_100), .Y(n_1569) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_101), .A2(n_332), .B1(n_694), .B2(n_696), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_101), .A2(n_332), .B1(n_711), .B2(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g1441 ( .A(n_103), .Y(n_1441) );
INVx1_ASAP7_75t_L g917 ( .A(n_104), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_104), .A2(n_198), .B1(n_866), .B2(n_869), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_105), .A2(n_162), .B1(n_683), .B2(n_684), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_105), .A2(n_162), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g1603 ( .A1(n_106), .A2(n_302), .B1(n_1581), .B2(n_1584), .Y(n_1603) );
CKINVDCx5p33_ASAP7_75t_R g1856 ( .A(n_107), .Y(n_1856) );
INVx1_ASAP7_75t_L g549 ( .A(n_108), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_108), .A2(n_290), .B1(n_629), .B2(n_630), .C(n_633), .Y(n_628) );
INVx1_ASAP7_75t_L g890 ( .A(n_109), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_109), .A2(n_113), .B1(n_835), .B2(n_836), .Y(n_895) );
INVx1_ASAP7_75t_L g1226 ( .A(n_110), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_111), .A2(n_205), .B1(n_711), .B2(n_1071), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_111), .Y(n_1082) );
INVxp33_ASAP7_75t_L g1055 ( .A(n_112), .Y(n_1055) );
INVx1_ASAP7_75t_L g889 ( .A(n_113), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g1616 ( .A1(n_114), .A2(n_274), .B1(n_1552), .B2(n_1560), .Y(n_1616) );
AO221x1_ASAP7_75t_L g1023 ( .A1(n_115), .A2(n_201), .B1(n_433), .B2(n_719), .C(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1038 ( .A(n_115), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_116), .A2(n_275), .B1(n_483), .B2(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1374 ( .A(n_116), .Y(n_1374) );
INVx1_ASAP7_75t_L g955 ( .A(n_117), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_117), .A2(n_223), .B1(n_591), .B2(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g958 ( .A(n_119), .Y(n_958) );
AO22x2_ASAP7_75t_L g934 ( .A1(n_122), .A2(n_935), .B1(n_936), .B2(n_990), .Y(n_934) );
INVxp67_ASAP7_75t_SL g935 ( .A(n_122), .Y(n_935) );
INVx1_ASAP7_75t_L g1250 ( .A(n_125), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1264 ( .A1(n_125), .A2(n_642), .B1(n_661), .B2(n_1265), .C(n_1268), .Y(n_1264) );
INVx1_ASAP7_75t_L g1611 ( .A(n_126), .Y(n_1611) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_127), .A2(n_285), .B1(n_694), .B2(n_1000), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_127), .A2(n_285), .B1(n_769), .B2(n_1019), .C(n_1020), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_128), .A2(n_203), .B1(n_629), .B2(n_630), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_128), .A2(n_203), .B1(n_694), .B2(n_696), .Y(n_981) );
INVx1_ASAP7_75t_L g883 ( .A(n_129), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g1202 ( .A(n_130), .Y(n_1202) );
OA22x2_ASAP7_75t_L g1430 ( .A1(n_132), .A2(n_1431), .B1(n_1487), .B2(n_1488), .Y(n_1430) );
INVxp67_ASAP7_75t_SL g1488 ( .A(n_132), .Y(n_1488) );
INVx1_ASAP7_75t_L g1179 ( .A(n_134), .Y(n_1179) );
OAI22xp33_ASAP7_75t_L g1189 ( .A1(n_134), .A2(n_200), .B1(n_866), .B2(n_869), .Y(n_1189) );
XNOR2xp5_ASAP7_75t_L g528 ( .A(n_135), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g1404 ( .A(n_136), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_137), .A2(n_170), .B1(n_474), .B2(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g519 ( .A(n_137), .Y(n_519) );
INVx1_ASAP7_75t_L g1349 ( .A(n_139), .Y(n_1349) );
INVx1_ASAP7_75t_L g1157 ( .A(n_140), .Y(n_1157) );
OAI221xp5_ASAP7_75t_L g1168 ( .A1(n_140), .A2(n_642), .B1(n_661), .B2(n_1169), .C(n_1171), .Y(n_1168) );
INVx1_ASAP7_75t_L g1500 ( .A(n_141), .Y(n_1500) );
INVx1_ASAP7_75t_L g1113 ( .A(n_142), .Y(n_1113) );
AOI22xp33_ASAP7_75t_SL g1131 ( .A1(n_142), .A2(n_309), .B1(n_696), .B2(n_985), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_143), .A2(n_164), .B1(n_591), .B2(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g732 ( .A(n_143), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g1862 ( .A(n_144), .Y(n_1862) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_145), .A2(n_199), .B1(n_590), .B2(n_591), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_145), .A2(n_199), .B1(n_664), .B2(n_666), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_146), .Y(n_553) );
INVx1_ASAP7_75t_L g742 ( .A(n_147), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_148), .Y(n_1442) );
INVx1_ASAP7_75t_L g1504 ( .A(n_149), .Y(n_1504) );
CKINVDCx5p33_ASAP7_75t_R g1517 ( .A(n_150), .Y(n_1517) );
INVx1_ASAP7_75t_L g962 ( .A(n_151), .Y(n_962) );
INVx1_ASAP7_75t_L g1557 ( .A(n_153), .Y(n_1557) );
OAI22xp33_ASAP7_75t_L g1211 ( .A1(n_154), .A2(n_325), .B1(n_828), .B2(n_830), .Y(n_1211) );
INVx1_ASAP7_75t_L g1230 ( .A(n_154), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1824 ( .A1(n_156), .A2(n_256), .B1(n_630), .B2(n_1825), .Y(n_1824) );
AOI22xp33_ASAP7_75t_L g1833 ( .A1(n_156), .A2(n_256), .B1(n_985), .B2(n_1291), .Y(n_1833) );
INVx1_ASAP7_75t_L g1108 ( .A(n_157), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_157), .A2(n_195), .B1(n_480), .B2(n_555), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_158), .A2(n_340), .B1(n_821), .B2(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1216 ( .A(n_158), .Y(n_1216) );
AOI221xp5_ASAP7_75t_L g1550 ( .A1(n_159), .A2(n_246), .B1(n_1551), .B2(n_1558), .C(n_1561), .Y(n_1550) );
INVx1_ASAP7_75t_L g1392 ( .A(n_161), .Y(n_1392) );
INVx1_ASAP7_75t_L g1056 ( .A(n_163), .Y(n_1056) );
INVx1_ASAP7_75t_L g733 ( .A(n_164), .Y(n_733) );
INVx1_ASAP7_75t_L g1243 ( .A(n_165), .Y(n_1243) );
INVx1_ASAP7_75t_L g1555 ( .A(n_166), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_166), .B(n_1568), .Y(n_1573) );
AOI221xp5_ASAP7_75t_L g1514 ( .A1(n_167), .A2(n_301), .B1(n_715), .B2(n_1515), .C(n_1516), .Y(n_1514) );
INVx1_ASAP7_75t_L g1525 ( .A(n_167), .Y(n_1525) );
INVx1_ASAP7_75t_L g1209 ( .A(n_168), .Y(n_1209) );
OAI211xp5_ASAP7_75t_SL g1223 ( .A1(n_168), .A2(n_613), .B(n_1224), .C(n_1229), .Y(n_1223) );
INVx1_ASAP7_75t_L g391 ( .A(n_169), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_169), .A2(n_190), .B1(n_453), .B2(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g494 ( .A(n_170), .Y(n_494) );
INVx2_ASAP7_75t_L g361 ( .A(n_171), .Y(n_361) );
AO221x2_ASAP7_75t_L g1591 ( .A1(n_172), .A2(n_218), .B1(n_1552), .B2(n_1592), .C(n_1593), .Y(n_1591) );
INVx1_ASAP7_75t_L g1101 ( .A(n_173), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_174), .A2(n_207), .B1(n_830), .B2(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1184 ( .A(n_174), .Y(n_1184) );
INVx1_ASAP7_75t_L g918 ( .A(n_175), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_176), .A2(n_272), .B1(n_715), .B2(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_176), .A2(n_272), .B1(n_576), .B2(n_591), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g1461 ( .A(n_177), .Y(n_1461) );
BUFx3_ASAP7_75t_L g381 ( .A(n_178), .Y(n_381) );
INVx1_ASAP7_75t_L g397 ( .A(n_178), .Y(n_397) );
INVx1_ASAP7_75t_L g1227 ( .A(n_179), .Y(n_1227) );
OAI22xp33_ASAP7_75t_L g1233 ( .A1(n_179), .A2(n_270), .B1(n_543), .B2(n_1188), .Y(n_1233) );
CKINVDCx5p33_ASAP7_75t_R g1452 ( .A(n_180), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_181), .Y(n_1027) );
INVx1_ASAP7_75t_L g1061 ( .A(n_182), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_183), .Y(n_1443) );
OAI22xp5_ASAP7_75t_L g1872 ( .A1(n_184), .A2(n_314), .B1(n_835), .B2(n_836), .Y(n_1872) );
INVx1_ASAP7_75t_L g1882 ( .A(n_184), .Y(n_1882) );
INVx1_ASAP7_75t_L g690 ( .A(n_185), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g1102 ( .A1(n_186), .A2(n_254), .B1(n_684), .B2(n_1103), .C(n_1104), .Y(n_1102) );
INVx1_ASAP7_75t_L g1111 ( .A(n_186), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_187), .A2(n_233), .B1(n_784), .B2(n_785), .Y(n_783) );
INVx1_ASAP7_75t_L g1159 ( .A(n_188), .Y(n_1159) );
OAI211xp5_ASAP7_75t_SL g1174 ( .A1(n_188), .A2(n_613), .B(n_1175), .C(n_1183), .Y(n_1174) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_189), .Y(n_1009) );
INVx1_ASAP7_75t_L g416 ( .A(n_190), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_191), .A2(n_342), .B1(n_555), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1013 ( .A(n_191), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g1409 ( .A(n_192), .Y(n_1409) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_193), .A2(n_202), .B1(n_1291), .B2(n_1292), .C(n_1293), .Y(n_1290) );
INVx1_ASAP7_75t_L g1347 ( .A(n_193), .Y(n_1347) );
AOI221xp5_ASAP7_75t_L g858 ( .A1(n_194), .A2(n_343), .B1(n_438), .B2(n_633), .C(n_769), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_194), .A2(n_289), .B1(n_866), .B2(n_869), .Y(n_865) );
INVx1_ASAP7_75t_L g1109 ( .A(n_195), .Y(n_1109) );
INVx1_ASAP7_75t_L g408 ( .A(n_196), .Y(n_408) );
INVx1_ASAP7_75t_L g914 ( .A(n_198), .Y(n_914) );
INVx1_ASAP7_75t_L g1040 ( .A(n_201), .Y(n_1040) );
INVx1_ASAP7_75t_L g1344 ( .A(n_202), .Y(n_1344) );
INVx1_ASAP7_75t_L g422 ( .A(n_204), .Y(n_422) );
INVx1_ASAP7_75t_L g540 ( .A(n_204), .Y(n_540) );
INVxp33_ASAP7_75t_L g1086 ( .A(n_205), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_206), .A2(n_279), .B1(n_866), .B2(n_869), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_206), .A2(n_245), .B1(n_1019), .B2(n_1024), .C(n_1222), .Y(n_1277) );
INVx1_ASAP7_75t_L g1185 ( .A(n_207), .Y(n_1185) );
INVxp67_ASAP7_75t_L g1820 ( .A(n_208), .Y(n_1820) );
AOI22xp33_ASAP7_75t_L g1838 ( .A1(n_208), .A2(n_296), .B1(n_803), .B2(n_1204), .Y(n_1838) );
CKINVDCx5p33_ASAP7_75t_R g1465 ( .A(n_211), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1406 ( .A(n_212), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_213), .A2(n_320), .B1(n_696), .B2(n_1002), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1022 ( .A1(n_213), .A2(n_613), .B1(n_1023), .B2(n_1025), .C(n_1028), .Y(n_1022) );
INVx1_ASAP7_75t_L g817 ( .A(n_214), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g837 ( .A1(n_214), .A2(n_642), .B1(n_838), .B2(n_844), .C(n_847), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_215), .Y(n_1410) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_216), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_217), .Y(n_384) );
XOR2xp5_ASAP7_75t_L g1384 ( .A(n_218), .B(n_1385), .Y(n_1384) );
INVx1_ASAP7_75t_L g1105 ( .A(n_219), .Y(n_1105) );
INVx1_ASAP7_75t_L g1399 ( .A(n_220), .Y(n_1399) );
AOI221xp5_ASAP7_75t_L g1422 ( .A1(n_220), .A2(n_234), .B1(n_1291), .B2(n_1313), .C(n_1423), .Y(n_1422) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_221), .A2(n_283), .B1(n_1581), .B2(n_1584), .Y(n_1580) );
CKINVDCx5p33_ASAP7_75t_R g1496 ( .A(n_222), .Y(n_1496) );
INVx1_ASAP7_75t_L g954 ( .A(n_223), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g1871 ( .A(n_224), .Y(n_1871) );
OAI221xp5_ASAP7_75t_L g1883 ( .A1(n_224), .A2(n_561), .B1(n_570), .B2(n_595), .C(n_1884), .Y(n_1883) );
AOI22xp5_ASAP7_75t_L g1604 ( .A1(n_225), .A2(n_300), .B1(n_1560), .B2(n_1587), .Y(n_1604) );
INVx1_ASAP7_75t_L g1393 ( .A(n_226), .Y(n_1393) );
CKINVDCx5p33_ASAP7_75t_R g1494 ( .A(n_227), .Y(n_1494) );
INVx1_ASAP7_75t_L g893 ( .A(n_228), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g1245 ( .A(n_230), .Y(n_1245) );
INVx1_ASAP7_75t_L g1253 ( .A(n_231), .Y(n_1253) );
INVx1_ASAP7_75t_L g765 ( .A(n_232), .Y(n_765) );
INVx1_ASAP7_75t_L g1403 ( .A(n_234), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_235), .Y(n_1100) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_236), .A2(n_319), .B1(n_828), .B2(n_830), .Y(n_891) );
INVx1_ASAP7_75t_L g925 ( .A(n_236), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g1510 ( .A(n_237), .Y(n_1510) );
INVx1_ASAP7_75t_L g1612 ( .A(n_238), .Y(n_1612) );
CKINVDCx16_ASAP7_75t_R g1048 ( .A(n_240), .Y(n_1048) );
INVx1_ASAP7_75t_L g1197 ( .A(n_242), .Y(n_1197) );
CKINVDCx20_ASAP7_75t_R g1594 ( .A(n_243), .Y(n_1594) );
INVx1_ASAP7_75t_L g886 ( .A(n_244), .Y(n_886) );
OAI221xp5_ASAP7_75t_L g896 ( .A1(n_244), .A2(n_642), .B1(n_847), .B2(n_897), .C(n_903), .Y(n_896) );
INVx1_ASAP7_75t_L g653 ( .A(n_247), .Y(n_653) );
INVx1_ASAP7_75t_L g1241 ( .A(n_248), .Y(n_1241) );
INVx1_ASAP7_75t_L g412 ( .A(n_249), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_249), .A2(n_333), .B1(n_432), .B2(n_436), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g1864 ( .A(n_251), .Y(n_1864) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_252), .A2(n_276), .B1(n_1435), .B2(n_1437), .Y(n_1434) );
INVx1_ASAP7_75t_L g1471 ( .A(n_252), .Y(n_1471) );
INVx1_ASAP7_75t_L g1201 ( .A(n_253), .Y(n_1201) );
AOI21xp33_ASAP7_75t_L g1221 ( .A1(n_253), .A2(n_1020), .B(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1112 ( .A(n_254), .Y(n_1112) );
AOI21xp33_ASAP7_75t_L g1859 ( .A1(n_255), .A2(n_610), .B(n_1020), .Y(n_1859) );
INVx1_ASAP7_75t_L g516 ( .A(n_257), .Y(n_516) );
INVx1_ASAP7_75t_L g1331 ( .A(n_258), .Y(n_1331) );
OAI211xp5_ASAP7_75t_L g1438 ( .A1(n_260), .A2(n_645), .B(n_968), .C(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1468 ( .A(n_260), .Y(n_1468) );
INVx1_ASAP7_75t_L g1052 ( .A(n_261), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1325 ( .A(n_262), .Y(n_1325) );
XNOR2xp5_ASAP7_75t_L g1194 ( .A(n_263), .B(n_1195), .Y(n_1194) );
INVxp33_ASAP7_75t_L g1817 ( .A(n_264), .Y(n_1817) );
INVx1_ASAP7_75t_L g877 ( .A(n_265), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g1210 ( .A1(n_266), .A2(n_291), .B1(n_803), .B2(n_1079), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_266), .A2(n_291), .B1(n_664), .B2(n_666), .Y(n_1213) );
BUFx3_ASAP7_75t_L g382 ( .A(n_267), .Y(n_382) );
INVx1_ASAP7_75t_L g419 ( .A(n_267), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g1497 ( .A(n_268), .Y(n_1497) );
INVx1_ASAP7_75t_L g1261 ( .A(n_269), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_271), .Y(n_1008) );
AO22x2_ASAP7_75t_L g1093 ( .A1(n_273), .A2(n_1094), .B1(n_1133), .B2(n_1134), .Y(n_1093) );
INVxp67_ASAP7_75t_L g1133 ( .A(n_273), .Y(n_1133) );
XNOR2xp5_ASAP7_75t_L g1236 ( .A(n_274), .B(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1366 ( .A(n_275), .Y(n_1366) );
INVx1_ASAP7_75t_L g1470 ( .A(n_276), .Y(n_1470) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_277), .Y(n_357) );
INVx1_ASAP7_75t_L g465 ( .A(n_277), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_277), .B(n_327), .Y(n_609) );
AND2x2_ASAP7_75t_L g617 ( .A(n_277), .B(n_464), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_278), .Y(n_1026) );
INVx1_ASAP7_75t_L g1275 ( .A(n_279), .Y(n_1275) );
AOI21xp33_ASAP7_75t_L g1865 ( .A1(n_280), .A2(n_433), .B(n_1024), .Y(n_1865) );
INVx1_ASAP7_75t_L g1886 ( .A(n_280), .Y(n_1886) );
XNOR2xp5_ASAP7_75t_L g676 ( .A(n_281), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g378 ( .A(n_282), .Y(n_378) );
OR2x2_ASAP7_75t_L g539 ( .A(n_282), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g1799 ( .A(n_283), .Y(n_1799) );
AOI22xp33_ASAP7_75t_L g1843 ( .A1(n_283), .A2(n_1844), .B1(n_1848), .B2(n_1888), .Y(n_1843) );
CKINVDCx5p33_ASAP7_75t_R g1328 ( .A(n_284), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_286), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g1855 ( .A(n_287), .Y(n_1855) );
CKINVDCx5p33_ASAP7_75t_R g1457 ( .A(n_288), .Y(n_1457) );
INVx1_ASAP7_75t_L g853 ( .A(n_289), .Y(n_853) );
INVx1_ASAP7_75t_L g541 ( .A(n_290), .Y(n_541) );
INVx1_ASAP7_75t_L g857 ( .A(n_292), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_292), .A2(n_343), .B1(n_536), .B2(n_543), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g1861 ( .A(n_293), .Y(n_1861) );
INVx1_ASAP7_75t_L g822 ( .A(n_294), .Y(n_822) );
INVx1_ASAP7_75t_L g950 ( .A(n_295), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_295), .A2(n_308), .B1(n_704), .B2(n_842), .Y(n_973) );
INVx1_ASAP7_75t_L g1818 ( .A(n_296), .Y(n_1818) );
CKINVDCx5p33_ASAP7_75t_R g1466 ( .A(n_297), .Y(n_1466) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_298), .A2(n_313), .B1(n_696), .B2(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g735 ( .A(n_298), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g1807 ( .A1(n_299), .A2(n_326), .B1(n_684), .B2(n_940), .Y(n_1807) );
OAI22xp5_ASAP7_75t_L g1815 ( .A1(n_299), .A2(n_326), .B1(n_502), .B2(n_730), .Y(n_1815) );
AOI22x1_ASAP7_75t_L g992 ( .A1(n_300), .A2(n_993), .B1(n_994), .B2(n_1041), .Y(n_992) );
INVxp67_ASAP7_75t_SL g1041 ( .A(n_300), .Y(n_1041) );
INVx1_ASAP7_75t_L g1523 ( .A(n_301), .Y(n_1523) );
INVx1_ASAP7_75t_L g946 ( .A(n_303), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_304), .A2(n_328), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1167 ( .A1(n_304), .A2(n_328), .B1(n_835), .B2(n_836), .Y(n_1167) );
INVx1_ASAP7_75t_L g1138 ( .A(n_305), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_306), .A2(n_338), .B1(n_711), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_306), .A2(n_338), .B1(n_401), .B2(n_694), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_307), .Y(n_568) );
INVx1_ASAP7_75t_L g949 ( .A(n_308), .Y(n_949) );
INVx1_ASAP7_75t_L g1118 ( .A(n_309), .Y(n_1118) );
INVx1_ASAP7_75t_L g1181 ( .A(n_310), .Y(n_1181) );
OAI22xp33_ASAP7_75t_L g1256 ( .A1(n_311), .A2(n_331), .B1(n_828), .B2(n_830), .Y(n_1256) );
INVx1_ASAP7_75t_L g1280 ( .A(n_311), .Y(n_1280) );
INVx1_ASAP7_75t_L g659 ( .A(n_312), .Y(n_659) );
INVx1_ASAP7_75t_L g727 ( .A(n_313), .Y(n_727) );
INVx1_ASAP7_75t_L g1881 ( .A(n_314), .Y(n_1881) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
AND3x2_ASAP7_75t_L g1556 ( .A(n_315), .B(n_349), .C(n_1557), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_315), .B(n_349), .Y(n_1566) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_316), .Y(n_832) );
INVx2_ASAP7_75t_L g362 ( .A(n_317), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_318), .Y(n_881) );
INVx1_ASAP7_75t_L g923 ( .A(n_319), .Y(n_923) );
INVx1_ASAP7_75t_L g1021 ( .A(n_320), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_321), .Y(n_745) );
XNOR2xp5_ASAP7_75t_L g871 ( .A(n_322), .B(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g599 ( .A(n_323), .Y(n_599) );
INVx1_ASAP7_75t_L g686 ( .A(n_324), .Y(n_686) );
INVx1_ASAP7_75t_L g1231 ( .A(n_325), .Y(n_1231) );
INVx1_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
INVx2_ASAP7_75t_L g464 ( .A(n_327), .Y(n_464) );
AO22x2_ASAP7_75t_L g1490 ( .A1(n_329), .A2(n_1491), .B1(n_1539), .B2(n_1540), .Y(n_1490) );
INVxp67_ASAP7_75t_SL g1539 ( .A(n_329), .Y(n_1539) );
CKINVDCx5p33_ASAP7_75t_R g1433 ( .A(n_330), .Y(n_1433) );
INVx1_ASAP7_75t_L g1279 ( .A(n_331), .Y(n_1279) );
INVx1_ASAP7_75t_L g399 ( .A(n_333), .Y(n_399) );
INVx1_ASAP7_75t_L g1870 ( .A(n_334), .Y(n_1870) );
HB1xp67_ASAP7_75t_L g1884 ( .A(n_334), .Y(n_1884) );
OAI211xp5_ASAP7_75t_L g1447 ( .A1(n_335), .A2(n_747), .B(n_1448), .C(n_1449), .Y(n_1447) );
INVx1_ASAP7_75t_L g1485 ( .A(n_335), .Y(n_1485) );
INVx1_ASAP7_75t_L g860 ( .A(n_336), .Y(n_860) );
OAI211xp5_ASAP7_75t_SL g612 ( .A1(n_337), .A2(n_613), .B(n_618), .C(n_635), .Y(n_612) );
INVx1_ASAP7_75t_L g1147 ( .A(n_339), .Y(n_1147) );
INVx1_ASAP7_75t_L g1218 ( .A(n_340), .Y(n_1218) );
INVxp33_ASAP7_75t_SL g1172 ( .A(n_341), .Y(n_1172) );
INVx1_ASAP7_75t_L g1014 ( .A(n_342), .Y(n_1014) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_365), .B(n_1543), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_352), .Y(n_346) );
AND2x4_ASAP7_75t_L g1842 ( .A(n_347), .B(n_353), .Y(n_1842) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_SL g1847 ( .A(n_348), .Y(n_1847) );
NAND2xp5_ASAP7_75t_L g1891 ( .A(n_348), .B(n_350), .Y(n_1891) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g1846 ( .A(n_350), .B(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_358), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g522 ( .A(n_355), .B(n_489), .Y(n_522) );
OR2x6_ASAP7_75t_L g736 ( .A(n_355), .B(n_489), .Y(n_736) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g430 ( .A(n_356), .B(n_364), .Y(n_430) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_357), .B(n_511), .Y(n_1020) );
INVx8_ASAP7_75t_L g518 ( .A(n_358), .Y(n_518) );
OR2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_363), .Y(n_358) );
OR2x6_ASAP7_75t_L g521 ( .A(n_359), .B(n_510), .Y(n_521) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_359), .Y(n_652) );
INVx2_ASAP7_75t_SL g906 ( .A(n_359), .Y(n_906) );
INVx1_ASAP7_75t_L g913 ( .A(n_359), .Y(n_913) );
BUFx2_ASAP7_75t_L g1271 ( .A(n_359), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_359), .B(n_1335), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g435 ( .A(n_361), .B(n_362), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_361), .Y(n_440) );
INVx2_ASAP7_75t_L g445 ( .A(n_361), .Y(n_445) );
AND2x4_ASAP7_75t_L g451 ( .A(n_361), .B(n_441), .Y(n_451) );
INVx1_ASAP7_75t_L g507 ( .A(n_361), .Y(n_507) );
INVx2_ASAP7_75t_L g441 ( .A(n_362), .Y(n_441) );
INVx1_ASAP7_75t_L g447 ( .A(n_362), .Y(n_447) );
INVx1_ASAP7_75t_L g504 ( .A(n_362), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_362), .B(n_445), .Y(n_622) );
INVx1_ASAP7_75t_L g648 ( .A(n_362), .Y(n_648) );
AND2x4_ASAP7_75t_L g503 ( .A(n_363), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g505 ( .A(n_364), .B(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g730 ( .A(n_364), .B(n_506), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_1380), .B2(n_1381), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
XNOR2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_1042), .Y(n_367) );
XNOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_673), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_525), .B1(n_671), .B2(n_672), .Y(n_369) );
INVx2_ASAP7_75t_L g671 ( .A(n_370), .Y(n_671) );
INVx1_ASAP7_75t_L g524 ( .A(n_371), .Y(n_524) );
AOI211x1_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_420), .B(n_425), .C(n_492), .Y(n_371) );
NAND4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_383), .C(n_398), .D(n_411), .Y(n_372) );
BUFx2_ASAP7_75t_L g1529 ( .A(n_373), .Y(n_1529) );
NAND4xp25_ASAP7_75t_L g1801 ( .A(n_373), .B(n_1802), .C(n_1805), .D(n_1808), .Y(n_1801) );
INVx5_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_374), .A2(n_680), .B(n_681), .C(n_682), .Y(n_679) );
CKINVDCx8_ASAP7_75t_R g747 ( .A(n_374), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_374), .B(n_939), .Y(n_938) );
AOI211xp5_ASAP7_75t_L g1081 ( .A1(n_374), .A2(n_1082), .B(n_1083), .C(n_1084), .Y(n_1081) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_379), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g1104 ( .A1(n_375), .A2(n_476), .B(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x6_ASAP7_75t_L g417 ( .A(n_376), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g753 ( .A(n_376), .Y(n_753) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_376), .B(n_401), .Y(n_1083) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x6_ASAP7_75t_L g409 ( .A(n_377), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_378), .Y(n_387) );
INVx1_ASAP7_75t_L g394 ( .A(n_378), .Y(n_394) );
AND2x2_ASAP7_75t_L g470 ( .A(n_378), .B(n_422), .Y(n_470) );
INVx2_ASAP7_75t_L g491 ( .A(n_378), .Y(n_491) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_379), .Y(n_476) );
INVx2_ASAP7_75t_L g697 ( .A(n_379), .Y(n_697) );
INVx1_ASAP7_75t_L g798 ( .A(n_379), .Y(n_798) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_380), .Y(n_585) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx2_ASAP7_75t_L g389 ( .A(n_381), .Y(n_389) );
AND2x4_ASAP7_75t_L g418 ( .A(n_381), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g390 ( .A(n_382), .Y(n_390) );
AND2x4_ASAP7_75t_L g396 ( .A(n_382), .B(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_391), .B2(n_392), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_384), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_385), .A2(n_413), .B1(n_686), .B2(n_687), .Y(n_685) );
INVx4_ASAP7_75t_L g755 ( .A(n_385), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_385), .A2(n_413), .B1(n_946), .B2(n_947), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_385), .A2(n_1056), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1099 ( .A1(n_385), .A2(n_417), .B1(n_1100), .B2(n_1101), .C(n_1102), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_385), .A2(n_392), .B1(n_1494), .B2(n_1525), .Y(n_1524) );
AOI22xp5_ASAP7_75t_SL g1802 ( .A1(n_385), .A2(n_1087), .B1(n_1803), .B2(n_1804), .Y(n_1802) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AND2x4_ASAP7_75t_L g404 ( .A(n_386), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_SL g1453 ( .A(n_386), .B(n_405), .Y(n_1453) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx6_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
INVx2_ASAP7_75t_L g484 ( .A(n_388), .Y(n_484) );
BUFx2_ASAP7_75t_L g582 ( .A(n_388), .Y(n_582) );
AND2x2_ASAP7_75t_L g602 ( .A(n_388), .B(n_566), .Y(n_602) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g410 ( .A(n_389), .Y(n_410) );
INVx1_ASAP7_75t_L g407 ( .A(n_390), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_392), .A2(n_417), .B1(n_689), .B2(n_690), .Y(n_688) );
INVx4_ASAP7_75t_L g750 ( .A(n_392), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_392), .A2(n_417), .B1(n_949), .B2(n_950), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_392), .A2(n_417), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_392), .A2(n_413), .B1(n_1097), .B2(n_1098), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g1808 ( .A1(n_392), .A2(n_417), .B1(n_1809), .B2(n_1810), .Y(n_1808) );
AND2x6_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AND2x4_ASAP7_75t_L g413 ( .A(n_393), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_393), .B(n_414), .Y(n_1087) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g941 ( .A(n_394), .B(n_942), .Y(n_941) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_395), .Y(n_1006) );
BUFx6f_ASAP7_75t_L g1079 ( .A(n_395), .Y(n_1079) );
INVx2_ASAP7_75t_L g1163 ( .A(n_395), .Y(n_1163) );
BUFx6f_ASAP7_75t_L g1204 ( .A(n_395), .Y(n_1204) );
INVx1_ASAP7_75t_L g1472 ( .A(n_395), .Y(n_1472) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_396), .Y(n_481) );
INVx1_ASAP7_75t_L g537 ( .A(n_396), .Y(n_537) );
INVx2_ASAP7_75t_L g580 ( .A(n_396), .Y(n_580) );
INVx1_ASAP7_75t_L g780 ( .A(n_396), .Y(n_780) );
INVx1_ASAP7_75t_L g546 ( .A(n_397), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_402), .B2(n_403), .C1(n_408), .C2(n_409), .Y(n_398) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_401), .Y(n_681) );
HB1xp67_ASAP7_75t_L g1416 ( .A(n_401), .Y(n_1416) );
AOI222xp33_ASAP7_75t_L g1526 ( .A1(n_403), .A2(n_409), .B1(n_1512), .B2(n_1513), .C1(n_1517), .C2(n_1527), .Y(n_1526) );
BUFx4f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g683 ( .A(n_404), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_404), .A2(n_409), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g942 ( .A(n_406), .Y(n_942) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g563 ( .A(n_407), .Y(n_563) );
INVx3_ASAP7_75t_L g684 ( .A(n_409), .Y(n_684) );
AOI322xp5_ASAP7_75t_L g1449 ( .A1(n_409), .A2(n_1442), .A3(n_1443), .B1(n_1450), .B2(n_1451), .C1(n_1452), .C2(n_1453), .Y(n_1449) );
BUFx3_ASAP7_75t_L g572 ( .A(n_410), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_416), .B2(n_417), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_413), .A2(n_417), .B1(n_1522), .B2(n_1523), .Y(n_1521) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_415), .Y(n_588) );
INVx2_ASAP7_75t_L g695 ( .A(n_415), .Y(n_695) );
INVx1_ASAP7_75t_L g985 ( .A(n_415), .Y(n_985) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_415), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1877 ( .A(n_415), .Y(n_1877) );
CKINVDCx6p67_ASAP7_75t_R g749 ( .A(n_417), .Y(n_749) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_418), .Y(n_479) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_418), .Y(n_487) );
INVx2_ASAP7_75t_SL g556 ( .A(n_418), .Y(n_556) );
BUFx2_ASAP7_75t_L g576 ( .A(n_418), .Y(n_576) );
BUFx3_ASAP7_75t_L g803 ( .A(n_418), .Y(n_803) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_418), .Y(n_821) );
BUFx2_ASAP7_75t_L g987 ( .A(n_418), .Y(n_987) );
BUFx6f_ASAP7_75t_L g1450 ( .A(n_418), .Y(n_1450) );
INVx1_ASAP7_75t_L g547 ( .A(n_419), .Y(n_547) );
AO211x2_ASAP7_75t_L g677 ( .A1(n_420), .A2(n_678), .B(n_691), .C(n_725), .Y(n_677) );
BUFx6f_ASAP7_75t_L g951 ( .A(n_420), .Y(n_951) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
AND2x4_ASAP7_75t_L g756 ( .A(n_421), .B(n_423), .Y(n_756) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g490 ( .A(n_422), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g1036 ( .A(n_423), .Y(n_1036) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g429 ( .A(n_424), .Y(n_429) );
OR2x6_ASAP7_75t_L g1364 ( .A(n_424), .B(n_1020), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_466), .Y(n_425) );
AOI33xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_431), .A3(n_442), .B1(n_452), .B2(n_457), .B3(n_458), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_428), .B(n_714), .C(n_717), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g1822 ( .A(n_428), .B(n_1823), .C(n_1824), .Y(n_1822) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OR2x6_ASAP7_75t_L g468 ( .A(n_429), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g604 ( .A(n_429), .Y(n_604) );
BUFx2_ASAP7_75t_L g670 ( .A(n_429), .Y(n_670) );
OR2x2_ASAP7_75t_L g700 ( .A(n_429), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g767 ( .A(n_429), .B(n_430), .Y(n_767) );
OR2x2_ASAP7_75t_L g800 ( .A(n_429), .B(n_469), .Y(n_800) );
AND2x2_ASAP7_75t_L g1831 ( .A(n_429), .B(n_634), .Y(n_1831) );
INVx1_ASAP7_75t_L g655 ( .A(n_430), .Y(n_655) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g610 ( .A(n_434), .Y(n_610) );
INVx2_ASAP7_75t_SL g1222 ( .A(n_434), .Y(n_1222) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_435), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g726 ( .A1(n_436), .A2(n_498), .B(n_727), .C(n_728), .Y(n_726) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g959 ( .A(n_437), .Y(n_959) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx6f_ASAP7_75t_L g1065 ( .A(n_438), .Y(n_1065) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g497 ( .A(n_439), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_439), .B(n_499), .Y(n_498) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_439), .Y(n_719) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_439), .Y(n_1019) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_439), .Y(n_1116) );
INVx1_ASAP7_75t_L g1826 ( .A(n_439), .Y(n_1826) );
AND2x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_444), .Y(n_455) );
AND2x4_ASAP7_75t_L g509 ( .A(n_444), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g665 ( .A(n_444), .B(n_617), .Y(n_665) );
INVx1_ASAP7_75t_L g705 ( .A(n_444), .Y(n_705) );
BUFx2_ASAP7_75t_L g715 ( .A(n_444), .Y(n_715) );
BUFx6f_ASAP7_75t_L g1017 ( .A(n_444), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g1829 ( .A(n_444), .Y(n_1829) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g640 ( .A(n_445), .Y(n_640) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_449), .A2(n_658), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
OAI221xp5_ASAP7_75t_L g1224 ( .A1(n_449), .A2(n_1225), .B1(n_1226), .B2(n_1227), .C(n_1228), .Y(n_1224) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_449), .A2(n_1274), .B1(n_1275), .B2(n_1276), .C(n_1277), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_449), .A2(n_1301), .B1(n_1328), .B2(n_1370), .Y(n_1375) );
INVx2_ASAP7_75t_L g1515 ( .A(n_449), .Y(n_1515) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g456 ( .A(n_450), .Y(n_456) );
INVx2_ASAP7_75t_SL g1373 ( .A(n_450), .Y(n_1373) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g515 ( .A(n_451), .Y(n_515) );
INVx1_ASAP7_75t_L g627 ( .A(n_451), .Y(n_627) );
INVx3_ASAP7_75t_L g709 ( .A(n_451), .Y(n_709) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_455), .B(n_1343), .Y(n_1350) );
AOI33xp33_ASAP7_75t_L g766 ( .A1(n_458), .A2(n_767), .A3(n_768), .B1(n_772), .B2(n_773), .B3(n_774), .Y(n_766) );
AOI33xp33_ASAP7_75t_L g1063 ( .A1(n_458), .A2(n_767), .A3(n_1064), .B1(n_1066), .B2(n_1068), .B3(n_1070), .Y(n_1063) );
INVx2_ASAP7_75t_L g1486 ( .A(n_458), .Y(n_1486) );
INVx6_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx5_ASAP7_75t_L g712 ( .A(n_459), .Y(n_712) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_460), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g538 ( .A(n_461), .B(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g1343 ( .A(n_461), .B(n_617), .Y(n_1343) );
INVx2_ASAP7_75t_L g634 ( .A(n_462), .Y(n_634) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_462), .Y(n_1024) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g511 ( .A(n_464), .Y(n_511) );
AOI33xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_471), .A3(n_477), .B1(n_482), .B2(n_485), .B3(n_488), .Y(n_466) );
AOI33xp33_ASAP7_75t_L g775 ( .A1(n_467), .A2(n_488), .A3(n_776), .B1(n_781), .B2(n_783), .B3(n_786), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g574 ( .A(n_468), .Y(n_574) );
OAI22xp5_ASAP7_75t_SL g1144 ( .A1(n_468), .A2(n_1145), .B1(n_1153), .B2(n_1155), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1530 ( .A1(n_468), .A2(n_1153), .B1(n_1531), .B2(n_1537), .Y(n_1530) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g701 ( .A(n_470), .Y(n_701) );
INVx2_ASAP7_75t_SL g1315 ( .A(n_470), .Y(n_1315) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_473), .Y(n_784) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_476), .Y(n_785) );
INVx1_ASAP7_75t_L g1312 ( .A(n_476), .Y(n_1312) );
AND2x4_ASAP7_75t_L g1321 ( .A(n_476), .B(n_1322), .Y(n_1321) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_SL g778 ( .A(n_479), .Y(n_778) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_479), .B(n_1300), .Y(n_1299) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g878 ( .A(n_481), .Y(n_878) );
INVx1_ASAP7_75t_L g1242 ( .A(n_481), .Y(n_1242) );
BUFx3_ASAP7_75t_L g1317 ( .A(n_481), .Y(n_1317) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_SL g551 ( .A(n_484), .Y(n_551) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx4f_ASAP7_75t_L g590 ( .A(n_487), .Y(n_590) );
INVx1_ASAP7_75t_L g870 ( .A(n_487), .Y(n_870) );
INVx4_ASAP7_75t_L g826 ( .A(n_488), .Y(n_826) );
BUFx4f_ASAP7_75t_L g1154 ( .A(n_488), .Y(n_1154) );
AOI221xp5_ASAP7_75t_L g1874 ( .A1(n_488), .A2(n_574), .B1(n_1875), .B2(n_1879), .C(n_1883), .Y(n_1874) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AND2x4_ASAP7_75t_L g592 ( .A(n_489), .B(n_490), .Y(n_592) );
AND2x4_ASAP7_75t_L g601 ( .A(n_489), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g1294 ( .A(n_490), .Y(n_1294) );
AND2x4_ASAP7_75t_L g566 ( .A(n_491), .B(n_567), .Y(n_566) );
AOI31xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_508), .A3(n_517), .B(n_522), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_498), .C(n_501), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g629 ( .A(n_496), .Y(n_629) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g614 ( .A(n_497), .B(n_615), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_498), .B(n_759), .C(n_762), .Y(n_758) );
CKINVDCx11_ASAP7_75t_R g968 ( .A(n_498), .Y(n_968) );
AOI211xp5_ASAP7_75t_L g1812 ( .A1(n_498), .A2(n_1813), .B(n_1814), .C(n_1815), .Y(n_1812) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g965 ( .A(n_500), .Y(n_965) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g729 ( .A(n_503), .Y(n_729) );
INVx2_ASAP7_75t_L g760 ( .A(n_503), .Y(n_760) );
AOI222xp33_ASAP7_75t_L g1110 ( .A1(n_503), .A2(n_963), .B1(n_1111), .B2(n_1112), .C1(n_1113), .C2(n_1114), .Y(n_1110) );
AOI322xp5_ASAP7_75t_L g1439 ( .A1(n_503), .A2(n_963), .A3(n_1436), .B1(n_1440), .B2(n_1441), .C1(n_1442), .C2(n_1443), .Y(n_1439) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_504), .Y(n_637) );
INVx1_ASAP7_75t_L g1033 ( .A(n_504), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1869 ( .A1(n_504), .A2(n_1358), .B1(n_1870), .B2(n_1871), .Y(n_1869) );
INVx1_ASAP7_75t_L g964 ( .A(n_506), .Y(n_964) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g647 ( .A(n_507), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_507), .B(n_648), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_512), .B1(n_513), .B2(n_516), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_509), .A2(n_513), .B1(n_732), .B2(n_733), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_509), .A2(n_513), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_509), .A2(n_954), .B1(n_955), .B2(n_956), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_509), .A2(n_956), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_509), .A2(n_956), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
AOI22xp33_ASAP7_75t_SL g1816 ( .A1(n_509), .A2(n_518), .B1(n_1817), .B2(n_1818), .Y(n_1816) );
AND2x4_ASAP7_75t_L g513 ( .A(n_510), .B(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g956 ( .A(n_510), .B(n_514), .Y(n_956) );
INVx1_ASAP7_75t_L g1436 ( .A(n_510), .Y(n_1436) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx5_ASAP7_75t_SL g1437 ( .A(n_513), .Y(n_1437) );
AOI22xp33_ASAP7_75t_SL g1819 ( .A1(n_513), .A2(n_520), .B1(n_1804), .B2(n_1820), .Y(n_1819) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_515), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_518), .A2(n_520), .B1(n_687), .B2(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_518), .A2(n_520), .B1(n_947), .B2(n_967), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_518), .A2(n_1055), .B1(n_1056), .B2(n_1057), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_518), .A2(n_1057), .B1(n_1100), .B2(n_1118), .Y(n_1117) );
AOI211xp5_ASAP7_75t_L g1432 ( .A1(n_518), .A2(n_1433), .B(n_1434), .C(n_1438), .Y(n_1432) );
INVx5_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx4_ASAP7_75t_L g1057 ( .A(n_521), .Y(n_1057) );
OAI211xp5_ASAP7_75t_L g1431 ( .A1(n_522), .A2(n_1432), .B(n_1444), .C(n_1454), .Y(n_1431) );
AOI31xp33_ASAP7_75t_L g1811 ( .A1(n_522), .A2(n_1812), .A3(n_1816), .B(n_1819), .Y(n_1811) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g672 ( .A(n_528), .Y(n_672) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_598), .C(n_611), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_557), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_548), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_541), .B2(n_542), .Y(n_533) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_534), .A2(n_553), .B1(n_619), .B2(n_623), .C(n_628), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g1037 ( .A1(n_535), .A2(n_550), .B1(n_601), .B2(n_1026), .C1(n_1029), .C2(n_1038), .Y(n_1037) );
AOI22xp5_ASAP7_75t_L g1887 ( .A1(n_535), .A2(n_542), .B1(n_1862), .B2(n_1864), .Y(n_1887) );
CKINVDCx6p67_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_537), .A2(n_802), .B1(n_889), .B2(n_890), .Y(n_888) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_537), .B(n_538), .Y(n_1188) );
INVx2_ASAP7_75t_L g1419 ( .A(n_537), .Y(n_1419) );
OR2x6_ASAP7_75t_L g543 ( .A(n_538), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g552 ( .A(n_538), .Y(n_552) );
OR2x2_ASAP7_75t_L g866 ( .A(n_538), .B(n_867), .Y(n_866) );
OR2x2_ASAP7_75t_L g869 ( .A(n_538), .B(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g1300 ( .A(n_539), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_539), .B(n_754), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_539), .B(n_580), .Y(n_1330) );
INVx1_ASAP7_75t_L g567 ( .A(n_540), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_542), .A2(n_554), .B1(n_1027), .B2(n_1040), .Y(n_1039) );
CKINVDCx6p67_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g814 ( .A1(n_544), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_814) );
BUFx3_ASAP7_75t_L g882 ( .A(n_544), .Y(n_882) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g812 ( .A(n_545), .Y(n_812) );
BUFx4f_ASAP7_75t_L g1151 ( .A(n_545), .Y(n_1151) );
INVx1_ASAP7_75t_L g1208 ( .A(n_545), .Y(n_1208) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
OR2x2_ASAP7_75t_L g754 ( .A(n_546), .B(n_547), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_553), .B2(n_554), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g1885 ( .A1(n_550), .A2(n_554), .B1(n_601), .B2(n_1861), .C1(n_1867), .C2(n_1886), .Y(n_1885) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g554 ( .A(n_552), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g724 ( .A(n_556), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_556), .A2(n_1470), .B1(n_1471), .B2(n_1472), .Y(n_1469) );
INVx2_ASAP7_75t_SL g1835 ( .A(n_556), .Y(n_1835) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_573), .C(n_593), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_568), .B2(n_569), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_559), .A2(n_568), .B1(n_636), .B2(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g1165 ( .A(n_560), .Y(n_1165) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g829 ( .A(n_561), .Y(n_829) );
NAND2x1p5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g1305 ( .A(n_563), .Y(n_1305) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OR2x6_ASAP7_75t_L g570 ( .A(n_565), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g597 ( .A(n_565), .Y(n_597) );
OR2x2_ASAP7_75t_L g830 ( .A(n_565), .B(n_571), .Y(n_830) );
AND2x4_ASAP7_75t_L g1304 ( .A(n_566), .B(n_1305), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_566), .B(n_572), .Y(n_1307) );
INVx1_ASAP7_75t_L g1323 ( .A(n_566), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_569), .A2(n_796), .B1(n_829), .B2(n_1008), .C(n_1009), .Y(n_1007) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI33xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .A3(n_581), .B1(n_586), .B2(n_589), .B3(n_592), .Y(n_573) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g591 ( .A(n_578), .Y(n_591) );
INVx2_ASAP7_75t_SL g806 ( .A(n_578), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g1880 ( .A1(n_578), .A2(n_1460), .B1(n_1881), .B2(n_1882), .Y(n_1880) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g1298 ( .A(n_579), .Y(n_1298) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g1463 ( .A(n_580), .Y(n_1463) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g743 ( .A(n_584), .Y(n_743) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_585), .Y(n_596) );
BUFx3_ASAP7_75t_L g782 ( .A(n_585), .Y(n_782) );
BUFx4f_ASAP7_75t_L g1000 ( .A(n_585), .Y(n_1000) );
INVx1_ASAP7_75t_L g1077 ( .A(n_585), .Y(n_1077) );
AND2x4_ASAP7_75t_L g1319 ( .A(n_585), .B(n_1300), .Y(n_1319) );
INVx1_ASAP7_75t_L g1528 ( .A(n_585), .Y(n_1528) );
INVx4_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g722 ( .A(n_588), .Y(n_722) );
INVx1_ASAP7_75t_L g1292 ( .A(n_588), .Y(n_1292) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_592), .B(n_721), .C(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g989 ( .A(n_592), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g996 ( .A1(n_592), .A2(n_997), .A3(n_998), .B1(n_999), .B2(n_1001), .B3(n_1005), .Y(n_996) );
AOI33xp33_ASAP7_75t_L g1072 ( .A1(n_592), .A2(n_997), .A3(n_1073), .B1(n_1074), .B2(n_1075), .B3(n_1078), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1130 ( .A(n_592), .B(n_1131), .C(n_1132), .Y(n_1130) );
NAND3xp33_ASAP7_75t_L g1836 ( .A(n_592), .B(n_1837), .C(n_1838), .Y(n_1836) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g1536 ( .A(n_596), .Y(n_1536) );
AND2x2_ASAP7_75t_L g796 ( .A(n_597), .B(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_600), .B(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_600), .B(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_600), .B(n_1141), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_600), .B(n_1197), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_600), .B(n_1261), .Y(n_1260) );
OR2x6_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx2_ASAP7_75t_L g1336 ( .A(n_601), .Y(n_1336) );
NOR2xp67_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g862 ( .A(n_604), .Y(n_862) );
INVx1_ASAP7_75t_L g1495 ( .A(n_605), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_610), .Y(n_605) );
AND2x2_ASAP7_75t_L g636 ( .A(n_606), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g924 ( .A(n_606), .B(n_637), .Y(n_924) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x6_ASAP7_75t_L g639 ( .A(n_607), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g661 ( .A(n_607), .B(n_662), .Y(n_661) );
OR2x6_ASAP7_75t_L g847 ( .A(n_607), .B(n_662), .Y(n_847) );
INVx1_ASAP7_75t_L g1034 ( .A(n_607), .Y(n_1034) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g711 ( .A(n_610), .Y(n_711) );
OAI31xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_641), .A3(n_663), .B(n_668), .Y(n_611) );
INVx8_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g1493 ( .A1(n_614), .A2(n_643), .B1(n_1494), .B2(n_1495), .C1(n_1496), .C2(n_1497), .Y(n_1493) );
AND2x4_ASAP7_75t_L g667 ( .A(n_615), .B(n_626), .Y(n_667) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g643 ( .A(n_617), .B(n_632), .Y(n_643) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g658 ( .A(n_621), .Y(n_658) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_621), .Y(n_840) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g852 ( .A(n_622), .Y(n_852) );
INVx1_ASAP7_75t_L g900 ( .A(n_622), .Y(n_900) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g716 ( .A(n_625), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g1477 ( .A1(n_625), .A2(n_850), .B1(n_1457), .B2(n_1461), .Y(n_1477) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g1028 ( .A1(n_630), .A2(n_1029), .B(n_1030), .C(n_1034), .Y(n_1028) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g1440 ( .A(n_631), .Y(n_1440) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g769 ( .A(n_632), .Y(n_769) );
INVx1_ASAP7_75t_L g915 ( .A(n_633), .Y(n_915) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_636), .A2(n_638), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_636), .A2(n_638), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_636), .A2(n_638), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1511 ( .A1(n_636), .A2(n_638), .B1(n_1512), .B2(n_1513), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_638), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_638), .A2(n_924), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
CKINVDCx11_ASAP7_75t_R g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g1358 ( .A(n_640), .Y(n_1358) );
CKINVDCx6p67_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_643), .A2(n_1016), .B1(n_1018), .B2(n_1021), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B1(n_650), .B2(n_653), .C(n_654), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g1170 ( .A(n_646), .Y(n_1170) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g662 ( .A(n_647), .Y(n_662) );
INVx2_ASAP7_75t_L g761 ( .A(n_647), .Y(n_761) );
INVx3_ASAP7_75t_L g904 ( .A(n_647), .Y(n_904) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_650), .A2(n_654), .B1(n_1147), .B2(n_1148), .C(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_652), .A2(n_654), .B1(n_810), .B2(n_813), .C(n_845), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g1474 ( .A1(n_652), .A2(n_1465), .B1(n_1466), .B2(n_1475), .Y(n_1474) );
OAI22xp33_ASAP7_75t_L g1483 ( .A1(n_652), .A2(n_909), .B1(n_1484), .B2(n_1485), .Y(n_1483) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_654), .A2(n_881), .B1(n_883), .B2(n_904), .C(n_905), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_654), .A2(n_904), .B1(n_1245), .B2(n_1248), .C(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_658), .A2(n_707), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g1854 ( .A1(n_658), .A2(n_921), .B1(n_1855), .B2(n_1856), .Y(n_1854) );
OAI22xp5_ASAP7_75t_L g1860 ( .A1(n_658), .A2(n_707), .B1(n_1861), .B2(n_1862), .Y(n_1860) );
INVx1_ASAP7_75t_L g902 ( .A(n_660), .Y(n_902) );
INVx1_ASAP7_75t_L g1476 ( .A(n_662), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1868 ( .A(n_662), .B(n_1869), .Y(n_1868) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g835 ( .A(n_665), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_665), .A2(n_667), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_665), .A2(n_667), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx3_ASAP7_75t_L g836 ( .A(n_667), .Y(n_836) );
OAI31xp33_ASAP7_75t_L g894 ( .A1(n_668), .A2(n_895), .A3(n_896), .B(n_907), .Y(n_894) );
OAI31xp33_ASAP7_75t_L g1262 ( .A1(n_668), .A2(n_1263), .A3(n_1264), .B(n_1272), .Y(n_1262) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
CKINVDCx8_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
AOI221x1_ASAP7_75t_SL g1491 ( .A1(n_670), .A2(n_951), .B1(n_1492), .B2(n_1520), .C(n_1530), .Y(n_1491) );
XNOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_930), .Y(n_673) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_790), .Y(n_674) );
XNOR2x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_737), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_685), .C(n_688), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_702), .C(n_713), .D(n_720), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_698), .C(n_699), .Y(n_692) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g980 ( .A(n_699), .B(n_981), .C(n_982), .Y(n_980) );
NAND3xp33_ASAP7_75t_L g1127 ( .A(n_699), .B(n_1128), .C(n_1129), .Y(n_1127) );
NAND3xp33_ASAP7_75t_L g1832 ( .A(n_699), .B(n_1833), .C(n_1834), .Y(n_1832) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_710), .C(n_712), .Y(n_702) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g1067 ( .A(n_707), .Y(n_1067) );
INVx1_ASAP7_75t_L g1267 ( .A(n_707), .Y(n_1267) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g843 ( .A(n_708), .Y(n_843) );
INVx2_ASAP7_75t_L g921 ( .A(n_708), .Y(n_921) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_709), .Y(n_856) );
INVx3_ASAP7_75t_L g978 ( .A(n_709), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g971 ( .A(n_712), .B(n_972), .C(n_973), .Y(n_971) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_712), .B(n_1124), .C(n_1126), .Y(n_1123) );
CKINVDCx8_ASAP7_75t_R g1378 ( .A(n_712), .Y(n_1378) );
INVx1_ASAP7_75t_L g1180 ( .A(n_716), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g771 ( .A(n_719), .Y(n_771) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_719), .Y(n_1071) );
AOI31xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_731), .A3(n_734), .B(n_736), .Y(n_725) );
INVx1_ASAP7_75t_L g961 ( .A(n_729), .Y(n_961) );
AO21x1_ASAP7_75t_SL g757 ( .A1(n_736), .A2(n_758), .B(n_763), .Y(n_757) );
CKINVDCx16_ASAP7_75t_R g969 ( .A(n_736), .Y(n_969) );
AND4x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_757), .C(n_766), .D(n_775), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g789 ( .A(n_739), .B(n_757), .C(n_766), .D(n_775), .Y(n_789) );
OAI31xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_748), .A3(n_751), .B(n_756), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .C(n_747), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g1451 ( .A(n_753), .Y(n_1451) );
BUFx2_ASAP7_75t_L g809 ( .A(n_754), .Y(n_809) );
INVx1_ASAP7_75t_L g816 ( .A(n_754), .Y(n_816) );
INVx2_ASAP7_75t_L g868 ( .A(n_754), .Y(n_868) );
INVx1_ASAP7_75t_SL g1091 ( .A(n_756), .Y(n_1091) );
OAI31xp33_ASAP7_75t_SL g1444 ( .A1(n_756), .A2(n_1445), .A3(n_1446), .B(n_1447), .Y(n_1444) );
AOI211xp5_ASAP7_75t_L g1800 ( .A1(n_756), .A2(n_1801), .B(n_1811), .C(n_1821), .Y(n_1800) );
OAI22xp33_ASAP7_75t_L g1408 ( .A1(n_761), .A2(n_912), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
OAI21xp5_ASAP7_75t_SL g1516 ( .A1(n_761), .A2(n_1517), .B(n_1518), .Y(n_1516) );
OAI21xp33_ASAP7_75t_L g1863 ( .A1(n_761), .A2(n_1864), .B(n_1865), .Y(n_1863) );
NAND3xp33_ASAP7_75t_L g974 ( .A(n_767), .B(n_975), .C(n_979), .Y(n_974) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_767), .B(n_1121), .C(n_1122), .Y(n_1120) );
A2O1A1Ixp33_ASAP7_75t_L g1866 ( .A1(n_769), .A2(n_1034), .B(n_1867), .C(n_1868), .Y(n_1866) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_778), .A2(n_1253), .B1(n_1254), .B2(n_1255), .Y(n_1252) );
INVx1_ASAP7_75t_L g1296 ( .A(n_778), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1878 ( .A1(n_778), .A2(n_780), .B1(n_1855), .B2(n_1856), .Y(n_1878) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g787 ( .A(n_780), .Y(n_787) );
INVx1_ASAP7_75t_L g824 ( .A(n_780), .Y(n_824) );
INVx1_ASAP7_75t_L g1533 ( .A(n_787), .Y(n_1533) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B1(n_871), .B2(n_929), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AND4x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_831), .C(n_833), .D(n_863), .Y(n_793) );
NOR3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_799), .C(n_827), .Y(n_794) );
NOR3xp33_ASAP7_75t_SL g873 ( .A(n_795), .B(n_874), .C(n_891), .Y(n_873) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_796), .Y(n_1143) );
NOR3xp33_ASAP7_75t_SL g1198 ( .A(n_796), .B(n_1199), .C(n_1211), .Y(n_1198) );
NOR3xp33_ASAP7_75t_SL g1238 ( .A(n_796), .B(n_1239), .C(n_1256), .Y(n_1238) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1291 ( .A(n_798), .Y(n_1291) );
OAI33xp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .A3(n_808), .B1(n_814), .B2(n_819), .B3(n_826), .Y(n_799) );
OAI33xp33_ASAP7_75t_L g874 ( .A1(n_800), .A2(n_826), .A3(n_875), .B1(n_880), .B2(n_884), .B3(n_888), .Y(n_874) );
INVx1_ASAP7_75t_SL g997 ( .A(n_800), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_800), .A2(n_1153), .B1(n_1200), .B2(n_1205), .Y(n_1199) );
OAI33xp33_ASAP7_75t_L g1239 ( .A1(n_800), .A2(n_826), .A3(n_1240), .B1(n_1244), .B2(n_1249), .B3(n_1252), .Y(n_1239) );
OAI33xp33_ASAP7_75t_L g1455 ( .A1(n_800), .A2(n_826), .A3(n_1456), .B1(n_1464), .B2(n_1467), .B3(n_1469), .Y(n_1455) );
OAI22xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_804), .B1(n_805), .B2(n_807), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
BUFx3_ASAP7_75t_L g1161 ( .A(n_803), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_804), .A2(n_807), .B1(n_839), .B2(n_841), .Y(n_838) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_811), .B2(n_813), .Y(n_808) );
OAI22xp33_ASAP7_75t_L g880 ( .A1(n_809), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g1200 ( .A1(n_809), .A2(n_1158), .B1(n_1201), .B2(n_1202), .C(n_1203), .Y(n_1200) );
OAI221xp5_ASAP7_75t_L g1205 ( .A1(n_809), .A2(n_1206), .B1(n_1207), .B2(n_1209), .C(n_1210), .Y(n_1205) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g944 ( .A(n_812), .Y(n_944) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_815), .Y(n_1146) );
OAI221xp5_ASAP7_75t_L g1537 ( .A1(n_815), .A2(n_1246), .B1(n_1496), .B2(n_1497), .C(n_1538), .Y(n_1537) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_822), .B1(n_823), .B2(n_825), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g876 ( .A(n_821), .Y(n_876) );
BUFx2_ASAP7_75t_L g1310 ( .A(n_821), .Y(n_1310) );
BUFx3_ASAP7_75t_L g1423 ( .A(n_821), .Y(n_1423) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI31xp33_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_837), .A3(n_848), .B(n_862), .Y(n_833) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g910 ( .A(n_845), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_845), .B(n_1031), .Y(n_1030) );
BUFx3_ASAP7_75t_L g1220 ( .A(n_845), .Y(n_1220) );
BUFx3_ASAP7_75t_L g1401 ( .A(n_845), .Y(n_1401) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g1519 ( .A(n_847), .Y(n_1519) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_853), .B1(n_854), .B2(n_857), .C(n_858), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_852), .B(n_1436), .Y(n_1435) );
BUFx2_ASAP7_75t_L g1507 ( .A(n_852), .Y(n_1507) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g1125 ( .A(n_856), .Y(n_1125) );
INVx2_ASAP7_75t_SL g1481 ( .A(n_856), .Y(n_1481) );
OAI31xp33_ASAP7_75t_L g1166 ( .A1(n_862), .A2(n_1167), .A3(n_1168), .B(n_1174), .Y(n_1166) );
INVx1_ASAP7_75t_L g1412 ( .A(n_862), .Y(n_1412) );
OAI31xp33_ASAP7_75t_L g1852 ( .A1(n_862), .A2(n_1853), .A3(n_1872), .B(n_1873), .Y(n_1852) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g885 ( .A(n_868), .Y(n_885) );
INVx2_ASAP7_75t_L g1156 ( .A(n_868), .Y(n_1156) );
INVx1_ASAP7_75t_L g929 ( .A(n_871), .Y(n_929) );
AND4x1_ASAP7_75t_L g872 ( .A(n_873), .B(n_892), .C(n_894), .D(n_926), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_877), .B1(n_878), .B2(n_879), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_876), .A2(n_1241), .B1(n_1242), .B2(n_1243), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_877), .A2(n_879), .B1(n_898), .B2(n_901), .Y(n_897) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_882), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_884) );
OAI22xp33_ASAP7_75t_L g1467 ( .A1(n_882), .A2(n_885), .B1(n_1433), .B2(n_1468), .Y(n_1467) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_885), .A2(n_1245), .B1(n_1246), .B2(n_1248), .Y(n_1244) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_885), .A2(n_1158), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
OAI22xp33_ASAP7_75t_SL g1464 ( .A1(n_885), .A2(n_1207), .B1(n_1465), .B2(n_1466), .Y(n_1464) );
OAI22xp5_ASAP7_75t_SL g916 ( .A1(n_898), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_898), .A2(n_1216), .B1(n_1217), .B2(n_1218), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1265 ( .A1(n_898), .A2(n_1241), .B1(n_1243), .B2(n_1266), .Y(n_1265) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g1225 ( .A(n_899), .Y(n_1225) );
INVx2_ASAP7_75t_L g1274 ( .A(n_899), .Y(n_1274) );
INVx2_ASAP7_75t_SL g1479 ( .A(n_899), .Y(n_1479) );
BUFx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g1178 ( .A(n_900), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_901), .A2(n_1370), .B1(n_1403), .B2(n_1404), .Y(n_1402) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OAI21xp5_ASAP7_75t_L g1857 ( .A1(n_904), .A2(n_1858), .B(n_1859), .Y(n_1857) );
BUFx2_ASAP7_75t_L g1377 ( .A(n_905), .Y(n_1377) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_911), .B1(n_912), .B2(n_914), .C(n_915), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g1367 ( .A(n_910), .Y(n_1367) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_912), .A2(n_1366), .B1(n_1367), .B2(n_1368), .Y(n_1365) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g1398 ( .A(n_913), .Y(n_1398) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g1069 ( .A(n_921), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
OAI22x1_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B1(n_991), .B2(n_992), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g990 ( .A(n_936), .Y(n_990) );
AOI221x1_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_951), .B1(n_952), .B2(n_969), .C(n_970), .Y(n_936) );
NAND3xp33_ASAP7_75t_L g937 ( .A(n_938), .B(n_945), .C(n_948), .Y(n_937) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g1103 ( .A(n_941), .Y(n_1103) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
AOI221x1_ASAP7_75t_L g1094 ( .A1(n_951), .A2(n_969), .B1(n_1095), .B2(n_1106), .C(n_1119), .Y(n_1094) );
NAND4xp25_ASAP7_75t_SL g952 ( .A(n_953), .B(n_957), .C(n_966), .D(n_968), .Y(n_952) );
AOI222xp33_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_959), .B1(n_960), .B2(n_961), .C1(n_962), .C2(n_963), .Y(n_957) );
AOI222xp33_ASAP7_75t_L g1058 ( .A1(n_959), .A2(n_961), .B1(n_963), .B2(n_1059), .C1(n_1060), .C2(n_1061), .Y(n_1058) );
AND2x4_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_964), .A2(n_1008), .B1(n_1009), .B2(n_1032), .Y(n_1031) );
NAND4xp25_ASAP7_75t_SL g1050 ( .A(n_968), .B(n_1051), .C(n_1054), .D(n_1058), .Y(n_1050) );
NAND4xp25_ASAP7_75t_SL g1106 ( .A(n_968), .B(n_1107), .C(n_1110), .D(n_1117), .Y(n_1106) );
AOI211xp5_ASAP7_75t_L g1049 ( .A1(n_969), .A2(n_1050), .B(n_1062), .C(n_1080), .Y(n_1049) );
NAND4xp25_ASAP7_75t_L g970 ( .A(n_971), .B(n_974), .C(n_980), .D(n_983), .Y(n_970) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AND2x4_ASAP7_75t_L g1342 ( .A(n_978), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1509 ( .A(n_978), .Y(n_1509) );
NAND3xp33_ASAP7_75t_L g983 ( .A(n_984), .B(n_986), .C(n_988), .Y(n_983) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_SL g991 ( .A(n_992), .Y(n_991) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NAND4xp75_ASAP7_75t_L g994 ( .A(n_995), .B(n_1010), .C(n_1037), .D(n_1039), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_996), .B(n_1007), .Y(n_995) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
OAI21xp5_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1022), .B(n_1035), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1015), .Y(n_1011) );
AND2x6_ASAP7_75t_L g1345 ( .A(n_1019), .B(n_1343), .Y(n_1345) );
NAND2x1p5_ASAP7_75t_L g1360 ( .A(n_1019), .B(n_1355), .Y(n_1360) );
BUFx2_ASAP7_75t_L g1814 ( .A(n_1019), .Y(n_1814) );
NAND2x1_ASAP7_75t_SL g1354 ( .A(n_1032), .B(n_1355), .Y(n_1354) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
OAI31xp33_ASAP7_75t_L g1212 ( .A1(n_1035), .A2(n_1213), .A3(n_1214), .B(n_1223), .Y(n_1212) );
BUFx8_ASAP7_75t_SL g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1036), .Y(n_1287) );
XNOR2xp5_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1191), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B1(n_1136), .B2(n_1190), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
OA22x2_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1092), .B1(n_1093), .B2(n_1135), .Y(n_1046) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1047), .Y(n_1135) );
XNOR2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1049), .Y(n_1047) );
NAND2xp5_ASAP7_75t_SL g1062 ( .A(n_1063), .B(n_1072), .Y(n_1062) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
AOI31xp33_ASAP7_75t_SL g1080 ( .A1(n_1081), .A2(n_1085), .A3(n_1088), .B(n_1091), .Y(n_1080) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1083), .Y(n_1448) );
AOI21xp5_ASAP7_75t_L g1805 ( .A1(n_1083), .A2(n_1806), .B(n_1807), .Y(n_1805) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1094), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1099), .Y(n_1095) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
NAND4xp25_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1123), .C(n_1127), .D(n_1130), .Y(n_1119) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1125), .Y(n_1217) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1136), .Y(n_1190) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
XNOR2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1139), .Y(n_1137) );
AND4x1_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1142), .C(n_1166), .D(n_1186), .Y(n_1139) );
NOR3xp33_ASAP7_75t_SL g1142 ( .A(n_1143), .B(n_1144), .C(n_1164), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1147), .B1(n_1148), .B2(n_1149), .C(n_1152), .Y(n_1145) );
OAI221xp5_ASAP7_75t_L g1531 ( .A1(n_1146), .A2(n_1510), .B1(n_1532), .B2(n_1533), .C(n_1534), .Y(n_1531) );
BUFx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1151), .Y(n_1158) );
CKINVDCx5p33_ASAP7_75t_R g1153 ( .A(n_1154), .Y(n_1153) );
OAI221xp5_ASAP7_75t_L g1155 ( .A1(n_1156), .A2(n_1157), .B1(n_1158), .B2(n_1159), .C(n_1160), .Y(n_1155) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
OAI221xp5_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1179), .B1(n_1180), .B2(n_1181), .C(n_1182), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1189), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_1192), .A2(n_1193), .B1(n_1282), .B2(n_1379), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
AO22x2_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1235), .B1(n_1236), .B2(n_1281), .Y(n_1193) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1194), .Y(n_1281) );
AND4x1_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1198), .C(n_1212), .D(n_1232), .Y(n_1195) );
OAI21xp33_ASAP7_75t_L g1219 ( .A1(n_1202), .A2(n_1220), .B(n_1221), .Y(n_1219) );
INVx2_ASAP7_75t_SL g1254 ( .A(n_1204), .Y(n_1254) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1208), .Y(n_1247) );
OAI22xp33_ASAP7_75t_L g1376 ( .A1(n_1220), .A2(n_1320), .B1(n_1325), .B2(n_1377), .Y(n_1376) );
AND2x4_ASAP7_75t_L g1348 ( .A(n_1222), .B(n_1343), .Y(n_1348) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1225), .Y(n_1371) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
AND4x1_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1257), .C(n_1260), .D(n_1262), .Y(n_1237) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1259), .Y(n_1257) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_1270), .Y(n_1269) );
INVx2_ASAP7_75t_SL g1270 ( .A(n_1271), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1283), .Y(n_1379) );
XNOR2x1_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1285), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1337), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1288), .B1(n_1331), .B2(n_1332), .Y(n_1286) );
NAND3xp33_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1308), .C(n_1324), .Y(n_1288) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1295), .B1(n_1299), .B2(n_1301), .C(n_1302), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
AOI221xp5_ASAP7_75t_L g1414 ( .A1(n_1299), .A2(n_1406), .B1(n_1415), .B2(n_1417), .C(n_1420), .Y(n_1414) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx2_ASAP7_75t_SL g1306 ( .A(n_1307), .Y(n_1306) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1316), .B1(n_1318), .B2(n_1320), .C(n_1321), .Y(n_1308) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
AOI221xp5_ASAP7_75t_L g1421 ( .A1(n_1318), .A2(n_1321), .B1(n_1410), .B2(n_1422), .C(n_1424), .Y(n_1421) );
BUFx6f_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_SL g1322 ( .A(n_1323), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1326), .B1(n_1328), .B2(n_1329), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_1326), .A2(n_1329), .B1(n_1407), .B2(n_1409), .Y(n_1425) );
INVx6_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx4_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_1332), .A2(n_1412), .B1(n_1413), .B2(n_1426), .Y(n_1411) );
INVx5_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
AND2x4_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1336), .Y(n_1333) );
INVx3_ASAP7_75t_L g1355 ( .A(n_1335), .Y(n_1355) );
NOR3xp33_ASAP7_75t_SL g1337 ( .A(n_1338), .B(n_1351), .C(n_1361), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1346), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_1340), .A2(n_1341), .B1(n_1344), .B2(n_1345), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_1341), .A2(n_1345), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
BUFx2_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_1347), .A2(n_1348), .B1(n_1349), .B2(n_1350), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_1348), .A2(n_1350), .B1(n_1392), .B2(n_1393), .Y(n_1391) );
INVx2_ASAP7_75t_SL g1352 ( .A(n_1353), .Y(n_1352) );
INVx2_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
NAND2x1p5_ASAP7_75t_L g1357 ( .A(n_1355), .B(n_1358), .Y(n_1357) );
BUFx4f_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
BUFx2_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
OAI33xp33_ASAP7_75t_L g1361 ( .A1(n_1362), .A2(n_1365), .A3(n_1369), .B1(n_1375), .B2(n_1376), .B3(n_1378), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
OAI33xp33_ASAP7_75t_L g1395 ( .A1(n_1364), .A2(n_1378), .A3(n_1396), .B1(n_1402), .B2(n_1405), .B3(n_1408), .Y(n_1395) );
OAI33xp33_ASAP7_75t_L g1473 ( .A1(n_1364), .A2(n_1474), .A3(n_1477), .B1(n_1478), .B2(n_1483), .B3(n_1486), .Y(n_1473) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_1370), .A2(n_1372), .B1(n_1373), .B2(n_1374), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_1370), .A2(n_1373), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
INVx2_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_1382), .A2(n_1427), .B1(n_1541), .B2(n_1542), .Y(n_1381) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1382), .Y(n_1541) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1411), .Y(n_1385) );
NOR3xp33_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1394), .C(n_1395), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .Y(n_1387) );
OAI22xp33_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1398), .B1(n_1399), .B2(n_1400), .Y(n_1396) );
BUFx3_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
OAI21xp5_ASAP7_75t_L g1503 ( .A1(n_1401), .A2(n_1504), .B(n_1505), .Y(n_1503) );
NAND3xp33_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1421), .C(n_1425), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVxp67_ASAP7_75t_SL g1542 ( .A(n_1427), .Y(n_1542) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1429), .B1(n_1489), .B2(n_1490), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
HB1xp67_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1431), .Y(n_1487) );
INVx2_ASAP7_75t_L g1460 ( .A(n_1450), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g1478 ( .A1(n_1452), .A2(n_1479), .B1(n_1480), .B2(n_1482), .Y(n_1478) );
NOR2xp33_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1473), .Y(n_1454) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_1457), .A2(n_1458), .B1(n_1461), .B2(n_1462), .Y(n_1456) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1460), .Y(n_1535) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx2_ASAP7_75t_SL g1489 ( .A(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1491), .Y(n_1540) );
NAND3xp33_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1498), .C(n_1501), .Y(n_1492) );
NOR3xp33_ASAP7_75t_L g1501 ( .A(n_1502), .B(n_1514), .C(n_1519), .Y(n_1501) );
OAI21xp5_ASAP7_75t_SL g1502 ( .A1(n_1503), .A2(n_1506), .B(n_1511), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g1506 ( .A1(n_1507), .A2(n_1508), .B1(n_1509), .B2(n_1510), .Y(n_1506) );
NAND4xp25_ASAP7_75t_SL g1520 ( .A(n_1521), .B(n_1524), .C(n_1526), .D(n_1529), .Y(n_1520) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
OAI221xp5_ASAP7_75t_SL g1543 ( .A1(n_1544), .A2(n_1794), .B1(n_1796), .B2(n_1839), .C(n_1843), .Y(n_1543) );
AND4x1_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1760), .C(n_1779), .D(n_1784), .Y(n_1544) );
AOI211xp5_ASAP7_75t_L g1545 ( .A1(n_1546), .A2(n_1574), .B(n_1707), .C(n_1744), .Y(n_1545) );
OAI221xp5_ASAP7_75t_L g1707 ( .A1(n_1546), .A2(n_1708), .B1(n_1723), .B2(n_1739), .C(n_1893), .Y(n_1707) );
INVx3_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
O2A1O1Ixp33_ASAP7_75t_L g1760 ( .A1(n_1547), .A2(n_1761), .B(n_1766), .C(n_1770), .Y(n_1760) );
INVx2_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1750 ( .A(n_1549), .B(n_1607), .Y(n_1750) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
NOR2xp33_ASAP7_75t_L g1755 ( .A(n_1550), .B(n_1717), .Y(n_1755) );
NOR3xp33_ASAP7_75t_L g1778 ( .A(n_1550), .B(n_1631), .C(n_1656), .Y(n_1778) );
BUFx3_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1552), .Y(n_1610) );
AND2x4_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1556), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1553), .B(n_1556), .Y(n_1587) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
AND2x4_ASAP7_75t_L g1560 ( .A(n_1554), .B(n_1556), .Y(n_1560) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1555), .B(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1557), .Y(n_1568) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx2_ASAP7_75t_L g1592 ( .A(n_1559), .Y(n_1592) );
OAI22xp5_ASAP7_75t_SL g1609 ( .A1(n_1559), .A2(n_1610), .B1(n_1611), .B2(n_1612), .Y(n_1609) );
INVx2_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
OAI22xp33_ASAP7_75t_L g1561 ( .A1(n_1562), .A2(n_1563), .B1(n_1569), .B2(n_1570), .Y(n_1561) );
BUFx3_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
OAI22xp33_ASAP7_75t_L g1593 ( .A1(n_1564), .A2(n_1594), .B1(n_1595), .B2(n_1596), .Y(n_1593) );
BUFx6f_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
OR2x2_ASAP7_75t_L g1565 ( .A(n_1566), .B(n_1567), .Y(n_1565) );
OR2x2_ASAP7_75t_L g1572 ( .A(n_1566), .B(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1566), .Y(n_1583) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1567), .Y(n_1582) );
HB1xp67_ASAP7_75t_L g1795 ( .A(n_1570), .Y(n_1795) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
HB1xp67_ASAP7_75t_L g1596 ( .A(n_1572), .Y(n_1596) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1573), .Y(n_1585) );
NAND5xp2_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1627), .C(n_1667), .D(n_1680), .E(n_1696), .Y(n_1574) );
AOI21xp5_ASAP7_75t_L g1575 ( .A1(n_1576), .A2(n_1605), .B(n_1617), .Y(n_1575) );
INVx2_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1588), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1578), .B(n_1623), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1578), .B(n_1638), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1578), .B(n_1625), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1578), .B(n_1591), .Y(n_1689) );
OR2x2_ASAP7_75t_L g1710 ( .A(n_1578), .B(n_1711), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1578), .B(n_1640), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1578), .B(n_1733), .Y(n_1776) );
CKINVDCx5p33_ASAP7_75t_R g1578 ( .A(n_1579), .Y(n_1578) );
HB1xp67_ASAP7_75t_L g1642 ( .A(n_1579), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1579), .B(n_1590), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1579), .B(n_1659), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1579), .B(n_1640), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1579), .B(n_1638), .Y(n_1679) );
OR2x2_ASAP7_75t_L g1698 ( .A(n_1579), .B(n_1699), .Y(n_1698) );
OR2x2_ASAP7_75t_L g1720 ( .A(n_1579), .B(n_1659), .Y(n_1720) );
NOR2xp33_ASAP7_75t_L g1726 ( .A(n_1579), .B(n_1727), .Y(n_1726) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1579), .B(n_1598), .Y(n_1730) );
NOR2xp33_ASAP7_75t_L g1738 ( .A(n_1579), .B(n_1656), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1579), .B(n_1656), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1579), .B(n_1625), .Y(n_1769) );
AND2x4_ASAP7_75t_SL g1579 ( .A(n_1580), .B(n_1586), .Y(n_1579) );
AND2x4_ASAP7_75t_L g1581 ( .A(n_1582), .B(n_1583), .Y(n_1581) );
AND2x4_ASAP7_75t_L g1584 ( .A(n_1583), .B(n_1585), .Y(n_1584) );
HB1xp67_ASAP7_75t_L g1890 ( .A(n_1585), .Y(n_1890) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1597), .Y(n_1588) );
NOR2xp33_ASAP7_75t_L g1623 ( .A(n_1589), .B(n_1624), .Y(n_1623) );
INVxp67_ASAP7_75t_L g1655 ( .A(n_1589), .Y(n_1655) );
HB1xp67_ASAP7_75t_L g1670 ( .A(n_1589), .Y(n_1670) );
NOR2x1p5_ASAP7_75t_L g1733 ( .A(n_1589), .B(n_1734), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1589), .B(n_1738), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1746 ( .A(n_1589), .B(n_1662), .Y(n_1746) );
INVx2_ASAP7_75t_SL g1589 ( .A(n_1590), .Y(n_1589) );
BUFx3_ASAP7_75t_L g1631 ( .A(n_1590), .Y(n_1631) );
BUFx2_ASAP7_75t_L g1675 ( .A(n_1590), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1719 ( .A(n_1590), .B(n_1619), .Y(n_1719) );
NOR2xp33_ASAP7_75t_L g1731 ( .A(n_1590), .B(n_1663), .Y(n_1731) );
INVx2_ASAP7_75t_SL g1590 ( .A(n_1591), .Y(n_1590) );
INVx2_ASAP7_75t_L g1734 ( .A(n_1597), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1597), .B(n_1650), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1601), .Y(n_1597) );
INVxp67_ASAP7_75t_SL g1626 ( .A(n_1598), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1598), .B(n_1602), .Y(n_1638) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1598), .Y(n_1641) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1598), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1600), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1601), .B(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1601), .Y(n_1656) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1602), .B(n_1626), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1604), .Y(n_1602) );
AOI221xp5_ASAP7_75t_L g1723 ( .A1(n_1605), .A2(n_1724), .B1(n_1732), .B2(n_1733), .C(n_1735), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1613), .Y(n_1605) );
NAND2xp5_ASAP7_75t_SL g1683 ( .A(n_1606), .B(n_1662), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1606), .B(n_1663), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1606), .B(n_1676), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1606), .B(n_1619), .Y(n_1774) );
O2A1O1Ixp33_ASAP7_75t_L g1792 ( .A1(n_1606), .A2(n_1664), .B(n_1720), .C(n_1793), .Y(n_1792) );
CKINVDCx6p67_ASAP7_75t_R g1606 ( .A(n_1607), .Y(n_1606) );
OR2x2_ASAP7_75t_L g1644 ( .A(n_1607), .B(n_1613), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1607), .B(n_1655), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1607), .B(n_1662), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1607), .B(n_1647), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1607), .B(n_1613), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1607), .B(n_1614), .Y(n_1702) );
CKINVDCx5p33_ASAP7_75t_R g1732 ( .A(n_1607), .Y(n_1732) );
OR2x2_ASAP7_75t_L g1759 ( .A(n_1607), .B(n_1633), .Y(n_1759) );
OR2x6_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
OR2x2_ASAP7_75t_L g1765 ( .A(n_1608), .B(n_1609), .Y(n_1765) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1613), .Y(n_1717) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1614), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1614), .B(n_1619), .Y(n_1653) );
BUFx6f_ASAP7_75t_L g1672 ( .A(n_1614), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1614), .B(n_1663), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1622), .Y(n_1617) );
NAND2xp67_ASAP7_75t_L g1786 ( .A(n_1618), .B(n_1649), .Y(n_1786) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1633 ( .A(n_1619), .B(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1619), .Y(n_1648) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1619), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1622), .Y(n_1789) );
OR2x2_ASAP7_75t_L g1711 ( .A(n_1624), .B(n_1675), .Y(n_1711) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1625), .B(n_1650), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1625), .B(n_1689), .Y(n_1703) );
AOI321xp33_ASAP7_75t_L g1627 ( .A1(n_1628), .A2(n_1635), .A3(n_1642), .B1(n_1643), .B2(n_1645), .C(n_1651), .Y(n_1627) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1628), .Y(n_1793) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1632), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_1630), .B(n_1640), .Y(n_1791) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1631), .B(n_1658), .Y(n_1657) );
A2O1A1Ixp33_ASAP7_75t_L g1712 ( .A1(n_1631), .A2(n_1713), .B(n_1714), .C(n_1716), .Y(n_1712) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1631), .B(n_1662), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1631), .B(n_1715), .Y(n_1772) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
INVx2_ASAP7_75t_L g1666 ( .A(n_1633), .Y(n_1666) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1633), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1634), .B(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1639), .Y(n_1636) );
OR2x2_ASAP7_75t_L g1687 ( .A(n_1637), .B(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1638), .B(n_1706), .Y(n_1705) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1640), .B(n_1650), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1643), .B(n_1737), .Y(n_1736) );
AOI222xp33_ASAP7_75t_L g1739 ( .A1(n_1643), .A2(n_1653), .B1(n_1740), .B2(n_1741), .C1(n_1742), .C2(n_1743), .Y(n_1739) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVxp67_ASAP7_75t_SL g1645 ( .A(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1649), .Y(n_1646) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1647), .Y(n_1749) );
INVx3_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1648), .B(n_1702), .Y(n_1701) );
OAI21xp33_ASAP7_75t_L g1724 ( .A1(n_1648), .A2(n_1725), .B(n_1728), .Y(n_1724) );
AOI32xp33_ASAP7_75t_L g1747 ( .A1(n_1648), .A2(n_1685), .A3(n_1711), .B1(n_1714), .B2(n_1748), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1648), .B(n_1772), .Y(n_1783) );
OAI321xp33_ASAP7_75t_L g1651 ( .A1(n_1652), .A2(n_1654), .A3(n_1656), .B1(n_1657), .B2(n_1660), .C(n_1664), .Y(n_1651) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
AOI221xp5_ASAP7_75t_SL g1696 ( .A1(n_1653), .A2(n_1697), .B1(n_1700), .B2(n_1703), .C(n_1704), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1653), .B(n_1665), .Y(n_1722) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1656), .Y(n_1659) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1666), .Y(n_1664) );
AOI21xp5_ASAP7_75t_L g1667 ( .A1(n_1668), .A2(n_1672), .B(n_1673), .Y(n_1667) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1671), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_1671), .B(n_1782), .Y(n_1781) );
AOI211xp5_ASAP7_75t_L g1708 ( .A1(n_1672), .A2(n_1709), .B(n_1712), .C(n_1721), .Y(n_1708) );
CKINVDCx14_ASAP7_75t_R g1787 ( .A(n_1672), .Y(n_1787) );
AOI21xp5_ASAP7_75t_L g1673 ( .A1(n_1674), .A2(n_1677), .B(n_1678), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1676), .Y(n_1674) );
INVx2_ASAP7_75t_L g1695 ( .A(n_1675), .Y(n_1695) );
NOR2xp33_ASAP7_75t_L g1697 ( .A(n_1675), .B(n_1698), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1725 ( .A(n_1675), .B(n_1726), .Y(n_1725) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1676), .Y(n_1713) );
OAI21xp33_ASAP7_75t_L g1757 ( .A1(n_1676), .A2(n_1709), .B(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1677), .Y(n_1743) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1679), .B(n_1695), .Y(n_1694) );
NOR2xp33_ASAP7_75t_L g1754 ( .A(n_1679), .B(n_1715), .Y(n_1754) );
AOI221xp5_ASAP7_75t_L g1680 ( .A1(n_1681), .A2(n_1682), .B1(n_1684), .B2(n_1690), .C(n_1691), .Y(n_1680) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
NAND2xp5_ASAP7_75t_SL g1684 ( .A(n_1685), .B(n_1687), .Y(n_1684) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVxp67_ASAP7_75t_SL g1742 ( .A(n_1687), .Y(n_1742) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1690), .Y(n_1767) );
INVxp67_ASAP7_75t_SL g1691 ( .A(n_1692), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1694), .Y(n_1692) );
OAI221xp5_ASAP7_75t_L g1744 ( .A1(n_1695), .A2(n_1745), .B1(n_1750), .B2(n_1751), .C(n_1757), .Y(n_1744) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1699), .Y(n_1727) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
OAI31xp33_ASAP7_75t_L g1779 ( .A1(n_1702), .A2(n_1709), .A3(n_1780), .B(n_1783), .Y(n_1779) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
AOI221xp5_ASAP7_75t_L g1784 ( .A1(n_1706), .A2(n_1785), .B1(n_1787), .B2(n_1788), .C(n_1792), .Y(n_1784) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
OAI21xp33_ASAP7_75t_L g1777 ( .A1(n_1715), .A2(n_1758), .B(n_1778), .Y(n_1777) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1718), .Y(n_1716) );
NOR2xp33_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1720), .Y(n_1718) );
INVxp67_ASAP7_75t_SL g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1727), .Y(n_1762) );
INVxp67_ASAP7_75t_SL g1741 ( .A(n_1728), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1731), .Y(n_1728) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
AOI21xp33_ASAP7_75t_SL g1745 ( .A1(n_1730), .A2(n_1746), .B(n_1747), .Y(n_1745) );
INVxp67_ASAP7_75t_SL g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1740), .Y(n_1764) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1749), .Y(n_1782) );
AOI22xp33_ASAP7_75t_L g1751 ( .A1(n_1752), .A2(n_1753), .B1(n_1755), .B2(n_1756), .Y(n_1751) );
INVxp33_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
O2A1O1Ixp33_ASAP7_75t_SL g1761 ( .A1(n_1762), .A2(n_1763), .B(n_1764), .C(n_1765), .Y(n_1761) );
NOR2xp33_ASAP7_75t_L g1766 ( .A(n_1767), .B(n_1768), .Y(n_1766) );
OAI221xp5_ASAP7_75t_L g1770 ( .A1(n_1767), .A2(n_1771), .B1(n_1773), .B2(n_1775), .C(n_1777), .Y(n_1770) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
CKINVDCx5p33_ASAP7_75t_R g1773 ( .A(n_1774), .Y(n_1773) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
NAND2xp5_ASAP7_75t_L g1788 ( .A(n_1789), .B(n_1790), .Y(n_1788) );
INVxp67_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
BUFx2_ASAP7_75t_SL g1794 ( .A(n_1795), .Y(n_1794) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
HB1xp67_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
XNOR2xp5_ASAP7_75t_L g1798 ( .A(n_1799), .B(n_1800), .Y(n_1798) );
NAND4xp25_ASAP7_75t_L g1821 ( .A(n_1822), .B(n_1827), .C(n_1832), .D(n_1836), .Y(n_1821) );
INVx2_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
NAND3xp33_ASAP7_75t_L g1827 ( .A(n_1828), .B(n_1830), .C(n_1831), .Y(n_1827) );
INVx2_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx2_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
CKINVDCx5p33_ASAP7_75t_R g1845 ( .A(n_1846), .Y(n_1845) );
OAI21xp5_ASAP7_75t_L g1889 ( .A1(n_1847), .A2(n_1890), .B(n_1891), .Y(n_1889) );
INVxp33_ASAP7_75t_SL g1848 ( .A(n_1849), .Y(n_1848) );
HB1xp67_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
NAND4xp25_ASAP7_75t_L g1851 ( .A(n_1852), .B(n_1874), .C(n_1885), .D(n_1887), .Y(n_1851) );
OAI221xp5_ASAP7_75t_L g1853 ( .A1(n_1854), .A2(n_1857), .B1(n_1860), .B2(n_1863), .C(n_1866), .Y(n_1853) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
BUFx2_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
endmodule