module real_jpeg_16174_n_15 (n_108, n_8, n_116, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_6, n_11, n_14, n_110, n_112, n_7, n_117, n_3, n_119, n_5, n_4, n_109, n_115, n_1, n_118, n_13, n_113, n_15);

input n_108;
input n_8;
input n_116;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_118;
input n_13;
input n_113;

output n_15;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

MAJx2_ASAP7_75t_L g60 ( 
.A(n_0),
.B(n_61),
.C(n_85),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_63),
.B(n_73),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_2),
.B(n_43),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_4),
.B(n_91),
.CON(n_90),
.SN(n_90)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

AOI322xp5_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_40),
.A3(n_53),
.B1(n_56),
.B2(n_94),
.C1(n_96),
.C2(n_119),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_6),
.Y(n_102)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_7),
.B(n_29),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_9),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_SL g74 ( 
.A(n_12),
.B(n_65),
.C(n_70),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_23),
.Y(n_15)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_99),
.B(n_103),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI31xp67_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_34),
.A3(n_60),
.B(n_89),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_39),
.C(n_46),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_35),
.B(n_48),
.C(n_95),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

OAI321xp33_ASAP7_75t_L g89 ( 
.A1(n_39),
.A2(n_46),
.A3(n_90),
.B1(n_92),
.B2(n_93),
.C(n_118),
.Y(n_89)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_79),
.C(n_80),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.C(n_69),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_108),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_109),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_110),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_111),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_112),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_113),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_114),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_115),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_116),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_117),
.Y(n_86)
);


endmodule