module real_jpeg_24623_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_29),
.B1(n_96),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_73),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_73),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx8_ASAP7_75t_SL g48 ( 
.A(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_9),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_82),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_9),
.A2(n_54),
.B(n_67),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_38),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_85),
.B1(n_166),
.B2(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_9),
.A2(n_25),
.B(n_181),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_92),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_19),
.B(n_92),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_63),
.C(n_78),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_20),
.A2(n_21),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_43),
.C(n_49),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_24),
.A2(n_31),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_26),
.B1(n_32),
.B2(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_26),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_32),
.A3(n_34),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_47),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_82),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_26),
.A2(n_46),
.A3(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_30),
.A2(n_38),
.B1(n_39),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_30),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_33),
.A2(n_34),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_33),
.B(n_36),
.Y(n_83)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_34),
.A2(n_69),
.B(n_82),
.C(n_140),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_44),
.A2(n_118),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_45),
.B(n_120),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_46),
.A2(n_47),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_57),
.Y(n_50)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_51),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_54),
.B1(n_67),
.B2(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_53),
.B(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_60),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_63),
.A2(n_78),
.B1(n_79),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_74),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_64),
.A2(n_70),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_75),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_65),
.A2(n_77),
.B1(n_138),
.B2(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_65),
.A2(n_72),
.B1(n_77),
.B2(n_146),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_70),
.B(n_82),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_80),
.B(n_84),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_81),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_98),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_97),
.B(n_123),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_169),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_85),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_85),
.A2(n_152),
.B1(n_157),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_87),
.B(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_110),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_100),
.B1(n_105),
.B2(n_106),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_190),
.B(n_196),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_175),
.B(n_189),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_153),
.B(n_174),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_147),
.C(n_148),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_162),
.B(n_173),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_160),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_167),
.B(n_172),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_177),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);


endmodule