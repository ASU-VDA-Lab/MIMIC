module real_jpeg_10826_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_326, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_326;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_25),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_2),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_2),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_67),
.B1(n_68),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_3),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_147),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_147),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_3),
.A2(n_25),
.B1(n_35),
.B2(n_147),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_25),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_4),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_4),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_52),
.B(n_65),
.C(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_52),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_10),
.A2(n_25),
.B1(n_35),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_10),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_10),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_60),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_67),
.B1(n_68),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_11),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_88),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_88),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_11),
.A2(n_25),
.B1(n_35),
.B2(n_88),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_67),
.B1(n_68),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_12),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_93),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_93),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_12),
.A2(n_25),
.B1(n_35),
.B2(n_93),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_14),
.A2(n_34),
.B1(n_52),
.B2(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_14),
.A2(n_34),
.B1(n_67),
.B2(n_68),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_15),
.A2(n_52),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_52),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_15),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_15),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_15),
.A2(n_30),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_15),
.B(n_30),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_15),
.B(n_32),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_15),
.A2(n_27),
.B(n_31),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_15),
.A2(n_25),
.B1(n_35),
.B2(n_113),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_16),
.A2(n_67),
.B1(n_68),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_16),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_129),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_129),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_16),
.A2(n_25),
.B1(n_35),
.B2(n_129),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_17),
.A2(n_52),
.B1(n_53),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_17),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_17),
.A2(n_67),
.B1(n_68),
.B2(n_100),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_17),
.A2(n_25),
.B1(n_35),
.B2(n_100),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B(n_33),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_23),
.A2(n_32),
.B1(n_37),
.B2(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_23),
.A2(n_32),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_24),
.A2(n_29),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_24),
.A2(n_29),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_24),
.A2(n_29),
.B1(n_210),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_24),
.A2(n_29),
.B1(n_235),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_24),
.A2(n_29),
.B1(n_253),
.B2(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_24),
.A2(n_29),
.B1(n_59),
.B2(n_274),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_25),
.A2(n_26),
.B(n_113),
.C(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_36),
.B(n_43),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_75),
.B(n_322),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_71),
.C(n_73),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_44),
.A2(n_45),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_57),
.C(n_63),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_46),
.A2(n_47),
.B1(n_63),
.B2(n_300),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_51),
.B(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_48),
.A2(n_51),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_48),
.A2(n_51),
.B1(n_138),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_48),
.A2(n_51),
.B1(n_155),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_48),
.A2(n_51),
.B1(n_195),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_48),
.A2(n_51),
.B1(n_206),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_48),
.A2(n_51),
.B1(n_232),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_48),
.A2(n_51),
.B1(n_250),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_48),
.A2(n_51),
.B1(n_55),
.B2(n_267),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_50),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_52),
.B(n_54),
.Y(n_142)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_53),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_57),
.A2(n_58),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_63),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_63),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_70),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_66),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_64),
.A2(n_66),
.B1(n_99),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_64),
.A2(n_66),
.B1(n_126),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_64),
.A2(n_66),
.B1(n_134),
.B2(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_64),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_64),
.A2(n_66),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_64),
.A2(n_66),
.B1(n_218),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_64),
.A2(n_66),
.B1(n_227),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_64),
.A2(n_66),
.B1(n_70),
.B2(n_259),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_71),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_315),
.B(n_321),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_292),
.A3(n_310),
.B1(n_313),
.B2(n_314),
.C(n_325),
.Y(n_76)
);

AOI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_243),
.A3(n_280),
.B1(n_286),
.B2(n_291),
.C(n_326),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_200),
.C(n_239),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_170),
.B(n_199),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_149),
.B(n_169),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_131),
.B(n_148),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_120),
.B(n_130),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_106),
.B(n_119),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_85),
.B(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_89),
.A2(n_90),
.B1(n_146),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_110),
.B1(n_111),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_105),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_114),
.B(n_118),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_111),
.B1(n_128),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_110),
.A2(n_111),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_110),
.A2(n_111),
.B1(n_181),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_110),
.A2(n_111),
.B1(n_215),
.B2(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_110),
.A2(n_111),
.B(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_132),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.CI(n_127),
.CON(n_123),
.SN(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.CI(n_139),
.CON(n_132),
.SN(n_132)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_162),
.B2(n_163),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_165),
.C(n_167),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_159),
.C(n_161),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_172),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_185),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_184),
.C(n_185),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_193),
.B2(n_194),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_193),
.C(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_201),
.A2(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_220),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_202),
.B(n_220),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_213),
.C(n_219),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_219),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_237),
.B2(n_238),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_228),
.C(n_238),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_226),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_233),
.C(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_231),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_262),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_244),
.B(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_255),
.C(n_261),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_246),
.B1(n_255),
.B2(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_251),
.C(n_254),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_257),
.B1(n_273),
.B2(n_275),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_256),
.A2(n_273),
.B(n_276),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_278),
.B2(n_279),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_270),
.C(n_279),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_268),
.B(n_269),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_268),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_294),
.C(n_302),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_269),
.B(n_294),
.CI(n_302),
.CON(n_312),
.SN(n_312)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_276),
.B2(n_277),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_287),
.B(n_290),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_303),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_303),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_296),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_300),
.C(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_305),
.C(n_309),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_299),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_320),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_317),
.Y(n_319)
);


endmodule