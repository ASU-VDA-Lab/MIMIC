module real_jpeg_7219_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_2),
.B(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_2),
.A2(n_210),
.B(n_259),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_2),
.B(n_187),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_2),
.B(n_369),
.C(n_372),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g374 ( 
.A1(n_2),
.A2(n_83),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_2),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_2),
.B(n_143),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_2),
.A2(n_32),
.B1(n_412),
.B2(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_3),
.A2(n_42),
.B1(n_45),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_50),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_50),
.B1(n_83),
.B2(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_50),
.B1(n_146),
.B2(n_229),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_4),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_126),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_4),
.A2(n_126),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_4),
.A2(n_126),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_6),
.A2(n_108),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_6),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_6),
.A2(n_192),
.B1(n_254),
.B2(n_291),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_6),
.A2(n_291),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_6),
.A2(n_291),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_82),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_33),
.B1(n_82),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_7),
.A2(n_82),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_59),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_54),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_8),
.A2(n_54),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_8),
.A2(n_54),
.B1(n_273),
.B2(n_275),
.Y(n_272)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_9),
.Y(n_307)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_11),
.Y(n_257)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_14),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_14),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_15),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_15),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_15),
.A2(n_148),
.B1(n_184),
.B2(n_281),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_15),
.A2(n_34),
.B1(n_184),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_15),
.A2(n_59),
.B1(n_184),
.B2(n_452),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_16),
.A2(n_108),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_16),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_16),
.A2(n_128),
.B1(n_288),
.B2(n_338),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_16),
.A2(n_59),
.B1(n_288),
.B2(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_16),
.A2(n_288),
.B1(n_413),
.B2(n_415),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_17),
.Y(n_371)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_493),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_483),
.B(n_492),
.Y(n_25)
);

OAI31xp33_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_216),
.A3(n_239),
.B(n_480),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_195),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_28),
.B(n_195),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_118),
.C(n_158),
.Y(n_28)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_29),
.B(n_118),
.CI(n_158),
.CON(n_357),
.SN(n_357)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_84),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_30),
.A2(n_31),
.B(n_86),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_51),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_31),
.A2(n_85),
.B1(n_86),
.B2(n_117),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_31),
.A2(n_51),
.B1(n_85),
.B2(n_349),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_41),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_32),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_32),
.A2(n_262),
.B1(n_268),
.B2(n_272),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_32),
.A2(n_272),
.B(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_32),
.A2(n_167),
.B(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_32),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_32),
.A2(n_306),
.B1(n_400),
.B2(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_32),
.A2(n_41),
.B(n_304),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_33),
.Y(n_264)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_36),
.Y(n_277)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_38),
.Y(n_332)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_38),
.Y(n_424)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_41),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_44),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_48),
.Y(n_414)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_49),
.Y(n_267)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_49),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_51),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_62),
.B(n_77),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_53),
.A2(n_63),
.B1(n_78),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_130)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_57),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_57),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_57),
.Y(n_388)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_62),
.B(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_62),
.A2(n_151),
.B(n_152),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_62),
.A2(n_77),
.B(n_152),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_62),
.A2(n_151),
.B1(n_156),
.B2(n_174),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_62),
.A2(n_464),
.B(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_63),
.A2(n_78),
.B1(n_374),
.B2(n_377),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_63),
.A2(n_78),
.B1(n_377),
.B2(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_63),
.A2(n_78),
.B1(n_386),
.B2(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_64)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_65),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_72),
.Y(n_372)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_105),
.B(n_110),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_87),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_87),
.A2(n_187),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_87),
.A2(n_187),
.B1(n_286),
.B2(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_88),
.A2(n_181),
.B(n_186),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_88),
.A2(n_116),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_88),
.A2(n_116),
.B1(n_181),
.B2(n_290),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_88),
.A2(n_489),
.B(n_490),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_100),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_100),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_100),
.Y(n_449)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_101),
.Y(n_284)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_101),
.Y(n_340)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_103),
.Y(n_441)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_104),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_105),
.B(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_107),
.Y(n_292)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_110),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_114),
.Y(n_238)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_116),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_116),
.A2(n_206),
.B(n_212),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_149),
.B(n_157),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_129),
.B1(n_143),
.B2(n_144),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_121),
.A2(n_130),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_137),
.B1(n_139),
.B2(n_141),
.Y(n_136)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_129),
.B(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_129),
.A2(n_144),
.B(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_129),
.A2(n_227),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_129),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_129),
.A2(n_143),
.B1(n_337),
.B2(n_448),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_129),
.A2(n_143),
.B(n_487),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_130),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_130),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_130),
.A2(n_299),
.B1(n_300),
.B2(n_336),
.Y(n_335)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_131),
.Y(n_376)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_132),
.Y(n_443)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_134),
.Y(n_437)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_143),
.B(n_191),
.Y(n_202)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g432 ( 
.A1(n_148),
.A2(n_433),
.A3(n_435),
.B1(n_438),
.B2(n_442),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_150),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_151),
.B(n_375),
.Y(n_410)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_153),
.Y(n_444)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_196),
.CI(n_215),
.CON(n_195),
.SN(n_195)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_179),
.C(n_188),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_159),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_171),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_160),
.A2(n_171),
.B1(n_172),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_160),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_162),
.A2(n_263),
.B(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_163),
.Y(n_308)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_169),
.Y(n_420)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_175),
.Y(n_452)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_177),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_179),
.A2(n_180),
.B1(n_188),
.B2(n_189),
.Y(n_351)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_186),
.B(n_212),
.Y(n_495)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_195),
.B(n_218),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_205),
.B2(n_214),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_204),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_199),
.B(n_224),
.C(n_232),
.Y(n_491)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_202),
.A2(n_228),
.B(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_205),
.B(n_219),
.C(n_222),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_217),
.A2(n_481),
.B(n_482),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_228),
.Y(n_487)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_234),
.Y(n_489)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_358),
.B(n_474),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_343),
.C(n_355),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_322),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_242),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_310),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_243),
.B(n_310),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_293),
.C(n_302),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_244),
.B(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_278),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_245),
.B(n_279),
.C(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_261),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_246),
.B(n_261),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_250),
.A3(n_251),
.B1(n_253),
.B2(n_258),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_266),
.Y(n_395)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_275),
.Y(n_401)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_276),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_302),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.C(n_298),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_294),
.B(n_295),
.CI(n_298),
.CON(n_324),
.SN(n_324)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

INVx3_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_313),
.C(n_315),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_320),
.C(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_341),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_323),
.B(n_341),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.C(n_326),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_324),
.B(n_472),
.Y(n_471)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_324),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_325),
.B(n_326),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_333),
.C(n_335),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_327),
.A2(n_328),
.B1(n_333),
.B2(n_334),
.Y(n_459)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_335),
.B(n_459),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

A2O1A1O1Ixp25_ASAP7_75t_L g474 ( 
.A1(n_343),
.A2(n_355),
.B(n_475),
.C(n_478),
.D(n_479),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_354),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_344),
.B(n_354),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_348),
.C(n_353),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_350),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_356),
.B(n_357),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_357),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_469),
.B(n_473),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_454),
.B(n_468),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_428),
.B(n_453),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_396),
.B(n_427),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_381),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_363),
.B(n_381),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_373),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_373),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_375),
.B(n_439),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_SL g448 ( 
.A1(n_375),
.A2(n_438),
.B(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_393),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_392),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_392),
.C(n_393),
.Y(n_429)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_385),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_408),
.B(n_426),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_407),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_407),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_401),
.B(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_418),
.B(n_425),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_410),
.B(n_411),
.Y(n_425)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_430),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_446),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_447),
.C(n_450),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_445),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_451),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_455),
.B(n_456),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_460),
.B2(n_461),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_463),
.C(n_466),
.Y(n_470)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_467),
.Y(n_461)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_462),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_463),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_471),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_485),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_485),
.B(n_495),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_485),
.Y(n_498)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_488),
.CI(n_491),
.CON(n_485),
.SN(n_485)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_495),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);


endmodule