module fake_jpeg_1521_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_18),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_8),
.B1(n_16),
.B2(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_17),
.B1(n_13),
.B2(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_58),
.B1(n_47),
.B2(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_32),
.B1(n_26),
.B2(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_58),
.B1(n_47),
.B2(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_23),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_21),
.B(n_17),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_62),
.B1(n_63),
.B2(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_69),
.B1(n_49),
.B2(n_71),
.Y(n_86)
);

NOR4xp25_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_21),
.C(n_42),
.D(n_23),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_81),
.B(n_74),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_71),
.C(n_66),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_39),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_86),
.B1(n_52),
.B2(n_45),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_78),
.B(n_75),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_83),
.B(n_39),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_82),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_95),
.B(n_90),
.Y(n_96)
);

OAI31xp33_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_97),
.A3(n_39),
.B(n_49),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_88),
.B(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_19),
.C(n_28),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.Y(n_101)
);


endmodule