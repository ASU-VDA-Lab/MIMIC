module real_aes_7713_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_726, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_726;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g463 ( .A1(n_0), .A2(n_201), .B(n_464), .C(n_467), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_1), .B(n_458), .Y(n_468) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g236 ( .A(n_3), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_4), .B(n_153), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_5), .A2(n_453), .B(n_541), .Y(n_540) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_6), .A2(n_176), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_7), .A2(n_37), .B1(n_146), .B2(n_170), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_8), .B(n_176), .Y(n_248) );
AND2x6_ASAP7_75t_L g161 ( .A(n_9), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_10), .A2(n_161), .B(n_444), .C(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_11), .B(n_38), .Y(n_117) );
INVx1_ASAP7_75t_L g716 ( .A(n_11), .Y(n_716) );
INVx1_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_13), .B(n_151), .Y(n_184) );
INVx1_ASAP7_75t_L g228 ( .A(n_14), .Y(n_228) );
OAI22xp33_ASAP7_75t_SL g701 ( .A1(n_15), .A2(n_702), .B1(n_707), .B2(n_708), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_15), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_16), .B(n_153), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_17), .B(n_177), .Y(n_215) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_18), .A2(n_175), .A3(n_176), .B1(n_199), .B2(n_203), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_19), .B(n_146), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_20), .B(n_177), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_21), .A2(n_53), .B1(n_146), .B2(n_170), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g173 ( .A1(n_22), .A2(n_80), .B1(n_146), .B2(n_151), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_23), .B(n_146), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_24), .A2(n_175), .B(n_444), .C(n_491), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_25), .A2(n_175), .B(n_444), .C(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_26), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_27), .B(n_138), .Y(n_257) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_28), .A2(n_90), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_28), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_29), .A2(n_453), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_30), .B(n_138), .Y(n_163) );
INVx2_ASAP7_75t_L g148 ( .A(n_31), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_32), .A2(n_450), .B(n_476), .C(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_33), .B(n_146), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_34), .B(n_138), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g705 ( .A1(n_35), .A2(n_42), .B1(n_434), .B2(n_706), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_35), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_36), .B(n_186), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_38), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_39), .B(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_40), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_41), .B(n_153), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_42), .A2(n_129), .B1(n_434), .B2(n_435), .Y(n_128) );
INVx1_ASAP7_75t_L g434 ( .A(n_42), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_43), .B(n_453), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_44), .A2(n_450), .B(n_476), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_45), .B(n_146), .Y(n_243) );
INVx1_ASAP7_75t_L g465 ( .A(n_46), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_47), .A2(n_91), .B1(n_170), .B2(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g528 ( .A(n_48), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_49), .B(n_146), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_50), .B(n_146), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_51), .B(n_453), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_52), .B(n_234), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g219 ( .A1(n_54), .A2(n_58), .B1(n_146), .B2(n_151), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_55), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_56), .B(n_146), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_57), .B(n_146), .Y(n_256) );
INVx1_ASAP7_75t_L g162 ( .A(n_59), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_60), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_61), .B(n_458), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_62), .A2(n_231), .B(n_234), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_63), .B(n_146), .Y(n_237) );
INVx1_ASAP7_75t_L g141 ( .A(n_64), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_65), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_66), .B(n_153), .Y(n_481) );
AO32x2_ASAP7_75t_L g167 ( .A1(n_67), .A2(n_168), .A3(n_174), .B1(n_175), .B2(n_176), .Y(n_167) );
AOI22xp5_ASAP7_75t_SL g118 ( .A1(n_68), .A2(n_114), .B1(n_119), .B2(n_697), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_69), .B(n_154), .Y(n_518) );
INVx1_ASAP7_75t_L g255 ( .A(n_70), .Y(n_255) );
INVx1_ASAP7_75t_L g149 ( .A(n_71), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_72), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_73), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_74), .B(n_480), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_75), .A2(n_444), .B(n_446), .C(n_450), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_76), .B(n_151), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_77), .Y(n_542) );
INVx1_ASAP7_75t_L g721 ( .A(n_78), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_79), .B(n_479), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_81), .B(n_170), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_82), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_83), .B(n_151), .Y(n_158) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
AOI22xp33_ASAP7_75t_SL g102 ( .A1(n_85), .A2(n_103), .B1(n_711), .B2(n_722), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_86), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_87), .B(n_172), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_88), .B(n_151), .Y(n_244) );
OR2x2_ASAP7_75t_L g113 ( .A(n_89), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_90), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_92), .A2(n_101), .B1(n_151), .B2(n_152), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_93), .B(n_453), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_94), .Y(n_478) );
INVxp67_ASAP7_75t_L g545 ( .A(n_95), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_96), .B(n_151), .Y(n_253) );
INVx1_ASAP7_75t_L g447 ( .A(n_97), .Y(n_447) );
INVx1_ASAP7_75t_L g514 ( .A(n_98), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_99), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g530 ( .A(n_100), .B(n_138), .Y(n_530) );
AOI22x1_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_108), .B1(n_118), .B2(n_700), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_109), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_109), .A2(n_701), .B(n_709), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g710 ( .A(n_113), .Y(n_710) );
NOR2x2_ASAP7_75t_L g699 ( .A(n_114), .B(n_127), .Y(n_699) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
NAND3xp33_ASAP7_75t_SL g718 ( .A(n_116), .B(n_127), .C(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_124), .B2(n_696), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
INVxp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g696 ( .A(n_126), .Y(n_696) );
AO22x2_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_128), .B1(n_436), .B2(n_695), .Y(n_126) );
INVx1_ASAP7_75t_L g695 ( .A(n_127), .Y(n_695) );
INVx1_ASAP7_75t_L g435 ( .A(n_129), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g703 ( .A1(n_129), .A2(n_435), .B1(n_704), .B2(n_705), .Y(n_703) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_355), .Y(n_129) );
NAND3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_304), .C(n_346), .Y(n_130) );
AOI211xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_209), .B(n_258), .C(n_280), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_164), .B(n_192), .C(n_204), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_134), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g367 ( .A(n_134), .B(n_284), .Y(n_367) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g269 ( .A(n_135), .B(n_195), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_135), .B(n_180), .Y(n_386) );
INVx1_ASAP7_75t_L g404 ( .A(n_135), .Y(n_404) );
AND2x2_ASAP7_75t_L g413 ( .A(n_135), .B(n_301), .Y(n_413) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g296 ( .A(n_136), .B(n_180), .Y(n_296) );
AND2x2_ASAP7_75t_L g354 ( .A(n_136), .B(n_301), .Y(n_354) );
INVx1_ASAP7_75t_L g398 ( .A(n_136), .Y(n_398) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g275 ( .A(n_137), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g283 ( .A(n_137), .Y(n_283) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_137), .Y(n_323) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_143), .B(n_163), .Y(n_137) );
INVx2_ASAP7_75t_L g174 ( .A(n_138), .Y(n_174) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_138), .A2(n_181), .B(n_191), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_138), .A2(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g497 ( .A(n_138), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_138), .A2(n_525), .B(n_526), .Y(n_524) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_L g177 ( .A(n_139), .B(n_140), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_156), .B(n_161), .Y(n_143) );
O2A1O1Ixp5_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_149), .B(n_150), .C(n_153), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_146), .Y(n_449) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
AND2x6_ASAP7_75t_L g444 ( .A(n_147), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g152 ( .A(n_148), .Y(n_152) );
INVx1_ASAP7_75t_L g235 ( .A(n_148), .Y(n_235) );
INVx2_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g201 ( .A(n_153), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_153), .A2(n_243), .B(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_153), .A2(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_153), .B(n_545), .Y(n_544) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_154), .A2(n_169), .B1(n_172), .B2(n_173), .Y(n_168) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_155), .Y(n_160) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
INVx1_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
INVx1_ASAP7_75t_L g445 ( .A(n_155), .Y(n_445) );
AND2x2_ASAP7_75t_L g454 ( .A(n_155), .B(n_235), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g231 ( .A(n_159), .Y(n_231) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g480 ( .A(n_160), .Y(n_480) );
BUFx3_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_161), .A2(n_182), .B(n_187), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_161), .A2(n_227), .B(n_232), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_161), .A2(n_242), .B(n_245), .Y(n_241) );
INVx4_ASAP7_75t_SL g451 ( .A(n_161), .Y(n_451) );
AND2x4_ASAP7_75t_L g453 ( .A(n_161), .B(n_454), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_161), .B(n_454), .Y(n_515) );
INVxp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_178), .Y(n_165) );
AND2x2_ASAP7_75t_L g262 ( .A(n_166), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g295 ( .A(n_166), .Y(n_295) );
OR2x2_ASAP7_75t_L g421 ( .A(n_166), .B(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_166), .B(n_180), .Y(n_425) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
INVx1_ASAP7_75t_L g207 ( .A(n_167), .Y(n_207) );
AND2x2_ASAP7_75t_L g284 ( .A(n_167), .B(n_197), .Y(n_284) );
AND2x2_ASAP7_75t_L g324 ( .A(n_167), .B(n_198), .Y(n_324) );
INVx2_ASAP7_75t_L g467 ( .A(n_171), .Y(n_467) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_171), .Y(n_482) );
INVx2_ASAP7_75t_L g190 ( .A(n_172), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_172), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_172), .A2(n_201), .B1(n_218), .B2(n_219), .Y(n_217) );
INVx4_ASAP7_75t_L g466 ( .A(n_172), .Y(n_466) );
INVx1_ASAP7_75t_L g494 ( .A(n_174), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g216 ( .A(n_175), .B(n_217), .C(n_220), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_175), .A2(n_251), .B(n_254), .Y(n_250) );
INVx4_ASAP7_75t_L g220 ( .A(n_176), .Y(n_220) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_176), .A2(n_241), .B(n_248), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_176), .A2(n_504), .B(n_505), .Y(n_503) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_176), .Y(n_539) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g203 ( .A(n_177), .Y(n_203) );
INVxp67_ASAP7_75t_L g366 ( .A(n_178), .Y(n_366) );
AND2x4_ASAP7_75t_L g391 ( .A(n_178), .B(n_284), .Y(n_391) );
BUFx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_179), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g196 ( .A(n_180), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g270 ( .A(n_180), .B(n_198), .Y(n_270) );
INVx1_ASAP7_75t_L g276 ( .A(n_180), .Y(n_276) );
INVx2_ASAP7_75t_L g302 ( .A(n_180), .Y(n_302) );
AND2x2_ASAP7_75t_L g318 ( .A(n_180), .B(n_319), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
O2A1O1Ixp5_ASAP7_75t_L g254 ( .A1(n_190), .A2(n_233), .B(n_255), .C(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_193), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_196), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx2_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
AND2x2_ASAP7_75t_L g381 ( .A(n_195), .B(n_197), .Y(n_381) );
AND2x2_ASAP7_75t_L g298 ( .A(n_196), .B(n_283), .Y(n_298) );
AND2x2_ASAP7_75t_L g397 ( .A(n_196), .B(n_398), .Y(n_397) );
NOR2xp67_ASAP7_75t_L g319 ( .A(n_197), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g422 ( .A(n_197), .B(n_283), .Y(n_422) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g208 ( .A(n_198), .Y(n_208) );
AND2x2_ASAP7_75t_L g301 ( .A(n_198), .B(n_302), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_233), .B(n_236), .C(n_237), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_201), .A2(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g225 ( .A(n_203), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_203), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
AND2x2_ASAP7_75t_L g347 ( .A(n_206), .B(n_282), .Y(n_347) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_207), .B(n_283), .Y(n_332) );
INVx2_ASAP7_75t_L g331 ( .A(n_208), .Y(n_331) );
OAI222xp33_ASAP7_75t_L g335 ( .A1(n_208), .A2(n_275), .B1(n_336), .B2(n_338), .C1(n_339), .C2(n_342), .Y(n_335) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g260 ( .A(n_213), .Y(n_260) );
OR2x2_ASAP7_75t_L g371 ( .A(n_213), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g293 ( .A(n_214), .Y(n_293) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_214), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g350 ( .A(n_214), .B(n_264), .Y(n_350) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g311 ( .A(n_215), .Y(n_311) );
AO21x1_ASAP7_75t_L g310 ( .A1(n_217), .A2(n_220), .B(n_311), .Y(n_310) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_220), .A2(n_442), .B(n_455), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_220), .B(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g458 ( .A(n_220), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_220), .B(n_484), .Y(n_483) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_220), .A2(n_513), .B(n_520), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_221), .A2(n_314), .B1(n_353), .B2(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_239), .Y(n_221) );
INVx3_ASAP7_75t_L g286 ( .A(n_222), .Y(n_286) );
OR2x2_ASAP7_75t_L g419 ( .A(n_222), .B(n_295), .Y(n_419) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g292 ( .A(n_223), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_223), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_223), .B(n_264), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_223), .B(n_240), .Y(n_372) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g263 ( .A(n_224), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g267 ( .A(n_224), .B(n_240), .Y(n_267) );
AND2x2_ASAP7_75t_L g343 ( .A(n_224), .B(n_290), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_224), .B(n_249), .Y(n_383) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_238), .Y(n_224) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_225), .A2(n_250), .B(n_257), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .C(n_231), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_229), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_229), .A2(n_518), .B(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_231), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_233), .A2(n_492), .B(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_239), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_239), .B(n_260), .Y(n_299) );
AND2x2_ASAP7_75t_L g303 ( .A(n_239), .B(n_293), .Y(n_303) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
INVx3_ASAP7_75t_L g264 ( .A(n_240), .Y(n_264) );
AND2x2_ASAP7_75t_L g289 ( .A(n_240), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g424 ( .A(n_240), .B(n_407), .Y(n_424) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_249), .Y(n_278) );
INVx2_ASAP7_75t_L g290 ( .A(n_249), .Y(n_290) );
AND2x2_ASAP7_75t_L g334 ( .A(n_249), .B(n_310), .Y(n_334) );
INVx1_ASAP7_75t_L g377 ( .A(n_249), .Y(n_377) );
OR2x2_ASAP7_75t_L g408 ( .A(n_249), .B(n_310), .Y(n_408) );
AND2x2_ASAP7_75t_L g428 ( .A(n_249), .B(n_264), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_261), .B(n_265), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g266 ( .A(n_260), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_260), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g385 ( .A(n_262), .Y(n_385) );
INVx2_ASAP7_75t_SL g279 ( .A(n_263), .Y(n_279) );
AND2x2_ASAP7_75t_L g399 ( .A(n_263), .B(n_293), .Y(n_399) );
INVx2_ASAP7_75t_L g345 ( .A(n_264), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_264), .B(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .B1(n_271), .B2(n_277), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_267), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g433 ( .A(n_267), .Y(n_433) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g358 ( .A(n_269), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_269), .B(n_301), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_270), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g374 ( .A(n_270), .B(n_323), .Y(n_374) );
INVx2_ASAP7_75t_L g430 ( .A(n_270), .Y(n_430) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g300 ( .A(n_273), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_273), .B(n_318), .Y(n_351) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_275), .B(n_295), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g412 ( .A(n_278), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_SL g362 ( .A1(n_279), .A2(n_363), .B(n_365), .C(n_368), .Y(n_362) );
OR2x2_ASAP7_75t_L g389 ( .A(n_279), .B(n_293), .Y(n_389) );
OAI221xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_285), .B1(n_287), .B2(n_294), .C(n_297), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_282), .B(n_331), .Y(n_338) );
AND2x2_ASAP7_75t_L g380 ( .A(n_282), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g416 ( .A(n_282), .Y(n_416) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
INVx1_ASAP7_75t_L g320 ( .A(n_283), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_286), .B(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g394 ( .A(n_286), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_286), .B(n_334), .Y(n_410) );
INVx2_ASAP7_75t_L g396 ( .A(n_287), .Y(n_396) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g337 ( .A(n_289), .B(n_308), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_289), .A2(n_305), .B(n_347), .C(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g315 ( .A(n_290), .B(n_310), .Y(n_315) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_294), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OR2x2_ASAP7_75t_L g363 ( .A(n_295), .B(n_364), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_300), .B2(n_303), .Y(n_297) );
INVx1_ASAP7_75t_L g417 ( .A(n_299), .Y(n_417) );
INVx1_ASAP7_75t_L g364 ( .A(n_301), .Y(n_364) );
INVx1_ASAP7_75t_L g415 ( .A(n_303), .Y(n_415) );
AOI211xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_308), .B(n_312), .C(n_335), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g327 ( .A(n_307), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g378 ( .A(n_308), .Y(n_378) );
AND2x2_ASAP7_75t_L g427 ( .A(n_308), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_317), .B(n_325), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_315), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g333 ( .A(n_316), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g409 ( .A(n_316), .Y(n_409) );
OAI32xp33_ASAP7_75t_L g420 ( .A1(n_316), .A2(n_368), .A3(n_375), .B1(n_416), .B2(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_SL g388 ( .A(n_318), .Y(n_388) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g328 ( .A(n_324), .Y(n_328) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B(n_333), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_327), .A2(n_375), .B1(n_401), .B2(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_331), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g361 ( .A(n_345), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_354), .A2(n_396), .B1(n_397), .B2(n_399), .C(n_400), .Y(n_395) );
NAND5xp2_ASAP7_75t_L g355 ( .A(n_356), .B(n_379), .C(n_395), .D(n_405), .E(n_423), .Y(n_355) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_359), .B(n_362), .C(n_369), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g426 ( .A(n_363), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_373), .B2(n_375), .Y(n_369) );
INVx1_ASAP7_75t_SL g402 ( .A(n_372), .Y(n_402) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI322xp33_ASAP7_75t_L g384 ( .A1(n_375), .A2(n_385), .A3(n_386), .B1(n_387), .B2(n_388), .C1(n_389), .C2(n_390), .Y(n_384) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g387 ( .A(n_377), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_377), .B(n_402), .Y(n_401) );
AOI211xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_382), .B(n_384), .C(n_392), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_388), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_414) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_413), .B1(n_414), .B2(n_418), .C(n_420), .Y(n_405) );
OAI211xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_409), .B(n_410), .C(n_411), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g432 ( .A(n_408), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_426), .B2(n_427), .C(n_429), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_431), .B(n_432), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_437), .B(n_638), .Y(n_436) );
AND4x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_578), .C(n_593), .D(n_618), .Y(n_437) );
NOR2xp33_ASAP7_75t_SL g438 ( .A(n_439), .B(n_551), .Y(n_438) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_469), .B(n_531), .Y(n_439) );
AND2x2_ASAP7_75t_L g581 ( .A(n_440), .B(n_486), .Y(n_581) );
AND2x2_ASAP7_75t_L g594 ( .A(n_440), .B(n_485), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_440), .B(n_470), .Y(n_644) );
INVx1_ASAP7_75t_L g648 ( .A(n_440), .Y(n_648) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_457), .Y(n_440) );
INVx2_ASAP7_75t_L g565 ( .A(n_441), .Y(n_565) );
BUFx2_ASAP7_75t_L g592 ( .A(n_441), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_452), .Y(n_442) );
INVx5_ASAP7_75t_L g462 ( .A(n_444), .Y(n_462) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g460 ( .A1(n_451), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_451), .A2(n_462), .B(n_542), .C(n_543), .Y(n_541) );
BUFx2_ASAP7_75t_L g489 ( .A(n_453), .Y(n_489) );
AND2x2_ASAP7_75t_L g532 ( .A(n_457), .B(n_486), .Y(n_532) );
INVx2_ASAP7_75t_L g548 ( .A(n_457), .Y(n_548) );
AND2x2_ASAP7_75t_L g557 ( .A(n_457), .B(n_485), .Y(n_557) );
AND2x2_ASAP7_75t_L g636 ( .A(n_457), .B(n_565), .Y(n_636) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_468), .Y(n_457) );
INVx2_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_498), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_470), .B(n_563), .Y(n_601) );
INVx1_ASAP7_75t_L g689 ( .A(n_470), .Y(n_689) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_485), .Y(n_470) );
AND2x2_ASAP7_75t_L g547 ( .A(n_471), .B(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g561 ( .A(n_471), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_471), .Y(n_590) );
OR2x2_ASAP7_75t_L g622 ( .A(n_471), .B(n_564), .Y(n_622) );
AND2x2_ASAP7_75t_L g630 ( .A(n_471), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g663 ( .A(n_471), .B(n_632), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_471), .B(n_532), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_471), .B(n_592), .Y(n_688) );
AND2x2_ASAP7_75t_L g694 ( .A(n_471), .B(n_581), .Y(n_694) );
INVx5_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g554 ( .A(n_472), .Y(n_554) );
AND2x2_ASAP7_75t_L g584 ( .A(n_472), .B(n_564), .Y(n_584) );
AND2x2_ASAP7_75t_L g617 ( .A(n_472), .B(n_577), .Y(n_617) );
AND2x2_ASAP7_75t_L g637 ( .A(n_472), .B(n_486), .Y(n_637) );
AND2x2_ASAP7_75t_L g671 ( .A(n_472), .B(n_537), .Y(n_671) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_481), .C(n_482), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_479), .A2(n_482), .B(n_528), .C(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g577 ( .A(n_485), .B(n_548), .Y(n_577) );
AND2x2_ASAP7_75t_L g588 ( .A(n_485), .B(n_584), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_485), .B(n_564), .Y(n_627) );
INVx2_ASAP7_75t_L g642 ( .A(n_485), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_485), .B(n_576), .Y(n_665) );
AND2x2_ASAP7_75t_L g684 ( .A(n_485), .B(n_636), .Y(n_684) );
INVx5_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
AND2x2_ASAP7_75t_L g591 ( .A(n_486), .B(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g632 ( .A(n_486), .B(n_548), .Y(n_632) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .Y(n_486) );
AOI21xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_490), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
AND2x2_ASAP7_75t_L g555 ( .A(n_500), .B(n_538), .Y(n_555) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_501), .B(n_512), .Y(n_535) );
OR2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_538), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_501), .B(n_538), .Y(n_573) );
AND2x2_ASAP7_75t_L g600 ( .A(n_501), .B(n_537), .Y(n_600) );
AND2x2_ASAP7_75t_L g652 ( .A(n_501), .B(n_511), .Y(n_652) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_502), .B(n_522), .Y(n_560) );
AND2x2_ASAP7_75t_L g596 ( .A(n_502), .B(n_512), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_509), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g586 ( .A(n_510), .B(n_568), .Y(n_586) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
OAI322xp33_ASAP7_75t_L g551 ( .A1(n_511), .A2(n_552), .A3(n_556), .B1(n_558), .B2(n_561), .C1(n_566), .C2(n_574), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_511), .B(n_537), .Y(n_559) );
OR2x2_ASAP7_75t_L g569 ( .A(n_511), .B(n_523), .Y(n_569) );
AND2x2_ASAP7_75t_L g571 ( .A(n_511), .B(n_523), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_511), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_511), .B(n_538), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_511), .B(n_667), .Y(n_666) );
INVx5_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_512), .B(n_555), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_522), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g549 ( .A(n_522), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_522), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g611 ( .A(n_522), .B(n_538), .Y(n_611) );
AOI211xp5_ASAP7_75t_SL g639 ( .A1(n_522), .A2(n_640), .B(n_643), .C(n_655), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_522), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g677 ( .A(n_522), .B(n_652), .Y(n_677) );
INVx5_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g605 ( .A(n_523), .B(n_538), .Y(n_605) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
AND2x2_ASAP7_75t_L g654 ( .A(n_523), .B(n_652), .Y(n_654) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_523), .B(n_555), .Y(n_685) );
AND2x2_ASAP7_75t_L g692 ( .A(n_523), .B(n_651), .Y(n_692) );
OR2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_530), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_547), .B2(n_549), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_532), .B(n_554), .Y(n_602) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g550 ( .A(n_535), .Y(n_550) );
OR2x2_ASAP7_75t_L g610 ( .A(n_535), .B(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g658 ( .A1(n_535), .A2(n_659), .B1(n_661), .B2(n_662), .C(n_664), .Y(n_658) );
INVx2_ASAP7_75t_L g597 ( .A(n_536), .Y(n_597) );
AND2x2_ASAP7_75t_L g570 ( .A(n_537), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g660 ( .A(n_537), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_537), .B(n_652), .Y(n_673) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_L g615 ( .A(n_538), .Y(n_615) );
AND2x2_ASAP7_75t_L g651 ( .A(n_538), .B(n_652), .Y(n_651) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_546), .Y(n_538) );
AND2x2_ASAP7_75t_L g653 ( .A(n_547), .B(n_592), .Y(n_653) );
AND2x2_ASAP7_75t_L g563 ( .A(n_548), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_548), .B(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_SL g634 ( .A(n_550), .B(n_597), .Y(n_634) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g640 ( .A(n_553), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OR2x2_ASAP7_75t_L g626 ( .A(n_554), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g691 ( .A(n_554), .B(n_636), .Y(n_691) );
INVx2_ASAP7_75t_L g624 ( .A(n_555), .Y(n_624) );
NAND4xp25_ASAP7_75t_SL g687 ( .A(n_556), .B(n_688), .C(n_689), .D(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_557), .B(n_621), .Y(n_656) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_SL g693 ( .A(n_560), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_SL g655 ( .A1(n_561), .A2(n_624), .B(n_628), .C(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g650 ( .A(n_563), .B(n_642), .Y(n_650) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_564), .Y(n_576) );
INVx1_ASAP7_75t_L g631 ( .A(n_564), .Y(n_631) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B(n_570), .C(n_572), .Y(n_566) );
AND2x2_ASAP7_75t_L g587 ( .A(n_567), .B(n_571), .Y(n_587) );
OAI322xp33_ASAP7_75t_SL g625 ( .A1(n_567), .A2(n_626), .A3(n_628), .B1(n_629), .B2(n_633), .C1(n_634), .C2(n_635), .Y(n_625) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g647 ( .A(n_569), .B(n_573), .Y(n_647) );
INVx1_ASAP7_75t_L g628 ( .A(n_571), .Y(n_628) );
INVx1_ASAP7_75t_SL g646 ( .A(n_573), .Y(n_646) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI222xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_585), .B1(n_587), .B2(n_588), .C1(n_589), .C2(n_726), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_582), .Y(n_579) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_580), .A2(n_642), .A3(n_647), .B1(n_669), .B2(n_670), .C1(n_672), .C2(n_673), .Y(n_668) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_581), .A2(n_595), .B1(n_619), .B2(n_623), .C(n_625), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_586), .A2(n_599), .B1(n_601), .B2(n_602), .C1(n_603), .C2(n_606), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_588), .A2(n_595), .B1(n_665), .B2(n_666), .Y(n_664) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_598), .C(n_609), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_595), .A2(n_632), .B(n_675), .C(n_678), .Y(n_674) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g604 ( .A(n_596), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g667 ( .A(n_600), .Y(n_667) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_607), .B(n_632), .Y(n_661) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B(n_616), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g678 ( .A1(n_610), .A2(n_679), .B1(n_680), .B2(n_681), .C(n_682), .Y(n_678) );
INVxp33_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_614), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_621), .B(n_632), .Y(n_672) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g683 ( .A(n_636), .B(n_642), .Y(n_683) );
AND4x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_657), .C(n_674), .D(n_686), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_645), .B1(n_647), .B2(n_648), .C(n_649), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g679 ( .A(n_650), .Y(n_679) );
INVx1_ASAP7_75t_SL g669 ( .A(n_654), .Y(n_669) );
NOR2xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_668), .Y(n_657) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_670), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_677), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx3_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g708 ( .A(n_702), .Y(n_708) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx3_ASAP7_75t_SL g724 ( .A(n_713), .Y(n_724) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx14_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
endmodule