module fake_jpeg_913_n_505 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_505);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_505;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_18),
.Y(n_121)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_55),
.Y(n_144)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_66),
.B(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_18),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_67),
.B(n_94),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_32),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_96),
.Y(n_103)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_93),
.Y(n_118)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_99),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_22),
.Y(n_151)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_22),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_39),
.B1(n_30),
.B2(n_43),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_107),
.A2(n_115),
.B1(n_136),
.B2(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_47),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_R g193 ( 
.A(n_108),
.B(n_121),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_114),
.B(n_142),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_30),
.B1(n_22),
.B2(n_16),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_35),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_46),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_44),
.B1(n_43),
.B2(n_35),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_41),
.B1(n_84),
.B2(n_82),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_68),
.A2(n_39),
.B1(n_44),
.B2(n_33),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_17),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_22),
.B1(n_33),
.B2(n_16),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_55),
.A2(n_46),
.B1(n_20),
.B2(n_41),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_147),
.B1(n_39),
.B2(n_77),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_63),
.A2(n_39),
.B1(n_21),
.B2(n_31),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_69),
.B1(n_92),
.B2(n_53),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_168),
.B1(n_187),
.B2(n_130),
.Y(n_213)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_115),
.A2(n_61),
.B1(n_64),
.B2(n_52),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_169),
.B(n_194),
.Y(n_231)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_42),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_173),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_31),
.B(n_42),
.C(n_21),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_104),
.B(n_22),
.Y(n_173)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_178),
.A2(n_202),
.B1(n_159),
.B2(n_122),
.Y(n_232)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_198),
.B1(n_160),
.B2(n_122),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_70),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_191),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_136),
.B1(n_107),
.B2(n_79),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_195),
.B1(n_196),
.B2(n_130),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_156),
.A2(n_93),
.B1(n_87),
.B2(n_81),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_0),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_93),
.B1(n_87),
.B2(n_34),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_139),
.A2(n_155),
.B1(n_152),
.B2(n_140),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_201),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_111),
.A2(n_34),
.B1(n_24),
.B2(n_12),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_129),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

AOI22x1_ASAP7_75t_SL g202 ( 
.A1(n_109),
.A2(n_24),
.B1(n_34),
.B2(n_10),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_0),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_137),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_207),
.Y(n_238)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_125),
.B1(n_120),
.B2(n_102),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_232),
.B1(n_221),
.B2(n_213),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_179),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_216),
.A2(n_221),
.B1(n_226),
.B2(n_234),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_173),
.C(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_239),
.C(n_214),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_175),
.A2(n_132),
.B1(n_154),
.B2(n_150),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_236),
.B1(n_226),
.B2(n_220),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_109),
.B1(n_112),
.B2(n_110),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_112),
.B1(n_110),
.B2(n_101),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_161),
.A2(n_184),
.B1(n_182),
.B2(n_190),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_239),
.B(n_183),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_101),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_197),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_253),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_245),
.B(n_250),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g278 ( 
.A(n_247),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_208),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_252),
.C(n_258),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_171),
.B1(n_187),
.B2(n_192),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_243),
.B1(n_241),
.B2(n_237),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_212),
.A2(n_172),
.B(n_193),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_255),
.B(n_263),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_174),
.B(n_202),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_257),
.B1(n_274),
.B2(n_230),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_165),
.C(n_191),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_189),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_233),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_214),
.A2(n_169),
.B(n_167),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_218),
.B(n_225),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_176),
.B(n_180),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_220),
.A2(n_201),
.B(n_200),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_230),
.B(n_233),
.Y(n_288)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_170),
.B(n_163),
.C(n_201),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_273),
.A2(n_234),
.B(n_216),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_219),
.A2(n_120),
.B1(n_125),
.B2(n_102),
.Y(n_274)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_235),
.A3(n_228),
.B1(n_227),
.B2(n_218),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_245),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_292),
.B(n_265),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_289),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_235),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_285),
.B(n_253),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_288),
.B(n_275),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_296),
.Y(n_311)
);

XOR2x1_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_211),
.Y(n_289)
);

AO22x1_ASAP7_75t_SL g292 ( 
.A1(n_257),
.A2(n_233),
.B1(n_228),
.B2(n_237),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_293),
.A2(n_299),
.B1(n_273),
.B2(n_209),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_250),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_305),
.B1(n_246),
.B2(n_256),
.Y(n_323)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_247),
.A2(n_240),
.B(n_215),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_243),
.B1(n_240),
.B2(n_229),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_265),
.B1(n_271),
.B2(n_269),
.Y(n_318)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_249),
.A2(n_206),
.B1(n_207),
.B2(n_117),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_259),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_297),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_319),
.Y(n_350)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_281),
.Y(n_315)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_326),
.B1(n_332),
.B2(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_254),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_278),
.A2(n_256),
.B1(n_268),
.B2(n_274),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_320),
.A2(n_334),
.B(n_299),
.Y(n_363)
);

A2O1A1O1Ixp25_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_252),
.B(n_258),
.C(n_244),
.D(n_261),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_286),
.B(n_285),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_329),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_263),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g361 ( 
.A1(n_324),
.A2(n_330),
.B(n_331),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_258),
.C(n_252),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_328),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_268),
.B1(n_255),
.B2(n_273),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_272),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_327),
.B(n_283),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_224),
.C(n_222),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_222),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_270),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_333),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_275),
.A2(n_209),
.B(n_215),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_229),
.B1(n_270),
.B2(n_209),
.Y(n_335)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_311),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_355),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_312),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_297),
.B1(n_282),
.B2(n_298),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_344),
.A2(n_363),
.B1(n_367),
.B2(n_306),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_346),
.B(n_358),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_308),
.A2(n_299),
.B1(n_285),
.B2(n_294),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_364),
.B1(n_312),
.B2(n_326),
.Y(n_374)
);

AOI32xp33_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_288),
.A3(n_276),
.B1(n_292),
.B2(n_290),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_366),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_292),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_354),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_304),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_SL g355 ( 
.A(n_322),
.B(n_291),
.C(n_301),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_291),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_356),
.B(n_359),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_324),
.B(n_300),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_365),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_300),
.C(n_305),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_303),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_306),
.Y(n_362)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_313),
.A2(n_299),
.B1(n_302),
.B2(n_164),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_333),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_309),
.B(n_302),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_312),
.A2(n_164),
.B1(n_177),
.B2(n_166),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_310),
.C(n_319),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_378),
.C(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_330),
.Y(n_370)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

XNOR2x1_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_361),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_318),
.Y(n_372)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_337),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_377),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_374),
.A2(n_391),
.B1(n_393),
.B2(n_367),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_345),
.B(n_321),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_354),
.C(n_356),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_342),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_388),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_334),
.C(n_321),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_323),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_392),
.Y(n_397)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_315),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_390),
.A2(n_395),
.B1(n_364),
.B2(n_349),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_343),
.A2(n_335),
.B1(n_331),
.B2(n_329),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_316),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_343),
.A2(n_317),
.B1(n_307),
.B2(n_177),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_307),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_150),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_344),
.A2(n_166),
.B1(n_203),
.B2(n_154),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_396),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_400),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_393),
.B1(n_382),
.B2(n_381),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_409),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_347),
.Y(n_406)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_370),
.Y(n_408)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_408),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_341),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_411),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_355),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_386),
.Y(n_412)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_412),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_381),
.B(n_362),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_10),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_199),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_392),
.C(n_394),
.Y(n_420)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_416),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_391),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_380),
.C(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_418),
.B(n_159),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_423),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_396),
.A2(n_390),
.B1(n_395),
.B2(n_383),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_403),
.Y(n_424)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_401),
.A2(n_374),
.B(n_371),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_426),
.A2(n_399),
.B(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_0),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_430),
.A2(n_431),
.B1(n_415),
.B2(n_397),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_382),
.B1(n_132),
.B2(n_162),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_433),
.B(n_439),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_427),
.B1(n_424),
.B2(n_431),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_437),
.A2(n_438),
.B1(n_410),
.B2(n_413),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_400),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_398),
.B(n_419),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_446),
.B(n_450),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_425),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_443),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_435),
.B(n_418),
.Y(n_443)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_411),
.B(n_409),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_414),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_453),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_421),
.A2(n_405),
.B(n_397),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_451),
.A2(n_452),
.B1(n_455),
.B2(n_456),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_414),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_417),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_3),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_1),
.B(n_2),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_2),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_3),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_428),
.C(n_423),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_459),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_429),
.C(n_422),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_429),
.C(n_438),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_464),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_3),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_467),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_440),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_454),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_34),
.C(n_4),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_SL g481 ( 
.A(n_468),
.B(n_9),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_3),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_472),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_4),
.Y(n_472)
);

AOI21xp33_ASAP7_75t_L g473 ( 
.A1(n_461),
.A2(n_450),
.B(n_446),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_473),
.A2(n_476),
.B(n_479),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_470),
.B(n_447),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_484),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_469),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_444),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_456),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_458),
.A2(n_34),
.B(n_5),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_SL g489 ( 
.A(n_480),
.B(n_468),
.C(n_465),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_4),
.C(n_5),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g497 ( 
.A(n_486),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_463),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g496 ( 
.A1(n_487),
.A2(n_490),
.B(n_7),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_483),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_4),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_489),
.A2(n_478),
.B(n_482),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_480),
.A2(n_9),
.B(n_5),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_491),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_493),
.A2(n_494),
.B(n_495),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_7),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_497),
.A2(n_492),
.B(n_485),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_498),
.A2(n_7),
.B(n_8),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_499),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_501),
.A2(n_500),
.B(n_7),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_502),
.C(n_7),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_8),
.Y(n_505)
);


endmodule