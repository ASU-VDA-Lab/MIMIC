module fake_netlist_5_811_n_779 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_779);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_779;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_666;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_401;
wire n_187;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_69),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_18),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_42),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_65),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_44),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_103),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_53),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_21),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_24),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_59),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_3),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_79),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_41),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_67),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_45),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_70),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_16),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_25),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_47),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_26),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_35),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_84),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_143),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_34),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_40),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_38),
.B(n_5),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_63),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_96),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_93),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_12),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_51),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_19),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_174),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_22),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_159),
.B(n_23),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_176),
.A2(n_0),
.B(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_155),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g244 ( 
.A1(n_171),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_27),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_165),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_167),
.B(n_2),
.Y(n_252)
);

CKINVDCx11_ASAP7_75t_R g253 ( 
.A(n_179),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_253),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_169),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g268 ( 
.A(n_233),
.B(n_185),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_217),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_249),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_249),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_251),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_217),
.Y(n_281)
);

AO21x2_ASAP7_75t_L g282 ( 
.A1(n_231),
.A2(n_197),
.B(n_184),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_216),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_R g286 ( 
.A(n_234),
.B(n_170),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_254),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_254),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_252),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_254),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_4),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_213),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_223),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

CKINVDCx11_ASAP7_75t_R g298 ( 
.A(n_213),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_213),
.B(n_220),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_223),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_220),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_220),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_235),
.C(n_228),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_280),
.B(n_231),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_231),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_218),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_230),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_173),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_R g316 ( 
.A(n_267),
.B(n_188),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_261),
.B(n_202),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_234),
.B1(n_244),
.B2(n_245),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_282),
.A2(n_234),
.B1(n_244),
.B2(n_245),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_256),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_218),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_230),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_276),
.B(n_175),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_181),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_270),
.B(n_203),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_182),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_214),
.Y(n_330)
);

NOR2x1p5_ASAP7_75t_L g331 ( 
.A(n_255),
.B(n_186),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_214),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_268),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_218),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_264),
.B(n_187),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_259),
.B(n_218),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_271),
.B(n_247),
.C(n_207),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_293),
.B(n_195),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_263),
.B(n_221),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_221),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_291),
.B(n_198),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_283),
.B(n_221),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_221),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_300),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_291),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_287),
.B(n_222),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_250),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_258),
.B(n_212),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_222),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_258),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_257),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_260),
.B(n_222),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_260),
.B(n_222),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_262),
.B(n_199),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_286),
.B(n_200),
.C(n_201),
.Y(n_362)
);

NOR3xp33_ASAP7_75t_L g363 ( 
.A(n_262),
.B(n_205),
.C(n_206),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_272),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_272),
.B(n_209),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_281),
.B(n_229),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_281),
.B(n_229),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_267),
.B(n_248),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

BUFx12f_ASAP7_75t_SL g370 ( 
.A(n_312),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_364),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

AND2x6_ASAP7_75t_SL g376 ( 
.A(n_352),
.B(n_4),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_332),
.B(n_229),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_332),
.B(n_229),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_305),
.B(n_212),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_316),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_304),
.B(n_225),
.Y(n_386)
);

BUFx4f_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_28),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_310),
.A2(n_240),
.B1(n_232),
.B2(n_225),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_324),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_SL g391 ( 
.A(n_316),
.B(n_232),
.C(n_240),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_248),
.C(n_241),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_314),
.B(n_5),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_330),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_339),
.B(n_29),
.Y(n_396)
);

NOR2x2_ASAP7_75t_L g397 ( 
.A(n_318),
.B(n_6),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_368),
.B(n_362),
.Y(n_398)
);

AO22x1_ASAP7_75t_L g399 ( 
.A1(n_354),
.A2(n_248),
.B1(n_8),
.B2(n_9),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_342),
.B(n_346),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_308),
.B(n_239),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_311),
.B(n_239),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

AO21x2_ASAP7_75t_L g406 ( 
.A1(n_340),
.A2(n_90),
.B(n_152),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_239),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_239),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_334),
.B(n_241),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_318),
.B(n_241),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_307),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_327),
.A2(n_329),
.B1(n_363),
.B2(n_319),
.Y(n_413)
);

BUFx10_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_319),
.B(n_241),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_321),
.A2(n_248),
.B1(n_8),
.B2(n_9),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

BUFx4f_ASAP7_75t_L g418 ( 
.A(n_309),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_336),
.B(n_30),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_354),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_306),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_315),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_345),
.B(n_7),
.Y(n_426)
);

A2O1A1Ixp33_ASAP7_75t_L g427 ( 
.A1(n_315),
.A2(n_7),
.B(n_10),
.C(n_11),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_326),
.B(n_335),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_335),
.B(n_361),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_337),
.B(n_10),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g433 ( 
.A(n_358),
.B(n_11),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_SL g436 ( 
.A(n_367),
.B(n_12),
.C(n_13),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_341),
.B(n_13),
.Y(n_437)
);

NAND2x1_ASAP7_75t_L g438 ( 
.A(n_343),
.B(n_31),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_347),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_386),
.A2(n_383),
.B(n_418),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_413),
.A2(n_405),
.B1(n_411),
.B2(n_415),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_375),
.B(n_348),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_427),
.A2(n_365),
.B(n_338),
.C(n_331),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_14),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_437),
.A2(n_14),
.B(n_15),
.C(n_32),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_377),
.B(n_15),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_387),
.B(n_39),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_377),
.A2(n_428),
.B1(n_408),
.B2(n_392),
.Y(n_455)
);

AOI33xp33_ASAP7_75t_L g456 ( 
.A1(n_395),
.A2(n_43),
.A3(n_46),
.B1(n_49),
.B2(n_50),
.B3(n_52),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_54),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_403),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_55),
.Y(n_459)
);

O2A1O1Ixp5_ASAP7_75t_SL g460 ( 
.A1(n_378),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_423),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_418),
.A2(n_60),
.B(n_61),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_62),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_64),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

OR2x6_ASAP7_75t_SL g469 ( 
.A(n_384),
.B(n_66),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_388),
.B(n_68),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_391),
.A2(n_71),
.B(n_72),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_423),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_73),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_381),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_416),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

BUFx8_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_432),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_387),
.B(n_77),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_398),
.A2(n_78),
.B(n_80),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_81),
.Y(n_484)
);

O2A1O1Ixp33_ASAP7_75t_SL g485 ( 
.A1(n_419),
.A2(n_82),
.B(n_83),
.C(n_85),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_414),
.B(n_86),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_414),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_88),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_436),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_417),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_94),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_404),
.A2(n_409),
.B(n_410),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_493),
.A2(n_489),
.B(n_440),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_396),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_474),
.A2(n_382),
.B(n_406),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_446),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_460),
.A2(n_438),
.B(n_389),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_453),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_431),
.B(n_393),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_477),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_441),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_477),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_479),
.Y(n_507)
);

CKINVDCx8_ASAP7_75t_R g508 ( 
.A(n_473),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_487),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_443),
.A2(n_430),
.B(n_379),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_459),
.B(n_423),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_457),
.A2(n_430),
.B(n_379),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_479),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_470),
.A2(n_420),
.B(n_373),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g517 ( 
.A1(n_474),
.A2(n_399),
.B(n_434),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_439),
.A2(n_434),
.B(n_420),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_476),
.A2(n_420),
.B(n_373),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_450),
.A2(n_373),
.B(n_434),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_448),
.A2(n_95),
.B(n_97),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_447),
.A2(n_98),
.B(n_99),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_444),
.B(n_433),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_468),
.B(n_433),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_455),
.A2(n_101),
.B(n_105),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_465),
.B(n_106),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_461),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_463),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_442),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_491),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_484),
.Y(n_534)
);

BUFx2_ASAP7_75t_R g535 ( 
.A(n_469),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_484),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_488),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_520),
.A2(n_483),
.B(n_462),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_472),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_495),
.A2(n_478),
.B1(n_464),
.B2(n_454),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_497),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_504),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_514),
.A2(n_475),
.B(n_478),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_504),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_505),
.Y(n_548)
);

BUFx2_ASAP7_75t_R g549 ( 
.A(n_508),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_525),
.Y(n_550)
);

NAND2x1p5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_482),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_525),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_519),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_512),
.B(n_456),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_533),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_533),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_530),
.Y(n_557)
);

NAND2x1p5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_525),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_492),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_532),
.Y(n_561)
);

OA21x2_ASAP7_75t_L g562 ( 
.A1(n_494),
.A2(n_490),
.B(n_485),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_534),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_527),
.A2(n_490),
.B1(n_486),
.B2(n_480),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_500),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_500),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_536),
.A2(n_480),
.B1(n_376),
.B2(n_449),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_536),
.A2(n_527),
.B1(n_537),
.B2(n_526),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_500),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_494),
.A2(n_451),
.B(n_108),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_524),
.B(n_107),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_506),
.Y(n_573)
);

INVx11_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_502),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_537),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_576)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_524),
.A2(n_511),
.B(n_510),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_532),
.Y(n_578)
);

NAND2x1p5_ASAP7_75t_L g579 ( 
.A(n_511),
.B(n_113),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_542),
.B(n_522),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_541),
.Y(n_581)
);

CKINVDCx14_ASAP7_75t_R g582 ( 
.A(n_545),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_554),
.B(n_517),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_R g584 ( 
.A(n_545),
.B(n_529),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_543),
.B(n_531),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_539),
.B(n_515),
.Y(n_586)
);

NAND2x1_ASAP7_75t_L g587 ( 
.A(n_550),
.B(n_502),
.Y(n_587)
);

NOR2x1_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_506),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_502),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_R g590 ( 
.A(n_573),
.B(n_522),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_554),
.B(n_496),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_R g592 ( 
.A(n_563),
.B(n_535),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_539),
.B(n_515),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_560),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_574),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_507),
.Y(n_596)
);

AO31x2_ASAP7_75t_L g597 ( 
.A1(n_577),
.A2(n_516),
.A3(n_528),
.B(n_496),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_574),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_507),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_555),
.B(n_507),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_SL g601 ( 
.A1(n_559),
.A2(n_528),
.B1(n_523),
.B2(n_496),
.Y(n_601)
);

NOR2x1_ASAP7_75t_SL g602 ( 
.A(n_559),
.B(n_518),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_R g603 ( 
.A(n_560),
.B(n_115),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_567),
.A2(n_528),
.B1(n_523),
.B2(n_518),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_540),
.A2(n_523),
.B1(n_501),
.B2(n_518),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_546),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_549),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_555),
.B(n_553),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_560),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_556),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_R g611 ( 
.A(n_550),
.B(n_520),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_553),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_560),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_560),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_551),
.B(n_521),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_548),
.B(n_501),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_564),
.A2(n_498),
.B1(n_521),
.B2(n_119),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_557),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_565),
.B(n_566),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_576),
.B(n_116),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_544),
.B(n_498),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_569),
.B(n_118),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_550),
.B(n_120),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_R g625 ( 
.A(n_552),
.B(n_121),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_575),
.B(n_124),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_578),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_551),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_SL g629 ( 
.A(n_552),
.B(n_128),
.Y(n_629)
);

NOR2x1_ASAP7_75t_L g630 ( 
.A(n_588),
.B(n_552),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_591),
.B(n_572),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_591),
.B(n_572),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_608),
.B(n_616),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_612),
.B(n_561),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_619),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_581),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_618),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_589),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_579),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_583),
.B(n_571),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_606),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_620),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_627),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_600),
.B(n_561),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_602),
.B(n_579),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_615),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_593),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_590),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_579),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_586),
.B(n_551),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_615),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_571),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_585),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_615),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_601),
.B(n_562),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_597),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_597),
.A2(n_562),
.A3(n_570),
.B(n_571),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_597),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_596),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_582),
.B(n_561),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_609),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_580),
.B(n_558),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_604),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_580),
.B(n_558),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_570),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_631),
.B(n_605),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_631),
.B(n_562),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_666),
.A2(n_628),
.B(n_668),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_632),
.B(n_571),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_632),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_654),
.B(n_607),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_636),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_638),
.B(n_614),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_648),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_633),
.B(n_570),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_652),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_649),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_643),
.B(n_613),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_651),
.B(n_603),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_664),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_633),
.B(n_617),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_637),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_639),
.B(n_594),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_643),
.B(n_607),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_647),
.Y(n_690)
);

NAND4xp25_ASAP7_75t_L g691 ( 
.A(n_642),
.B(n_584),
.C(n_592),
.D(n_625),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_639),
.B(n_594),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_647),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_650),
.B(n_626),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_650),
.B(n_623),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_635),
.B(n_624),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_644),
.B(n_598),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_682),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_688),
.B(n_655),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_684),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_682),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_675),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_678),
.B(n_655),
.Y(n_703)
);

AND3x1_ASAP7_75t_L g704 ( 
.A(n_674),
.B(n_663),
.C(n_646),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_673),
.B(n_653),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_690),
.B(n_646),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_678),
.B(n_656),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_677),
.B(n_644),
.Y(n_708)
);

NAND4xp25_ASAP7_75t_L g709 ( 
.A(n_691),
.B(n_640),
.C(n_653),
.D(n_662),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_688),
.B(n_640),
.Y(n_710)
);

NAND4xp25_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_661),
.C(n_665),
.D(n_667),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_669),
.B(n_656),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_690),
.B(n_693),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_684),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_669),
.B(n_658),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_673),
.B(n_658),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_670),
.B(n_658),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_680),
.B(n_645),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_670),
.B(n_658),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_698),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_713),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_713),
.Y(n_722)
);

OAI32xp33_ASAP7_75t_L g723 ( 
.A1(n_709),
.A2(n_696),
.A3(n_676),
.B1(n_693),
.B2(n_672),
.Y(n_723)
);

XOR2xp5_ASAP7_75t_L g724 ( 
.A(n_711),
.B(n_595),
.Y(n_724)
);

OR3x2_ASAP7_75t_L g725 ( 
.A(n_705),
.B(n_672),
.C(n_687),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_697),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_700),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_704),
.A2(n_683),
.B1(n_671),
.B2(n_685),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_718),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_706),
.A2(n_685),
.B1(n_712),
.B2(n_694),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_701),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_728),
.A2(n_714),
.B1(n_681),
.B2(n_708),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_720),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_725),
.A2(n_715),
.B1(n_712),
.B2(n_706),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_L g735 ( 
.A1(n_723),
.A2(n_724),
.B(n_726),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_731),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_733),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_736),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_734),
.B(n_727),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_732),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_737),
.Y(n_741)
);

NOR3xp33_ASAP7_75t_L g742 ( 
.A(n_740),
.B(n_735),
.C(n_729),
.Y(n_742)
);

OAI21xp5_ASAP7_75t_SL g743 ( 
.A1(n_739),
.A2(n_730),
.B(n_727),
.Y(n_743)
);

NAND4xp25_ASAP7_75t_L g744 ( 
.A(n_738),
.B(n_715),
.C(n_692),
.D(n_694),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_743),
.A2(n_714),
.B(n_721),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_629),
.B(n_722),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_741),
.A2(n_744),
.B1(n_706),
.B2(n_695),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_745),
.A2(n_702),
.B(n_630),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_747),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_746),
.A2(n_692),
.B1(n_695),
.B2(n_716),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_SL g751 ( 
.A(n_745),
.B(n_699),
.C(n_703),
.Y(n_751)
);

NOR2x1_ASAP7_75t_L g752 ( 
.A(n_751),
.B(n_675),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_749),
.B(n_713),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_750),
.B(n_679),
.Y(n_754)
);

NOR2x1_ASAP7_75t_L g755 ( 
.A(n_748),
.B(n_679),
.Y(n_755)
);

INVxp33_ASAP7_75t_L g756 ( 
.A(n_749),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_753),
.B(n_538),
.C(n_690),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_756),
.A2(n_660),
.B(n_687),
.Y(n_758)
);

OAI221xp5_ASAP7_75t_L g759 ( 
.A1(n_755),
.A2(n_686),
.B1(n_660),
.B2(n_703),
.C(n_716),
.Y(n_759)
);

AOI221x1_ASAP7_75t_L g760 ( 
.A1(n_754),
.A2(n_686),
.B1(n_657),
.B2(n_659),
.C(n_634),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_752),
.B(n_538),
.C(n_710),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_753),
.B(n_707),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_129),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_758),
.A2(n_634),
.B(n_645),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_760),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_765),
.A2(n_761),
.B1(n_757),
.B2(n_719),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_766),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_763),
.A2(n_645),
.B1(n_717),
.B2(n_719),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_764),
.A2(n_717),
.B1(n_707),
.B2(n_659),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_769),
.B1(n_767),
.B2(n_770),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_768),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_634),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_772),
.A2(n_657),
.B1(n_135),
.B2(n_136),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_774),
.Y(n_775)
);

AOI21xp33_ASAP7_75t_SL g776 ( 
.A1(n_775),
.A2(n_771),
.B(n_773),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_776),
.A2(n_611),
.B1(n_138),
.B2(n_139),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_777),
.A2(n_134),
.B1(n_140),
.B2(n_142),
.C(n_144),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_779)
);


endmodule