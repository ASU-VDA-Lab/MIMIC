module fake_jpeg_15382_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_9),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_29),
.B(n_31),
.C(n_25),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_32),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_59),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_32),
.B(n_22),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_31),
.B(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_33),
.B1(n_34),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_79),
.B(n_23),
.C(n_24),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_34),
.B1(n_33),
.B2(n_42),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_35),
.B(n_20),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_87),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_45),
.B1(n_44),
.B2(n_36),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_93),
.B1(n_97),
.B2(n_50),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_41),
.B(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_59),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_36),
.B1(n_45),
.B2(n_44),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_19),
.C(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_95),
.B(n_19),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_41),
.B1(n_43),
.B2(n_40),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_43),
.B1(n_40),
.B2(n_38),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_20),
.B1(n_35),
.B2(n_2),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_43),
.B1(n_40),
.B2(n_38),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_117),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_59),
.B(n_50),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_115),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_88),
.B1(n_93),
.B2(n_82),
.Y(n_145)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_88),
.B1(n_96),
.B2(n_90),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_26),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_120),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_19),
.B(n_1),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_51),
.B1(n_67),
.B2(n_43),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_75),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_51),
.B1(n_40),
.B2(n_38),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_73),
.B(n_92),
.C(n_91),
.D(n_74),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_128),
.A2(n_132),
.B(n_139),
.Y(n_177)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

AOI22x1_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_104),
.B1(n_107),
.B2(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_142),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_91),
.B(n_77),
.C(n_84),
.D(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_72),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_96),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_72),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_110),
.B1(n_125),
.B2(n_107),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_54),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_19),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_126),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_155),
.C(n_99),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_19),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_176),
.B1(n_181),
.B2(n_136),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_119),
.B(n_117),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_160),
.B(n_166),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_167),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_107),
.B(n_121),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_99),
.B1(n_107),
.B2(n_115),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_179),
.B1(n_186),
.B2(n_26),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_184),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_88),
.B(n_105),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_168),
.B(n_0),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_102),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_172),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_16),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_108),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_72),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_188),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_146),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_126),
.B(n_24),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_180),
.B(n_187),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_38),
.B1(n_69),
.B2(n_54),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_143),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_69),
.B1(n_54),
.B2(n_53),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_149),
.Y(n_191)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_26),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_35),
.B1(n_20),
.B2(n_38),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_53),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_193),
.B1(n_212),
.B2(n_214),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_128),
.B1(n_151),
.B2(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_148),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_18),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_180),
.B1(n_161),
.B2(n_158),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_187),
.B(n_177),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_129),
.Y(n_205)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_53),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_216),
.Y(n_217)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_182),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_35),
.B1(n_23),
.B2(n_26),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_17),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_184),
.C(n_178),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_23),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_176),
.B1(n_180),
.B2(n_161),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_235),
.B1(n_238),
.B2(n_208),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_228),
.C(n_233),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_166),
.C(n_177),
.Y(n_228)
);

AOI21x1_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_161),
.B(n_170),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_232),
.B(n_237),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_234),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_179),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_181),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_157),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_173),
.B1(n_167),
.B2(n_171),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_163),
.B(n_183),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_26),
.C(n_24),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_17),
.C(n_18),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_189),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_192),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_231),
.C(n_239),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_210),
.B1(n_200),
.B2(n_209),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_248),
.A2(n_261),
.B1(n_264),
.B2(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_222),
.B(n_206),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_258),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_203),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_217),
.B(n_240),
.C(n_226),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_236),
.B1(n_221),
.B2(n_232),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_263),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_223),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_221),
.A2(n_203),
.B1(n_212),
.B2(n_201),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_216),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_228),
.B(n_201),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_261),
.A2(n_235),
.B(n_238),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_278),
.B(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_283),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_237),
.B(n_241),
.C(n_217),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_264),
.B(n_244),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_266),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_17),
.C(n_18),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_254),
.C(n_259),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_256),
.A2(n_1),
.B(n_2),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_2),
.B(n_3),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_294),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_298),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_257),
.B(n_255),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_293),
.B(n_10),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_273),
.B1(n_280),
.B2(n_283),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_292),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_282),
.Y(n_292)
);

OAI321xp33_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_255),
.A3(n_245),
.B1(n_252),
.B2(n_246),
.C(n_259),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_252),
.C(n_18),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_18),
.C(n_5),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_11),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_303),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_273),
.B1(n_279),
.B2(n_277),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_304),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_278),
.B1(n_12),
.B2(n_6),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_308),
.C(n_12),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_310),
.B(n_7),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_284),
.B1(n_295),
.B2(n_298),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_10),
.B(n_15),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_4),
.Y(n_314)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_12),
.B(n_15),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_317),
.B1(n_319),
.B2(n_321),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_9),
.B(n_14),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_6),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_320),
.B(n_16),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_325),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_304),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_299),
.B1(n_308),
.B2(n_311),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_13),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_329),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_318),
.B(n_14),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_328),
.B(n_322),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_327),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_335),
.A3(n_332),
.B1(n_326),
.B2(n_333),
.C1(n_16),
.C2(n_4),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_4),
.B(n_5),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_5),
.Y(n_338)
);


endmodule