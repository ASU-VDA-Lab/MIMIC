module fake_jpeg_22456_n_58 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_36;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_0),
.B(n_25),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_27),
.B(n_33),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_41),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_43),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_30),
.B1(n_4),
.B2(n_6),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_47),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_41),
.B1(n_11),
.B2(n_12),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_8),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_13),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_52),
.CI(n_50),
.CON(n_53),
.SN(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_16),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_17),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_19),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_20),
.C(n_22),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_24),
.Y(n_58)
);


endmodule