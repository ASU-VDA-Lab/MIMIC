module real_aes_11149_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_397;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g621 ( .A(n_0), .B(n_204), .Y(n_621) );
INVx1_ASAP7_75t_L g181 ( .A(n_1), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_2), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_3), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_4), .B(n_222), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_5), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_6), .B(n_591), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_7), .B(n_147), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_8), .Y(n_617) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g120 ( .A(n_9), .B(n_88), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_10), .B(n_165), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_11), .B(n_151), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_12), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_13), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_14), .B(n_165), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_15), .B(n_168), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_16), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_17), .B(n_192), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_18), .B(n_165), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_19), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_20), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_21), .B(n_151), .Y(n_267) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_22), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_23), .B(n_147), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_24), .B(n_168), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_25), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_26), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_27), .B(n_192), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_28), .B(n_168), .Y(n_561) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_29), .Y(n_149) );
OAI21xp33_ASAP7_75t_L g244 ( .A1(n_30), .A2(n_154), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_31), .B(n_151), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_32), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_33), .B(n_546), .Y(n_557) );
NAND2xp33_ASAP7_75t_SL g575 ( .A(n_34), .B(n_190), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_35), .B(n_151), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_36), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_37), .B(n_172), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_38), .B(n_223), .Y(n_548) );
INVx1_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
OAI21x1_ASAP7_75t_L g160 ( .A1(n_40), .A2(n_70), .B(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_41), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_42), .B(n_151), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_43), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_44), .B(n_172), .Y(n_607) );
AND2x6_ASAP7_75t_L g174 ( .A(n_45), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_46), .B(n_569), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_47), .A2(n_84), .B1(n_222), .B2(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_48), .B(n_569), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_49), .B(n_192), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_50), .B(n_235), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_51), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_52), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_53), .Y(n_224) );
INVx1_ASAP7_75t_L g175 ( .A(n_54), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_55), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_56), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_57), .B(n_247), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_58), .B(n_247), .Y(n_264) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_59), .B(n_190), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_60), .B(n_172), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_61), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_62), .B(n_235), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_63), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g108 ( .A(n_64), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g193 ( .A(n_65), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g131 ( .A1(n_66), .A2(n_132), .B1(n_523), .B2(n_524), .Y(n_131) );
INVx1_ASAP7_75t_L g523 ( .A(n_66), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_66), .A2(n_523), .B1(n_529), .B2(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_67), .B(n_168), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_68), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_69), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_71), .B(n_151), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_72), .B(n_165), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_73), .B(n_192), .Y(n_603) );
INVx1_ASAP7_75t_L g184 ( .A(n_74), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_75), .B(n_172), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_76), .Y(n_170) );
BUFx10_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
INVx1_ASAP7_75t_L g157 ( .A(n_78), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_79), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_80), .B(n_165), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_81), .B(n_151), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_82), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_83), .B(n_263), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_85), .B(n_235), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_86), .B(n_165), .Y(n_602) );
INVx1_ASAP7_75t_L g195 ( .A(n_87), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_88), .B(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
INVx1_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g117 ( .A(n_90), .B(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_90), .B(n_119), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_91), .B(n_189), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_92), .B(n_546), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_93), .A2(n_529), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_93), .Y(n_895) );
INVx1_ASAP7_75t_L g109 ( .A(n_94), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_95), .B(n_147), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_96), .B(n_242), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_97), .Y(n_589) );
NAND2xp33_ASAP7_75t_L g289 ( .A(n_98), .B(n_235), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_112), .B(n_899), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx11_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx6_ASAP7_75t_SL g902 ( .A(n_103), .Y(n_902) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .C(n_111), .Y(n_106) );
INVx4_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g119 ( .A(n_110), .B(n_120), .Y(n_119) );
OR2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_121), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI21xp5_ASAP7_75t_SL g892 ( .A1(n_114), .A2(n_893), .B(n_896), .Y(n_892) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx5_ASAP7_75t_L g898 ( .A(n_116), .Y(n_898) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g129 ( .A(n_118), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g881 ( .A(n_118), .B(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_889), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_131), .B(n_527), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
AND2x6_ASAP7_75t_SL g880 ( .A(n_126), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx6_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_SL g887 ( .A(n_128), .Y(n_887) );
BUFx12f_ASAP7_75t_L g891 ( .A(n_128), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_130), .Y(n_882) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g526 ( .A(n_134), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_135), .B(n_412), .Y(n_134) );
AND4x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_349), .C(n_386), .D(n_406), .Y(n_135) );
NOR2xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_319), .Y(n_136) );
OAI21xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_252), .B(n_283), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_197), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_177), .Y(n_140) );
INVx2_ASAP7_75t_L g342 ( .A(n_141), .Y(n_342) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g301 ( .A(n_142), .B(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g315 ( .A(n_143), .Y(n_315) );
INVx1_ASAP7_75t_L g334 ( .A(n_143), .Y(n_334) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_162), .B(n_171), .Y(n_143) );
AO21x1_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_153), .B(n_156), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B1(n_150), .B2(n_152), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_147), .A2(n_220), .B(n_627), .C(n_628), .Y(n_626) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g629 ( .A(n_148), .Y(n_629) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_149), .Y(n_151) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx2_ASAP7_75t_L g223 ( .A(n_149), .Y(n_223) );
INVx2_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g276 ( .A(n_151), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_151), .A2(n_223), .B1(n_616), .B2(n_617), .Y(n_615) );
AOI21x1_ASAP7_75t_L g162 ( .A1(n_153), .A2(n_163), .B(n_166), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_187), .B(n_194), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_154), .Y(n_153) );
BUFx2_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_154), .B(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_154), .A2(n_241), .B1(n_244), .B2(n_246), .Y(n_240) );
INVx3_ASAP7_75t_L g277 ( .A(n_154), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_154), .A2(n_619), .B(n_620), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_154), .A2(n_631), .B(n_632), .Y(n_630) );
BUFx12f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx5_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
INVx5_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
INVxp67_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
INVx3_ASAP7_75t_L g172 ( .A(n_158), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_158), .B(n_195), .Y(n_194) );
AOI21xp33_ASAP7_75t_L g196 ( .A1(n_158), .A2(n_174), .B(n_194), .Y(n_196) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g236 ( .A(n_160), .Y(n_236) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx5_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_170), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_168), .B(n_184), .Y(n_183) );
INVxp67_ASAP7_75t_L g296 ( .A(n_168), .Y(n_296) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
INVx2_ASAP7_75t_L g546 ( .A(n_169), .Y(n_546) );
INVx2_ASAP7_75t_L g586 ( .A(n_169), .Y(n_586) );
INVx2_ASAP7_75t_L g591 ( .A(n_169), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_176), .Y(n_171) );
INVx2_ASAP7_75t_SL g214 ( .A(n_173), .Y(n_214) );
INVx8_ASAP7_75t_L g248 ( .A(n_173), .Y(n_248) );
INVx8_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g228 ( .A(n_174), .Y(n_228) );
INVx1_ASAP7_75t_L g300 ( .A(n_174), .Y(n_300) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_174), .A2(n_601), .B(n_604), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_174), .A2(n_213), .B(n_615), .C(n_618), .Y(n_614) );
OAI21x1_ASAP7_75t_SL g625 ( .A1(n_174), .A2(n_626), .B(n_630), .Y(n_625) );
INVx2_ASAP7_75t_L g307 ( .A(n_177), .Y(n_307) );
AND2x2_ASAP7_75t_L g329 ( .A(n_177), .B(n_305), .Y(n_329) );
AND2x2_ASAP7_75t_L g395 ( .A(n_177), .B(n_201), .Y(n_395) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g312 ( .A(n_178), .Y(n_312) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_186), .B(n_196), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B(n_185), .Y(n_179) );
NOR2x1_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g243 ( .A(n_190), .Y(n_243) );
INVx2_ASAP7_75t_L g245 ( .A(n_190), .Y(n_245) );
INVx2_ASAP7_75t_L g247 ( .A(n_190), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_192), .A2(n_222), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI221xp5_ASAP7_75t_SL g414 ( .A1(n_197), .A2(n_415), .B1(n_418), .B2(n_422), .C(n_424), .Y(n_414) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp33_ASAP7_75t_R g397 ( .A1(n_198), .A2(n_398), .B(n_402), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_198), .A2(n_425), .B(n_427), .Y(n_424) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_216), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_199), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g436 ( .A(n_199), .B(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_199), .A2(n_370), .B1(n_442), .B2(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g304 ( .A(n_201), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_201), .B(n_307), .Y(n_339) );
AND2x2_ASAP7_75t_L g430 ( .A(n_201), .B(n_238), .Y(n_430) );
AND2x2_ASAP7_75t_L g457 ( .A(n_201), .B(n_218), .Y(n_457) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx3_ASAP7_75t_L g328 ( .A(n_202), .Y(n_328) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B(n_215), .Y(n_202) );
OAI21x1_ASAP7_75t_SL g271 ( .A1(n_203), .A2(n_272), .B(n_282), .Y(n_271) );
OAI21x1_ASAP7_75t_L g641 ( .A1(n_203), .A2(n_642), .B(n_650), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_203), .A2(n_642), .B(n_650), .Y(n_665) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_204), .B(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
OAI21x1_ASAP7_75t_L g624 ( .A1(n_204), .A2(n_625), .B(n_633), .Y(n_624) );
OAI21x1_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_210), .B(n_214), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .Y(n_206) );
INVx2_ASAP7_75t_SL g213 ( .A(n_209), .Y(n_213) );
CKINVDCx6p67_ASAP7_75t_R g265 ( .A(n_209), .Y(n_265) );
INVx2_ASAP7_75t_SL g298 ( .A(n_209), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_209), .A2(n_557), .B(n_558), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_209), .A2(n_232), .B(n_572), .C(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_209), .A2(n_644), .B(n_645), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_213), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_213), .A2(n_575), .B(n_576), .Y(n_574) );
AOI21x1_ASAP7_75t_L g646 ( .A1(n_213), .A2(n_647), .B(n_648), .Y(n_646) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_214), .A2(n_571), .B(n_574), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_214), .A2(n_584), .B(n_588), .Y(n_583) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_214), .A2(n_643), .B(n_646), .Y(n_642) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g399 ( .A(n_217), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g410 ( .A(n_217), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g485 ( .A(n_217), .B(n_395), .Y(n_485) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_237), .Y(n_217) );
INVx2_ASAP7_75t_SL g305 ( .A(n_218), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_218), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g375 ( .A(n_218), .B(n_312), .Y(n_375) );
INVx1_ASAP7_75t_L g385 ( .A(n_218), .Y(n_385) );
AND2x2_ASAP7_75t_L g431 ( .A(n_218), .B(n_401), .Y(n_431) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_218), .Y(n_478) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_229), .B(n_234), .Y(n_218) );
OAI21xp33_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_227), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_220), .A2(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g281 ( .A(n_220), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_220), .A2(n_548), .B(n_549), .Y(n_547) );
O2A1O1Ixp5_ASAP7_75t_L g588 ( .A1(n_220), .A2(n_589), .B(n_590), .C(n_592), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_220), .A2(n_602), .B(n_603), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B1(n_225), .B2(n_226), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g232 ( .A(n_223), .Y(n_232) );
INVx2_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_225), .A2(n_231), .B1(n_232), .B2(n_233), .Y(n_230) );
INVx2_ASAP7_75t_L g239 ( .A(n_235), .Y(n_239) );
NOR2x1p5_ASAP7_75t_SL g299 ( .A(n_235), .B(n_300), .Y(n_299) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_235), .A2(n_542), .B(n_550), .Y(n_541) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_235), .A2(n_555), .B(n_562), .Y(n_554) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_235), .A2(n_583), .B(n_593), .Y(n_582) );
OA21x2_ASAP7_75t_L g613 ( .A1(n_235), .A2(n_614), .B(n_621), .Y(n_613) );
BUFx5_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g251 ( .A(n_236), .Y(n_251) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_236), .Y(n_563) );
INVx1_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g338 ( .A(n_238), .Y(n_338) );
INVx2_ASAP7_75t_L g355 ( .A(n_238), .Y(n_355) );
AND2x4_ASAP7_75t_L g359 ( .A(n_238), .B(n_328), .Y(n_359) );
AND2x2_ASAP7_75t_L g396 ( .A(n_238), .B(n_385), .Y(n_396) );
AO31x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .A3(n_248), .B(n_249), .Y(n_238) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_248), .A2(n_261), .B(n_266), .Y(n_260) );
OAI21x1_ASAP7_75t_SL g272 ( .A1(n_248), .A2(n_273), .B(n_278), .Y(n_272) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_248), .A2(n_543), .B(n_547), .Y(n_542) );
OAI21x1_ASAP7_75t_L g555 ( .A1(n_248), .A2(n_556), .B(n_559), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_SL g569 ( .A(n_251), .Y(n_569) );
INVx1_ASAP7_75t_L g634 ( .A(n_251), .Y(n_634) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_253), .A2(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g378 ( .A(n_255), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_270), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_256), .B(n_288), .Y(n_364) );
AND2x2_ASAP7_75t_L g367 ( .A(n_256), .B(n_316), .Y(n_367) );
INVx2_ASAP7_75t_L g405 ( .A(n_256), .Y(n_405) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g302 ( .A(n_257), .Y(n_302) );
OAI21x1_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_260), .B(n_269), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_265), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_265), .A2(n_291), .B(n_294), .C(n_299), .Y(n_290) );
AND2x4_ASAP7_75t_L g286 ( .A(n_270), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g363 ( .A(n_270), .Y(n_363) );
AND2x2_ASAP7_75t_L g391 ( .A(n_270), .B(n_288), .Y(n_391) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
AOI21x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B(n_277), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_281), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_303), .B1(n_309), .B2(n_313), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_301), .Y(n_285) );
BUFx2_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
AND2x4_ASAP7_75t_L g380 ( .A(n_286), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g403 ( .A(n_286), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g520 ( .A(n_286), .B(n_342), .Y(n_520) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_288), .B(n_315), .Y(n_322) );
AND2x2_ASAP7_75t_L g368 ( .A(n_288), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_SL g426 ( .A(n_288), .Y(n_426) );
INVx1_ASAP7_75t_L g455 ( .A(n_288), .Y(n_455) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_297), .C(n_298), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_298), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_298), .A2(n_585), .B(n_587), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_298), .A2(n_605), .B(n_606), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_301), .A2(n_421), .B1(n_433), .B2(n_441), .C(n_445), .Y(n_432) );
INVx3_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_304), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_307), .B(n_308), .Y(n_348) );
INVx2_ASAP7_75t_L g421 ( .A(n_307), .Y(n_421) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_308), .Y(n_508) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g388 ( .A(n_311), .Y(n_388) );
INVx2_ASAP7_75t_L g401 ( .A(n_312), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_313), .A2(n_407), .B(n_409), .Y(n_406) );
AND2x4_ASAP7_75t_SL g313 ( .A(n_314), .B(n_317), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g454 ( .A(n_315), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g489 ( .A(n_315), .Y(n_489) );
AND2x4_ASAP7_75t_L g323 ( .A(n_316), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_318), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_317), .B(n_367), .Y(n_423) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g345 ( .A(n_318), .B(n_324), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_318), .B(n_369), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_325), .B1(n_330), .B2(n_335), .C(n_340), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_321), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g377 ( .A(n_322), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_323), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g341 ( .A(n_323), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_323), .B(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_323), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g351 ( .A(n_324), .Y(n_351) );
BUFx2_ASAP7_75t_L g381 ( .A(n_324), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_324), .B(n_333), .Y(n_408) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx2_ASAP7_75t_L g383 ( .A(n_327), .Y(n_383) );
AND2x2_ASAP7_75t_L g409 ( .A(n_327), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_327), .B(n_399), .Y(n_515) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g354 ( .A(n_328), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_SL g353 ( .A(n_329), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_331), .B(n_362), .Y(n_504) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_332), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g369 ( .A(n_334), .Y(n_369) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
AND2x2_ASAP7_75t_L g373 ( .A(n_336), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g510 ( .A(n_337), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g384 ( .A(n_338), .B(n_385), .Y(n_384) );
OAI31xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .A3(n_344), .B(n_346), .Y(n_340) );
OR2x2_ASAP7_75t_L g442 ( .A(n_342), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_342), .Y(n_483) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B(n_356), .C(n_379), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_350), .A2(n_387), .B1(n_389), .B2(n_392), .C(n_397), .Y(n_386) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_351), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g429 ( .A(n_352), .Y(n_429) );
AND2x2_ASAP7_75t_L g464 ( .A(n_354), .B(n_374), .Y(n_464) );
AND2x4_ASAP7_75t_SL g499 ( .A(n_354), .B(n_421), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_354), .B(n_477), .Y(n_522) );
AND2x4_ASAP7_75t_L g437 ( .A(n_355), .B(n_401), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B1(n_365), .B2(n_370), .C(n_372), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_359), .Y(n_371) );
AND2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_359), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g479 ( .A(n_359), .Y(n_479) );
AND2x4_ASAP7_75t_L g497 ( .A(n_359), .B(n_374), .Y(n_497) );
AOI211xp5_ASAP7_75t_L g503 ( .A1(n_360), .A2(n_504), .B(n_505), .C(n_507), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g438 ( .A(n_363), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_363), .B(n_489), .Y(n_517) );
OR2x2_ASAP7_75t_L g446 ( .A(n_364), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x2_ASAP7_75t_L g468 ( .A(n_368), .B(n_405), .Y(n_468) );
INVx2_ASAP7_75t_L g447 ( .A(n_369), .Y(n_447) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g506 ( .A(n_377), .B(n_405), .Y(n_506) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx2_ASAP7_75t_L g444 ( .A(n_380), .Y(n_444) );
OR2x2_ASAP7_75t_L g416 ( .A(n_381), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g466 ( .A(n_381), .Y(n_466) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g440 ( .A(n_384), .B(n_421), .Y(n_440) );
NOR2x1_ASAP7_75t_SL g393 ( .A(n_387), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g443 ( .A(n_391), .Y(n_443) );
AND2x2_ASAP7_75t_L g461 ( .A(n_391), .B(n_405), .Y(n_461) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g411 ( .A(n_400), .Y(n_411) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI32xp33_ASAP7_75t_L g480 ( .A1(n_404), .A2(n_446), .A3(n_481), .B1(n_482), .B2(n_484), .Y(n_480) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_405), .B(n_426), .Y(n_490) );
OR2x2_ASAP7_75t_L g513 ( .A(n_405), .B(n_453), .Y(n_513) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g491 ( .A(n_410), .Y(n_491) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_470), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_432), .C(n_458), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g494 ( .A(n_417), .Y(n_494) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .C(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_428), .Y(n_434) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x6_ASAP7_75t_L g473 ( .A(n_429), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g449 ( .A(n_430), .Y(n_449) );
AOI21xp33_ASAP7_75t_SL g458 ( .A1(n_430), .A2(n_459), .B(n_462), .Y(n_458) );
INVx2_ASAP7_75t_L g450 ( .A(n_431), .Y(n_450) );
OAI22xp33_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B1(n_438), .B2(n_439), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp33_ASAP7_75t_L g469 ( .A(n_437), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_437), .B(n_457), .Y(n_481) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g487 ( .A(n_443), .B(n_488), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_451), .B2(n_456), .Y(n_445) );
INVx2_ASAP7_75t_L g474 ( .A(n_447), .Y(n_474) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B1(n_467), .B2(n_469), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_463), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_492), .C(n_509), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B(n_480), .C(n_486), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_490), .B(n_491), .Y(n_486) );
INVx2_ASAP7_75t_L g502 ( .A(n_487), .Y(n_502) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI211xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_495), .B(n_500), .C(n_503), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_497), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_514), .B2(n_516), .C(n_518), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_879), .B1(n_883), .B2(n_884), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g894 ( .A(n_531), .Y(n_894) );
AND3x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_749), .C(n_827), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_701), .C(n_723), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_670), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_594), .B1(n_635), .B2(n_651), .C1(n_660), .C2(n_666), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_536), .B(n_564), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_551), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g802 ( .A(n_539), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g655 ( .A(n_540), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g699 ( .A(n_540), .Y(n_699) );
INVx1_ASAP7_75t_L g722 ( .A(n_540), .Y(n_722) );
AND2x2_ASAP7_75t_L g744 ( .A(n_540), .B(n_657), .Y(n_744) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_551), .B(n_743), .Y(n_742) );
NOR2x1_ASAP7_75t_L g805 ( .A(n_551), .B(n_806), .Y(n_805) );
OR2x2_ASAP7_75t_L g813 ( .A(n_551), .B(n_654), .Y(n_813) );
INVx2_ASAP7_75t_SL g842 ( .A(n_551), .Y(n_842) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g678 ( .A(n_552), .B(n_679), .Y(n_678) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_552), .Y(n_700) );
AND2x2_ASAP7_75t_L g861 ( .A(n_552), .B(n_768), .Y(n_861) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g690 ( .A(n_553), .Y(n_690) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_578), .Y(n_564) );
AND2x4_ASAP7_75t_L g687 ( .A(n_565), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g780 ( .A(n_565), .B(n_744), .Y(n_780) );
INVx1_ASAP7_75t_L g825 ( .A(n_565), .Y(n_825) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g728 ( .A(n_566), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_566), .B(n_579), .Y(n_757) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_567), .B(n_580), .Y(n_659) );
INVx2_ASAP7_75t_L g668 ( .A(n_567), .Y(n_668) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_567), .Y(n_777) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g698 ( .A(n_568), .B(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_568), .Y(n_803) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_577), .Y(n_568) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_569), .A2(n_600), .B(n_607), .Y(n_599) );
INVx2_ASAP7_75t_L g669 ( .A(n_578), .Y(n_669) );
INVx1_ASAP7_75t_L g873 ( .A(n_578), .Y(n_873) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g830 ( .A(n_579), .Y(n_830) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g796 ( .A(n_580), .B(n_668), .Y(n_796) );
INVx2_ASAP7_75t_L g768 ( .A(n_581), .Y(n_768) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g657 ( .A(n_582), .Y(n_657) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_608), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_595), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g636 ( .A(n_597), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g664 ( .A(n_598), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g683 ( .A(n_598), .Y(n_683) );
AND2x2_ASAP7_75t_L g695 ( .A(n_598), .B(n_622), .Y(n_695) );
AND2x2_ASAP7_75t_L g705 ( .A(n_598), .B(n_623), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_598), .Y(n_790) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g718 ( .A(n_599), .B(n_665), .Y(n_718) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x6_ASAP7_75t_L g772 ( .A(n_610), .B(n_773), .Y(n_772) );
INVxp67_ASAP7_75t_L g876 ( .A(n_610), .Y(n_876) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g765 ( .A(n_611), .B(n_718), .Y(n_765) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_622), .Y(n_611) );
INVx1_ASAP7_75t_L g637 ( .A(n_612), .Y(n_637) );
AND2x2_ASAP7_75t_L g693 ( .A(n_612), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_612), .B(n_623), .Y(n_783) );
AND2x2_ASAP7_75t_L g801 ( .A(n_612), .B(n_690), .Y(n_801) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g663 ( .A(n_613), .B(n_624), .Y(n_663) );
INVx2_ASAP7_75t_L g674 ( .A(n_613), .Y(n_674) );
AND2x2_ASAP7_75t_L g791 ( .A(n_613), .B(n_694), .Y(n_791) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_623), .Y(n_639) );
AND2x2_ASAP7_75t_L g685 ( .A(n_623), .B(n_637), .Y(n_685) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_623), .Y(n_717) );
INVx1_ASAP7_75t_L g748 ( .A(n_623), .Y(n_748) );
INVx1_ASAP7_75t_L g821 ( .A(n_623), .Y(n_821) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g649 ( .A(n_629), .Y(n_649) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
AND2x2_ASAP7_75t_L g745 ( .A(n_636), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_639), .B(n_683), .Y(n_809) );
INVxp67_ASAP7_75t_R g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g694 ( .A(n_641), .Y(n_694) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_658), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g763 ( .A1(n_653), .A2(n_764), .B(n_765), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g766 ( .A1(n_653), .A2(n_692), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g815 ( .A(n_655), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g866 ( .A(n_655), .B(n_777), .Y(n_866) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_656), .Y(n_713) );
AND2x2_ASAP7_75t_L g721 ( .A(n_656), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g739 ( .A(n_656), .Y(n_739) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g680 ( .A(n_657), .Y(n_680) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_L g714 ( .A(n_659), .Y(n_714) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI21xp33_ASAP7_75t_L g715 ( .A1(n_662), .A2(n_716), .B(n_719), .Y(n_715) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_663), .B(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g773 ( .A(n_664), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_664), .B(n_748), .Y(n_812) );
INVx1_ASAP7_75t_L g860 ( .A(n_664), .Y(n_860) );
BUFx2_ASAP7_75t_L g747 ( .A(n_665), .Y(n_747) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
OR2x2_ASAP7_75t_L g676 ( .A(n_667), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g769 ( .A(n_667), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_667), .B(n_768), .Y(n_806) );
INVx1_ASAP7_75t_L g816 ( .A(n_667), .Y(n_816) );
INVx1_ASAP7_75t_L g851 ( .A(n_667), .Y(n_851) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g764 ( .A(n_668), .B(n_729), .Y(n_764) );
AND2x4_ASAP7_75t_L g753 ( .A(n_669), .B(n_754), .Y(n_753) );
AOI21xp33_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_675), .B(n_681), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g759 ( .A(n_673), .B(n_705), .Y(n_759) );
OAI311xp33_ASAP7_75t_L g760 ( .A1(n_673), .A2(n_724), .A3(n_761), .B1(n_763), .C1(n_766), .Y(n_760) );
INVx1_ASAP7_75t_L g833 ( .A(n_673), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_673), .B(n_709), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_673), .B(n_718), .Y(n_848) );
OR2x2_ASAP7_75t_L g859 ( .A(n_673), .B(n_860), .Y(n_859) );
OR2x2_ASAP7_75t_L g863 ( .A(n_673), .B(n_864), .Y(n_863) );
INVx4_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g817 ( .A(n_674), .B(n_737), .Y(n_817) );
AND2x2_ASAP7_75t_L g835 ( .A(n_674), .B(n_695), .Y(n_835) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g726 ( .A(n_678), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_679), .B(n_722), .Y(n_850) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_680), .B(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B1(n_691), .B2(n_696), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g870 ( .A(n_683), .Y(n_870) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g708 ( .A(n_685), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g854 ( .A(n_689), .Y(n_854) );
BUFx2_ASAP7_75t_L g720 ( .A(n_690), .Y(n_720) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx2_ASAP7_75t_L g707 ( .A(n_693), .Y(n_707) );
AND2x4_ASAP7_75t_L g709 ( .A(n_694), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g737 ( .A(n_694), .Y(n_737) );
AND2x2_ASAP7_75t_L g845 ( .A(n_695), .B(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_698), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g843 ( .A(n_698), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_698), .B(n_873), .Y(n_878) );
INVx1_ASAP7_75t_L g729 ( .A(n_699), .Y(n_729) );
NAND2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_715), .Y(n_701) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_708), .B(n_711), .Y(n_702) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
AND2x4_ASAP7_75t_L g736 ( .A(n_705), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g864 ( .A(n_705), .Y(n_864) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x6_ASAP7_75t_L g808 ( .A(n_707), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g734 ( .A(n_708), .Y(n_734) );
INVx1_ASAP7_75t_L g793 ( .A(n_709), .Y(n_793) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_714), .B(n_721), .Y(n_792) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g724 ( .A(n_718), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_718), .B(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
AND2x2_ASAP7_75t_L g762 ( .A(n_720), .B(n_744), .Y(n_762) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_721), .Y(n_733) );
AND2x2_ASAP7_75t_L g776 ( .A(n_721), .B(n_777), .Y(n_776) );
BUFx2_ASAP7_75t_L g754 ( .A(n_722), .Y(n_754) );
OAI211xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B(n_730), .C(n_740), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B1(n_735), .B2(n_738), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g862 ( .A1(n_735), .A2(n_863), .B(n_865), .C(n_867), .Y(n_862) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_736), .A2(n_798), .B1(n_807), .B2(n_810), .C(n_811), .Y(n_797) );
AND2x2_ASAP7_75t_L g832 ( .A(n_736), .B(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g758 ( .A(n_737), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g786 ( .A(n_737), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_739), .B(n_825), .Y(n_824) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g823 ( .A(n_742), .Y(n_823) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g795 ( .A(n_744), .B(n_796), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_745), .A2(n_802), .B(n_858), .C(n_861), .Y(n_857) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g846 ( .A(n_747), .Y(n_846) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_747), .Y(n_875) );
INVx1_ASAP7_75t_L g856 ( .A(n_748), .Y(n_856) );
AND4x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_770), .C(n_797), .D(n_814), .Y(n_749) );
O2A1O1Ixp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_755), .B(n_758), .C(n_760), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_752), .A2(n_779), .B1(n_781), .B2(n_784), .Y(n_778) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_754), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g826 ( .A(n_759), .Y(n_826) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AOI211x1_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_774), .B(n_778), .C(n_787), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_776), .Y(n_810) );
INVxp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_781), .B(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g785 ( .A(n_782), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_787) );
BUFx3_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g819 ( .A(n_789), .B(n_820), .Y(n_819) );
NAND2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_796), .A2(n_815), .B1(n_817), .B2(n_818), .C(n_822), .Y(n_814) );
OAI21xp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .B(n_804), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g838 ( .A(n_802), .Y(n_838) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_815), .B(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AOI21xp33_ASAP7_75t_SL g822 ( .A1(n_823), .A2(n_824), .B(n_826), .Y(n_822) );
NOR3xp33_ASAP7_75t_SL g827 ( .A(n_828), .B(n_847), .C(n_862), .Y(n_827) );
OAI211xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_831), .B(n_834), .C(n_844), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_830), .B(n_838), .Y(n_837) );
INVxp67_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_835), .A2(n_836), .B1(n_839), .B2(n_841), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_838), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NOR2xp67_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
AND2x2_ASAP7_75t_L g853 ( .A(n_843), .B(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_846), .B(n_856), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_852), .B2(n_855), .C(n_857), .Y(n_847) );
OR2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
INVxp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AOI22xp5_ASAP7_75t_SL g867 ( .A1(n_868), .A2(n_871), .B1(n_874), .B2(n_877), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
BUFx12f_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx4_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx6_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NOR2xp33_ASAP7_75t_SL g899 ( .A(n_900), .B(n_901), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_902), .Y(n_901) );
endmodule