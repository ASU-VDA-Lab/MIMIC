module fake_jpeg_8681_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_31),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_26),
.B1(n_32),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_20),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_76),
.B1(n_40),
.B2(n_41),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_41),
.B1(n_40),
.B2(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_41),
.B1(n_58),
.B2(n_54),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_93),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.C(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_33),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_64),
.B1(n_46),
.B2(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_57),
.C(n_61),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_107),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_97),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_36),
.B(n_21),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_117),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_110),
.B1(n_85),
.B2(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_108),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_60),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_85),
.B1(n_81),
.B2(n_36),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_41),
.B1(n_62),
.B2(n_36),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_115),
.B1(n_67),
.B2(n_93),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_66),
.A2(n_36),
.B1(n_64),
.B2(n_16),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_23),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_76),
.Y(n_143)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_75),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_144),
.B1(n_150),
.B2(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_137),
.B(n_143),
.Y(n_181)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_80),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_101),
.B1(n_113),
.B2(n_103),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_77),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_89),
.B1(n_82),
.B2(n_73),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_95),
.B(n_90),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_73),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_118),
.C(n_98),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_73),
.B1(n_83),
.B2(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_128),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_106),
.B(n_119),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_169),
.B(n_21),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_105),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_167),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_172),
.B1(n_176),
.B2(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_160),
.Y(n_202)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_179),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_18),
.B1(n_21),
.B2(n_2),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_111),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_101),
.B1(n_94),
.B2(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_135),
.B1(n_145),
.B2(n_148),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_0),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_125),
.A2(n_16),
.B1(n_31),
.B2(n_25),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_175),
.B1(n_178),
.B2(n_123),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_184),
.B(n_27),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_129),
.A2(n_23),
.B1(n_22),
.B2(n_17),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_17),
.B1(n_22),
.B2(n_33),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_137),
.B1(n_146),
.B2(n_136),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_13),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_18),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_145),
.B1(n_134),
.B2(n_18),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_22),
.B1(n_33),
.B2(n_24),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_72),
.B(n_24),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_172),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_200),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_189),
.A2(n_191),
.B(n_196),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_122),
.B1(n_29),
.B2(n_24),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_194),
.B1(n_199),
.B2(n_201),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_29),
.B1(n_97),
.B2(n_72),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_27),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_29),
.B1(n_72),
.B2(n_27),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_21),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_205),
.B(n_207),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_37),
.B(n_27),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_157),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_158),
.B1(n_159),
.B2(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_160),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_8),
.B(n_15),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_153),
.C(n_161),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_226),
.C(n_186),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_169),
.B(n_184),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_235),
.B(n_5),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_168),
.C(n_157),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_185),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_192),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_167),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_179),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_170),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_165),
.B1(n_169),
.B2(n_159),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_233),
.B1(n_237),
.B2(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_191),
.B(n_175),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_165),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_188),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_245),
.C(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_219),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_247),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_189),
.C(n_201),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_198),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_190),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_226),
.C(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_203),
.C(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_207),
.B1(n_190),
.B2(n_4),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_235),
.B1(n_223),
.B2(n_218),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_233),
.B1(n_216),
.B2(n_229),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_21),
.C(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_4),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_240),
.B(n_251),
.Y(n_267)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_232),
.B1(n_216),
.B2(n_222),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_223),
.B1(n_220),
.B2(n_7),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_244),
.B1(n_241),
.B2(n_246),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_238),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_282),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_275),
.A2(n_258),
.B1(n_268),
.B2(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_284),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_245),
.B(n_238),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_266),
.B(n_259),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_5),
.C(n_6),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_267),
.C(n_266),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_15),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_6),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_14),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_286),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_297),
.B(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_268),
.B1(n_261),
.B2(n_260),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_296),
.C(n_274),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_281),
.C(n_260),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_259),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_278),
.B(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_262),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_305),
.B(n_285),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_306),
.B(n_301),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_275),
.B(n_269),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_288),
.C(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_310),
.Y(n_314)
);

INVx11_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_311),
.B(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_308),
.C(n_309),
.Y(n_316)
);

AO221x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_314),
.B1(n_310),
.B2(n_312),
.C(n_273),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_7),
.C(n_11),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_12),
.C(n_306),
.Y(n_319)
);


endmodule