module fake_netlist_6_2225_n_2831 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2831);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2831;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_761;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g617 ( 
.A(n_132),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_360),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_0),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_134),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_587),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_258),
.Y(n_622)
);

BUFx5_ASAP7_75t_L g623 ( 
.A(n_79),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_99),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_215),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_258),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_366),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_395),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_606),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_251),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_597),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_0),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_48),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_574),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_464),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_46),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_217),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_580),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_146),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_229),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_514),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_44),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_482),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_360),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_80),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_260),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_267),
.Y(n_649)
);

BUFx5_ASAP7_75t_L g650 ( 
.A(n_354),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_428),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_118),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_244),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_246),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_225),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_403),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_460),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_412),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_498),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_86),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_544),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_566),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_179),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_613),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_77),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_556),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_356),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_543),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_478),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_193),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_459),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_189),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_549),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_215),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_24),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_71),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_475),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_551),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_149),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_73),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_139),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_281),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_413),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_419),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_462),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_602),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_433),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_264),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_435),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_478),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_462),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_167),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_367),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_338),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_431),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_567),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_535),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_235),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_13),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_581),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_483),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_269),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_90),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_446),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_256),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_357),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_569),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_392),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_511),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_600),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_189),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_196),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_471),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_410),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_60),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_486),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_573),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_205),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_287),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_34),
.Y(n_723)
);

BUFx8_ASAP7_75t_SL g724 ( 
.A(n_323),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_526),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_550),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_80),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_21),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_601),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_399),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_353),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_207),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_533),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_366),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_451),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_612),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_131),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_14),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_11),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_64),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_350),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_545),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_435),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_418),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_320),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_436),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_12),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_510),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_452),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_517),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_14),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_154),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_541),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_359),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_517),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_340),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_164),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_236),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_444),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_429),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_37),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_532),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_399),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_274),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_20),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_64),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_525),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_8),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_172),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_493),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_481),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_363),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_537),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_556),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_118),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_38),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_253),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_466),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_536),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_391),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_317),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_82),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_529),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_409),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_349),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_503),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_252),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_358),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_261),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_518),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_550),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_151),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_340),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_350),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_471),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_551),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_538),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_98),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_421),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_436),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_534),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_135),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_175),
.Y(n_803)
);

CKINVDCx14_ASAP7_75t_R g804 ( 
.A(n_220),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_7),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_546),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_337),
.Y(n_807)
);

BUFx5_ASAP7_75t_L g808 ( 
.A(n_538),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_326),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_67),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_18),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_542),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_594),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_595),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_343),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_344),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_314),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_172),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_519),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_509),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_335),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_110),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_246),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_193),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_66),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_521),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_288),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_577),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_540),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_443),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_196),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_204),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_582),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_303),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_13),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_500),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_301),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_374),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_43),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_304),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_122),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_464),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_358),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_9),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_455),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_496),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_509),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_562),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_30),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_315),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_525),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_522),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_214),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_500),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_200),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_558),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_238),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_327),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_623),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_623),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_623),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_630),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_630),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_724),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_724),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_623),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_623),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_804),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_623),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_719),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_623),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_796),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_710),
.B(n_1),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_636),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_650),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_635),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_650),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_820),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_650),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_650),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_650),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_618),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_650),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_650),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_715),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_710),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_635),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_759),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_715),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_715),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_715),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_715),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_642),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_715),
.Y(n_895)
);

CKINVDCx14_ASAP7_75t_R g896 ( 
.A(n_642),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_808),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_710),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_808),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_799),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_808),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_808),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_636),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_808),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_622),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_791),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_808),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_764),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_808),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_764),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_791),
.Y(n_911)
);

BUFx2_ASAP7_75t_SL g912 ( 
.A(n_640),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_791),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_642),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_656),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_656),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_677),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_677),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_695),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_695),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_646),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_704),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_674),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_704),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_764),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_774),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_774),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_774),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_774),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_798),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_798),
.Y(n_932)
);

CKINVDCx16_ASAP7_75t_R g933 ( 
.A(n_674),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_798),
.Y(n_934)
);

CKINVDCx16_ASAP7_75t_R g935 ( 
.A(n_674),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_798),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_826),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_826),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_625),
.Y(n_939)
);

INVxp33_ASAP7_75t_L g940 ( 
.A(n_617),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_826),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_841),
.Y(n_942)
);

BUFx2_ASAP7_75t_SL g943 ( 
.A(n_640),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_841),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_841),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_841),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_698),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_624),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_842),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_842),
.Y(n_950)
);

INVxp33_ASAP7_75t_SL g951 ( 
.A(n_634),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_842),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_842),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_626),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_698),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_627),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_626),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_848),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_628),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_944),
.B(n_945),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_934),
.Y(n_961)
);

INVx5_ASAP7_75t_L g962 ( 
.A(n_908),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_910),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_934),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_910),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_950),
.B(n_833),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_958),
.B(n_848),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_873),
.B(n_833),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_868),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_892),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_886),
.B(n_631),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_868),
.Y(n_972)
);

CKINVDCx11_ASAP7_75t_R g973 ( 
.A(n_862),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_937),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_874),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_912),
.B(n_664),
.Y(n_976)
);

AND2x2_ASAP7_75t_R g977 ( 
.A(n_896),
.B(n_857),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_874),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_892),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_937),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_876),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_870),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_952),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_942),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_908),
.B(n_898),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_912),
.B(n_633),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_863),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_863),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_906),
.B(n_707),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_952),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_942),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_908),
.B(n_717),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_943),
.B(n_633),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_903),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_911),
.B(n_729),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_953),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_874),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_874),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_943),
.B(n_621),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_903),
.B(n_662),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_953),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_915),
.B(n_707),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_864),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_870),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_874),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_915),
.B(n_686),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_893),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_916),
.B(n_697),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_882),
.B(n_856),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_917),
.B(n_919),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_925),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_926),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_913),
.B(n_638),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_893),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_920),
.B(n_701),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_927),
.Y(n_1016)
);

INVx5_ASAP7_75t_L g1017 ( 
.A(n_948),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_948),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_918),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_928),
.Y(n_1020)
);

BUFx8_ASAP7_75t_L g1021 ( 
.A(n_918),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_922),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_876),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_929),
.B(n_638),
.Y(n_1024)
);

CKINVDCx11_ASAP7_75t_R g1025 ( 
.A(n_862),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_SL g1026 ( 
.A1(n_981),
.A2(n_651),
.B1(n_679),
.B2(n_646),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_970),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1012),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_985),
.B(n_930),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1012),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_967),
.B(n_951),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_1009),
.B(n_951),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_986),
.B(n_882),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_1005),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_961),
.Y(n_1035)
);

AOI22x1_ASAP7_75t_SL g1036 ( 
.A1(n_1023),
.A2(n_679),
.B1(n_718),
.B2(n_651),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_970),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_971),
.A2(n_861),
.B(n_859),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_960),
.B(n_931),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_1019),
.B(n_894),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_961),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_985),
.B(n_932),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_994),
.B(n_900),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_960),
.B(n_936),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_994),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_970),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1019),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_979),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_979),
.Y(n_1049)
);

BUFx8_ASAP7_75t_L g1050 ( 
.A(n_972),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_993),
.A2(n_939),
.B1(n_956),
.B2(n_905),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_1005),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_964),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_972),
.B(n_793),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_998),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1019),
.B(n_914),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_979),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_1005),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_985),
.B(n_995),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_982),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_985),
.B(n_938),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_960),
.B(n_941),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_966),
.B(n_946),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1014),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_964),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_980),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1019),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_980),
.Y(n_1068)
);

AND2x6_ASAP7_75t_L g1069 ( 
.A(n_976),
.B(n_667),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_984),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_995),
.B(n_949),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_984),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1012),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1014),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_989),
.B(n_924),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_1019),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1014),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1014),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1006),
.B(n_947),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1019),
.B(n_923),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_1022),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_1007),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_966),
.B(n_866),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_1005),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_995),
.B(n_954),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_963),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_995),
.B(n_954),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_1005),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_963),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_991),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1007),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1021),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_975),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_996),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_996),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_966),
.B(n_867),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_965),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1001),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_965),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1001),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_983),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1007),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1007),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_983),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_966),
.B(n_957),
.Y(n_1106)
);

OA21x2_ASAP7_75t_L g1107 ( 
.A1(n_968),
.A2(n_871),
.B(n_869),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_990),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_989),
.B(n_922),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_999),
.B(n_905),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_990),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1007),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_976),
.B(n_667),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_974),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1043),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_1093),
.B(n_987),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1031),
.A2(n_1000),
.B1(n_1015),
.B2(n_1008),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1109),
.B(n_1022),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1080),
.B(n_1033),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1035),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_1038),
.A2(n_968),
.B(n_877),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1059),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1080),
.B(n_1022),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1041),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1041),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_1032),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1043),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1110),
.B(n_1022),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1059),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1053),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1109),
.B(n_1022),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1059),
.A2(n_968),
.B1(n_992),
.B2(n_897),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1029),
.B(n_968),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1051),
.B(n_1022),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1108),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1045),
.B(n_969),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1053),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1076),
.B(n_1106),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1029),
.B(n_1042),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1040),
.B(n_969),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_L g1142 ( 
.A(n_1069),
.B(n_856),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1065),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1065),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1107),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1108),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1060),
.B(n_982),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1029),
.B(n_1042),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1042),
.B(n_1061),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1107),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1061),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1066),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1061),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1076),
.B(n_956),
.C(n_939),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1056),
.B(n_1004),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1066),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1068),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1068),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1070),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1070),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1072),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1072),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1094),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1075),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1106),
.B(n_1021),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1107),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1106),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1075),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1091),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1069),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1091),
.Y(n_1171)
);

CKINVDCx6p67_ASAP7_75t_R g1172 ( 
.A(n_1093),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1081),
.B(n_1021),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1095),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1047),
.B(n_864),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1095),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1096),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1096),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1099),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1039),
.B(n_975),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1094),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1099),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1114),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1101),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1026),
.B(n_955),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1101),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1050),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1086),
.B(n_1002),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1027),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1027),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1086),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1055),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1037),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1044),
.B(n_975),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1062),
.B(n_997),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1094),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1084),
.A2(n_899),
.B(n_875),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1046),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1028),
.B(n_959),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1114),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1046),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1048),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1048),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1049),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1049),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1057),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1030),
.B(n_959),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1057),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1087),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1090),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1069),
.A2(n_992),
.B1(n_709),
.B2(n_720),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1073),
.B(n_978),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1086),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1088),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1098),
.B(n_933),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1088),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1100),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1102),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1105),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1111),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1069),
.A2(n_992),
.B1(n_712),
.B2(n_813),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1088),
.Y(n_1222)
);

INVx5_ASAP7_75t_L g1223 ( 
.A(n_1055),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1064),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1094),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1064),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1074),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1097),
.A2(n_1069),
.B1(n_1113),
.B2(n_1071),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1074),
.Y(n_1229)
);

NOR2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1050),
.B(n_865),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1063),
.B(n_978),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1078),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1078),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1079),
.Y(n_1234)
);

BUFx10_ASAP7_75t_L g1235 ( 
.A(n_1069),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1079),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1103),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1103),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1071),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1104),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1071),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1038),
.B(n_1002),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1104),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1112),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1094),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1113),
.Y(n_1246)
);

INVxp33_ASAP7_75t_SL g1247 ( 
.A(n_1036),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1112),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1113),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1050),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1036),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1115),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1147),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1226),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1226),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1136),
.B(n_1113),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1134),
.A2(n_1092),
.B(n_1077),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1189),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1147),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1227),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1227),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1120),
.B(n_1054),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1229),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1115),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1229),
.Y(n_1265)
);

XOR2xp5_ASAP7_75t_L g1266 ( 
.A(n_1187),
.B(n_888),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1172),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1189),
.Y(n_1268)
);

AND2x2_ASAP7_75t_SL g1269 ( 
.A(n_1185),
.B(n_935),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1232),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1123),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1232),
.Y(n_1272)
);

XNOR2xp5_ASAP7_75t_L g1273 ( 
.A(n_1230),
.B(n_888),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1234),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1234),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1190),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1128),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1128),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1172),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1198),
.Y(n_1280)
);

XOR2xp5_ASAP7_75t_L g1281 ( 
.A(n_1187),
.B(n_921),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1193),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1201),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1123),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1201),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1250),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1145),
.A2(n_1092),
.B(n_1077),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1127),
.B(n_1054),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_SL g1290 ( 
.A(n_1116),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1139),
.B(n_1054),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1208),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1208),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1151),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1140),
.A2(n_1092),
.B(n_1067),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1151),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1153),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1153),
.Y(n_1298)
);

XOR2xp5_ASAP7_75t_L g1299 ( 
.A(n_1250),
.B(n_921),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_SL g1300 ( 
.A(n_1127),
.B(n_1141),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1127),
.B(n_1054),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1198),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1202),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_1130),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1202),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1203),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1203),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1204),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_L g1309 ( 
.A(n_1154),
.B(n_987),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1204),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1155),
.B(n_872),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1205),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1119),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1205),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1206),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1206),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1136),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1146),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1188),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1139),
.B(n_878),
.Y(n_1320)
);

INVxp33_ASAP7_75t_L g1321 ( 
.A(n_1215),
.Y(n_1321)
);

XOR2xp5_ASAP7_75t_L g1322 ( 
.A(n_1118),
.B(n_865),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1146),
.Y(n_1323)
);

XOR2xp5_ASAP7_75t_L g1324 ( 
.A(n_1185),
.B(n_1247),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1224),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1224),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1233),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1233),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1188),
.B(n_889),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1236),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1199),
.B(n_988),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1236),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1130),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1119),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1217),
.B(n_1113),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1191),
.B(n_1082),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1116),
.B(n_988),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1137),
.B(n_1021),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1130),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1148),
.A2(n_1083),
.B(n_1052),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1207),
.B(n_1003),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1124),
.B(n_1003),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1174),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1116),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1216),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1163),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1174),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1176),
.Y(n_1348)
);

AND2x6_ASAP7_75t_L g1349 ( 
.A(n_1242),
.B(n_1034),
.Y(n_1349)
);

XNOR2xp5_ASAP7_75t_L g1350 ( 
.A(n_1230),
.B(n_1165),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1217),
.B(n_1209),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1176),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1177),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1177),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1178),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1178),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1184),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1184),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1186),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1186),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1239),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_SL g1362 ( 
.A(n_1170),
.B(n_718),
.Y(n_1362)
);

INVxp33_ASAP7_75t_L g1363 ( 
.A(n_1173),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1209),
.B(n_754),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1239),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1210),
.B(n_754),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1241),
.Y(n_1367)
);

XOR2xp5_ASAP7_75t_L g1368 ( 
.A(n_1247),
.B(n_1211),
.Y(n_1368)
);

XOR2xp5_ASAP7_75t_L g1369 ( 
.A(n_1221),
.B(n_973),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1210),
.B(n_940),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1241),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1149),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1216),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1218),
.B(n_1010),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1218),
.B(n_1013),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1219),
.B(n_778),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_1163),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1222),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1222),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1222),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1156),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1156),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1157),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1116),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1157),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1219),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1220),
.B(n_647),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1159),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1220),
.B(n_1013),
.Y(n_1389)
);

AND2x6_ASAP7_75t_L g1390 ( 
.A(n_1242),
.B(n_1034),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1159),
.Y(n_1391)
);

INVxp33_ASAP7_75t_SL g1392 ( 
.A(n_1251),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1167),
.B(n_1013),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1164),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1164),
.Y(n_1395)
);

NOR2xp67_ASAP7_75t_L g1396 ( 
.A(n_1135),
.B(n_1017),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1168),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1167),
.B(n_1013),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1175),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1168),
.Y(n_1400)
);

XNOR2xp5_ASAP7_75t_L g1401 ( 
.A(n_1132),
.B(n_1025),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1171),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1117),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1171),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1121),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1179),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1179),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1191),
.B(n_698),
.Y(n_1408)
);

XOR2xp5_ASAP7_75t_L g1409 ( 
.A(n_1213),
.B(n_778),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1182),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1182),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1213),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1129),
.Y(n_1413)
);

XOR2xp5_ASAP7_75t_L g1414 ( 
.A(n_1214),
.B(n_1133),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1121),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1125),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1125),
.Y(n_1417)
);

XNOR2x2_ASAP7_75t_L g1418 ( 
.A(n_1180),
.B(n_702),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1214),
.B(n_781),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1126),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1145),
.A2(n_1113),
.B(n_992),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1126),
.Y(n_1422)
);

XOR2x2_ASAP7_75t_L g1423 ( 
.A(n_1228),
.B(n_977),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1131),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1131),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1138),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1237),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1246),
.B(n_793),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1170),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1246),
.B(n_781),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1212),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1163),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1143),
.B(n_757),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1237),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1163),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1249),
.B(n_1024),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1143),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1144),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1145),
.A2(n_902),
.B(n_901),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1163),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1144),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1181),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1181),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1152),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1249),
.B(n_781),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1152),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1158),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1325),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_L g1449 ( 
.A(n_1342),
.B(n_1238),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1254),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1374),
.B(n_1313),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1423),
.A2(n_1142),
.B1(n_835),
.B2(n_847),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1351),
.B(n_1150),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1321),
.B(n_1150),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1330),
.Y(n_1455)
);

AO22x1_ASAP7_75t_L g1456 ( 
.A1(n_1311),
.A2(n_629),
.B1(n_637),
.B2(n_634),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1253),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1255),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1311),
.B(n_1166),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1372),
.A2(n_1142),
.B1(n_835),
.B2(n_784),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1334),
.B(n_1166),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1386),
.B(n_1158),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_L g1463 ( 
.A(n_1364),
.B(n_670),
.C(n_641),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1277),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_SL g1465 ( 
.A(n_1287),
.B(n_1253),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1362),
.B(n_1194),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1260),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1258),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1259),
.B(n_1160),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1268),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1362),
.B(n_1195),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1264),
.B(n_1300),
.Y(n_1472)
);

NOR2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1384),
.B(n_977),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1431),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1261),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1263),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1319),
.B(n_1238),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1370),
.B(n_1160),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1280),
.Y(n_1479)
);

CKINVDCx11_ASAP7_75t_R g1480 ( 
.A(n_1267),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1302),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1320),
.B(n_1024),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1317),
.A2(n_847),
.B1(n_853),
.B2(n_784),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1318),
.B(n_1161),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1264),
.B(n_1345),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1323),
.B(n_1161),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1412),
.B(n_1162),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1412),
.B(n_1162),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1291),
.B(n_1240),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1265),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1271),
.B(n_1169),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1329),
.B(n_1024),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1252),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1285),
.B(n_1235),
.Y(n_1494)
);

AND2x2_ASAP7_75t_SL g1495 ( 
.A(n_1269),
.B(n_1196),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1345),
.B(n_1235),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1270),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1272),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1403),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1271),
.B(n_1169),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1322),
.A2(n_853),
.B1(n_637),
.B2(n_748),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1304),
.B(n_1231),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1279),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1387),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1294),
.A2(n_815),
.B1(n_765),
.B2(n_708),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1252),
.B(n_1240),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1276),
.B(n_1243),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1274),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1364),
.B(n_1024),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_L g1510 ( 
.A(n_1432),
.B(n_1181),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1275),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1433),
.B(n_1244),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1278),
.B(n_1414),
.Y(n_1513)
);

BUFx5_ASAP7_75t_L g1514 ( 
.A(n_1349),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1405),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1426),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1345),
.B(n_1379),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1283),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1366),
.B(n_1248),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1366),
.B(n_1122),
.Y(n_1520)
);

NAND2xp33_ASAP7_75t_L g1521 ( 
.A(n_1435),
.B(n_1181),
.Y(n_1521)
);

INVx5_ASAP7_75t_L g1522 ( 
.A(n_1349),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1285),
.B(n_1181),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1326),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1278),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1296),
.A2(n_708),
.B1(n_713),
.B2(n_676),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1376),
.B(n_1409),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1291),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1282),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1284),
.B(n_1183),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1429),
.A2(n_1245),
.B1(n_1225),
.B2(n_1196),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1376),
.B(n_1183),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1408),
.B(n_1122),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1327),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1379),
.B(n_1245),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1286),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1439),
.A2(n_1245),
.B(n_1225),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1419),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1292),
.B(n_1200),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1293),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1331),
.B(n_1122),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1335),
.A2(n_1343),
.B(n_1348),
.C(n_1347),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1303),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1297),
.A2(n_713),
.B1(n_789),
.B2(n_676),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1305),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1379),
.B(n_1196),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1375),
.B(n_1200),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1285),
.B(n_1225),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1341),
.B(n_1200),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1262),
.B(n_957),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1336),
.B(n_1017),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1389),
.B(n_1011),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1306),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1298),
.B(n_1011),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1361),
.B(n_997),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1365),
.B(n_997),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1307),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1308),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1336),
.B(n_1017),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1367),
.B(n_1197),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1371),
.B(n_1197),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1418),
.B(n_748),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1430),
.B(n_736),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1401),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1445),
.B(n_814),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1398),
.B(n_1310),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1266),
.B(n_855),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1413),
.A2(n_828),
.B1(n_1018),
.B2(n_1017),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_SL g1569 ( 
.A(n_1337),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1281),
.A2(n_855),
.B1(n_643),
.B2(n_645),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1312),
.B(n_1018),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_SL g1572 ( 
.A(n_1337),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1363),
.B(n_632),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1328),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1314),
.B(n_1018),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1442),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1338),
.B(n_644),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1393),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1337),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1332),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1352),
.B(n_1018),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1399),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1344),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1353),
.Y(n_1585)
);

O2A1O1Ixp5_ASAP7_75t_L g1586 ( 
.A1(n_1256),
.A2(n_907),
.B(n_909),
.C(n_904),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1354),
.B(n_1018),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1355),
.B(n_1018),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1439),
.A2(n_1223),
.B(n_1192),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_L g1590 ( 
.A(n_1349),
.B(n_1192),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1442),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1436),
.A2(n_803),
.B1(n_789),
.B2(n_620),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1356),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1392),
.B(n_648),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1428),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1357),
.B(n_1034),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1428),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1335),
.A2(n_639),
.B(n_649),
.C(n_619),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1440),
.Y(n_1599)
);

NOR3xp33_ASAP7_75t_L g1600 ( 
.A(n_1289),
.B(n_1301),
.C(n_1309),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1289),
.B(n_653),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1346),
.A2(n_1223),
.B1(n_1192),
.B2(n_1052),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1373),
.B(n_1192),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1406),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1256),
.A2(n_655),
.B(n_659),
.C(n_652),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1301),
.B(n_654),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1358),
.B(n_1034),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1428),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1378),
.A2(n_1052),
.B1(n_1058),
.B2(n_1034),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1380),
.B(n_1223),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1359),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1407),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1410),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1411),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1333),
.B(n_1339),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1360),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1381),
.B(n_1052),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1393),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1382),
.B(n_657),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1383),
.B(n_658),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1415),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1416),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1385),
.B(n_1052),
.Y(n_1623)
);

BUFx12f_ASAP7_75t_L g1624 ( 
.A(n_1393),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1350),
.A2(n_1085),
.B1(n_1089),
.B2(n_1058),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1443),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1388),
.B(n_1058),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1421),
.A2(n_1223),
.B(n_1288),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1391),
.B(n_1058),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1394),
.B(n_1058),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1395),
.B(n_1085),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1417),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1397),
.B(n_1400),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1349),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1402),
.B(n_1085),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1404),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1346),
.A2(n_1089),
.B1(n_1085),
.B2(n_661),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1420),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1422),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1427),
.B(n_1085),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1377),
.B(n_1089),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1424),
.A2(n_666),
.B1(n_673),
.B2(n_665),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1451),
.A2(n_1377),
.B1(n_1421),
.B2(n_1434),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1474),
.B(n_1273),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1527),
.B(n_1299),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1459),
.B(n_1425),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1589),
.A2(n_1288),
.B(n_1257),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1459),
.B(n_1550),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1537),
.A2(n_1257),
.B(n_1340),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1586),
.A2(n_1295),
.B(n_1340),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1628),
.A2(n_1396),
.B(n_1295),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1478),
.B(n_1437),
.Y(n_1652)
);

NOR2xp67_ASAP7_75t_L g1653 ( 
.A(n_1583),
.B(n_1504),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1480),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1465),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1450),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1590),
.A2(n_1441),
.B(n_1438),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1482),
.B(n_1444),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1586),
.A2(n_1447),
.B(n_1446),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1509),
.B(n_1390),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1492),
.B(n_1454),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1522),
.B(n_1089),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1520),
.A2(n_1390),
.B(n_877),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1454),
.B(n_1390),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1562),
.A2(n_678),
.B(n_682),
.C(n_675),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1598),
.A2(n_1390),
.B(n_879),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1599),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1605),
.A2(n_879),
.B(n_860),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1510),
.A2(n_1083),
.B(n_1089),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1513),
.B(n_1368),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1466),
.B(n_1324),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1513),
.A2(n_1369),
.B1(n_1290),
.B2(n_663),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1458),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1495),
.A2(n_1578),
.B1(n_1606),
.B2(n_1601),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1521),
.A2(n_1083),
.B(n_998),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1457),
.B(n_1290),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1464),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1549),
.A2(n_668),
.B1(n_669),
.B2(n_660),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_L g1679 ( 
.A(n_1514),
.B(n_671),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1493),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1549),
.A2(n_680),
.B1(n_681),
.B2(n_672),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1472),
.B(n_1460),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1466),
.B(n_688),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1471),
.B(n_696),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1533),
.A2(n_880),
.B(n_860),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1604),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1471),
.B(n_699),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1519),
.B(n_1538),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_L g1689 ( 
.A(n_1463),
.B(n_737),
.C(n_714),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1602),
.A2(n_1083),
.B(n_998),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1532),
.B(n_723),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1532),
.A2(n_883),
.B(n_881),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1502),
.A2(n_998),
.B(n_1055),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1495),
.B(n_683),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1612),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1467),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1634),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1601),
.B(n_727),
.Y(n_1699)
);

INVxp33_ASAP7_75t_SL g1700 ( 
.A(n_1503),
.Y(n_1700)
);

INVx4_ASAP7_75t_SL g1701 ( 
.A(n_1634),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1472),
.B(n_684),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1475),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1613),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1606),
.B(n_731),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1452),
.A2(n_687),
.B(n_685),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1614),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1621),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1493),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1547),
.A2(n_884),
.B(n_883),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1594),
.A2(n_690),
.B1(n_691),
.B2(n_689),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1541),
.A2(n_693),
.B1(n_694),
.B2(n_692),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1453),
.A2(n_887),
.B(n_885),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1542),
.A2(n_887),
.B(n_885),
.Y(n_1714)
);

CKINVDCx8_ASAP7_75t_R g1715 ( 
.A(n_1599),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1552),
.A2(n_891),
.B(n_890),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1622),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1591),
.B(n_738),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1452),
.A2(n_742),
.B1(n_747),
.B2(n_741),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1619),
.B(n_749),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1542),
.A2(n_891),
.B(n_890),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1476),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1460),
.B(n_700),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1522),
.A2(n_895),
.B(n_962),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1494),
.A2(n_895),
.B(n_854),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1620),
.B(n_703),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1632),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1594),
.B(n_705),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1522),
.A2(n_962),
.B(n_974),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1522),
.A2(n_1641),
.B(n_1500),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1494),
.A2(n_852),
.B(n_752),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1449),
.A2(n_755),
.B(n_756),
.C(n_751),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1491),
.A2(n_962),
.B(n_974),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1563),
.A2(n_962),
.B(n_974),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1569),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1573),
.B(n_706),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1620),
.B(n_769),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1490),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1497),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1506),
.B(n_777),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1573),
.B(n_711),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1498),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1508),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1560),
.A2(n_792),
.B(n_783),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1506),
.B(n_1565),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1511),
.B(n_800),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1505),
.A2(n_802),
.B(n_805),
.C(n_801),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1531),
.A2(n_962),
.B(n_1016),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1566),
.A2(n_962),
.B(n_1016),
.Y(n_1749)
);

O2A1O1Ixp5_ASAP7_75t_L g1750 ( 
.A1(n_1496),
.A2(n_817),
.B(n_818),
.C(n_812),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1580),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1600),
.A2(n_721),
.B1(n_722),
.B2(n_716),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1599),
.Y(n_1753)
);

AO21x1_ASAP7_75t_L g1754 ( 
.A1(n_1600),
.A2(n_824),
.B(n_821),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1528),
.B(n_839),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1529),
.B(n_845),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1461),
.A2(n_726),
.B(n_725),
.Y(n_1757)
);

AO21x1_ASAP7_75t_L g1758 ( 
.A1(n_1561),
.A2(n_3),
.B(n_2),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1638),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1639),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1489),
.B(n_728),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1525),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1618),
.A2(n_732),
.B(n_733),
.C(n_730),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1591),
.B(n_1016),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1524),
.Y(n_1765)
);

AOI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1603),
.A2(n_1020),
.B(n_560),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1567),
.B(n_1469),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1633),
.A2(n_735),
.B1(n_739),
.B2(n_734),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1518),
.A2(n_1020),
.B(n_561),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1518),
.A2(n_1020),
.B(n_563),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1489),
.B(n_559),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1579),
.A2(n_743),
.B1(n_744),
.B2(n_740),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1536),
.B(n_745),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1540),
.B(n_746),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1585),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1534),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1523),
.A2(n_570),
.B(n_568),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1525),
.B(n_750),
.Y(n_1778)
);

CKINVDCx6p67_ASAP7_75t_R g1779 ( 
.A(n_1569),
.Y(n_1779)
);

NOR3xp33_ASAP7_75t_L g1780 ( 
.A(n_1456),
.B(n_758),
.C(n_753),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1501),
.B(n_760),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_L g1782 ( 
.A(n_1514),
.B(n_761),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1523),
.A2(n_572),
.B(n_571),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1597),
.B(n_762),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1570),
.B(n_763),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1599),
.Y(n_1786)
);

INVx5_ASAP7_75t_L g1787 ( 
.A(n_1634),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1584),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1473),
.A2(n_767),
.B1(n_768),
.B2(n_766),
.Y(n_1789)
);

AND2x2_ASAP7_75t_SL g1790 ( 
.A(n_1483),
.B(n_1),
.Y(n_1790)
);

INVx4_ASAP7_75t_L g1791 ( 
.A(n_1634),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1576),
.A2(n_576),
.B(n_575),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1535),
.A2(n_579),
.B(n_578),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1484),
.A2(n_771),
.B(n_770),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1595),
.B(n_583),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1593),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1546),
.A2(n_585),
.B(n_584),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1618),
.B(n_586),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1572),
.B(n_772),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1574),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1548),
.A2(n_589),
.B(n_588),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1551),
.A2(n_591),
.B(n_590),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1597),
.A2(n_775),
.B(n_779),
.C(n_773),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1559),
.A2(n_1486),
.B(n_1610),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1483),
.B(n_776),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1507),
.A2(n_593),
.B(n_592),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1581),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1487),
.B(n_780),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1608),
.B(n_782),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1579),
.A2(n_786),
.B1(n_787),
.B2(n_785),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1488),
.B(n_788),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1477),
.B(n_790),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1477),
.B(n_1505),
.Y(n_1813)
);

AO21x1_ASAP7_75t_L g1814 ( 
.A1(n_1615),
.A2(n_4),
.B(n_3),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1608),
.B(n_596),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1572),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1611),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1616),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1592),
.B(n_794),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1626),
.B(n_795),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1485),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1530),
.A2(n_599),
.B(n_598),
.Y(n_1822)
);

OAI21x1_ASAP7_75t_L g1823 ( 
.A1(n_1596),
.A2(n_604),
.B(n_603),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1647),
.A2(n_1539),
.B(n_1640),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1682),
.A2(n_1564),
.B(n_1636),
.C(n_1554),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1787),
.Y(n_1826)
);

OAI21xp33_ASAP7_75t_SL g1827 ( 
.A1(n_1674),
.A2(n_1517),
.B(n_1592),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1649),
.A2(n_1617),
.B(n_1607),
.Y(n_1828)
);

OR2x6_ASAP7_75t_SL g1829 ( 
.A(n_1735),
.B(n_797),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1745),
.B(n_1642),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1651),
.A2(n_1627),
.B(n_1623),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1817),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1701),
.B(n_1543),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1702),
.B(n_1642),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1728),
.B(n_1545),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1790),
.A2(n_1624),
.B1(n_1557),
.B2(n_1558),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1671),
.A2(n_1625),
.B1(n_1553),
.B2(n_1609),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_SL g1838 ( 
.A1(n_1736),
.A2(n_1568),
.B(n_1577),
.C(n_1544),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1679),
.A2(n_1782),
.B(n_1650),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1650),
.A2(n_1630),
.B(n_1629),
.Y(n_1840)
);

AO22x1_ASAP7_75t_L g1841 ( 
.A1(n_1741),
.A2(n_807),
.B1(n_809),
.B2(n_806),
.Y(n_1841)
);

A2O1A1Ixp33_ASAP7_75t_L g1842 ( 
.A1(n_1699),
.A2(n_1544),
.B(n_1526),
.C(n_1455),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1719),
.B(n_1448),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1688),
.B(n_1468),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1705),
.A2(n_1556),
.B(n_1555),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1655),
.B(n_1470),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1818),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1683),
.B(n_1479),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1663),
.A2(n_1635),
.B(n_1631),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1684),
.B(n_1481),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1648),
.A2(n_1462),
.B1(n_1515),
.B2(n_1499),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1677),
.Y(n_1852)
);

OAI21xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1663),
.A2(n_1813),
.B(n_1685),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1686),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1696),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1767),
.A2(n_1516),
.B1(n_1637),
.B2(n_1577),
.Y(n_1856)
);

O2A1O1Ixp33_ASAP7_75t_SL g1857 ( 
.A1(n_1720),
.A2(n_1582),
.B(n_1588),
.C(n_1587),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1645),
.B(n_810),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1737),
.A2(n_1575),
.B(n_1571),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1685),
.A2(n_1514),
.B(n_607),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1730),
.A2(n_1646),
.B(n_1657),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1693),
.A2(n_1514),
.B(n_608),
.Y(n_1862)
);

AND2x4_ASAP7_75t_SL g1863 ( 
.A(n_1654),
.B(n_1514),
.Y(n_1863)
);

OAI21xp33_ASAP7_75t_L g1864 ( 
.A1(n_1687),
.A2(n_816),
.B(n_811),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1695),
.B(n_819),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1690),
.B(n_1514),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1781),
.A2(n_823),
.B1(n_825),
.B2(n_822),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1766),
.A2(n_609),
.B(n_605),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1706),
.A2(n_829),
.B(n_827),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1680),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1704),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1656),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1726),
.B(n_830),
.Y(n_1873)
);

O2A1O1Ixp5_ASAP7_75t_L g1874 ( 
.A1(n_1754),
.A2(n_832),
.B(n_834),
.C(n_831),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1707),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1661),
.B(n_836),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1820),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1700),
.B(n_837),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1693),
.A2(n_616),
.B(n_615),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1673),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1780),
.A2(n_840),
.B1(n_843),
.B2(n_838),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1723),
.A2(n_846),
.B1(n_849),
.B2(n_844),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1658),
.B(n_1709),
.Y(n_1883)
);

AO21x1_ASAP7_75t_L g1884 ( 
.A1(n_1804),
.A2(n_2),
.B(n_4),
.Y(n_1884)
);

OA22x2_ASAP7_75t_L g1885 ( 
.A1(n_1789),
.A2(n_851),
.B1(n_858),
.B2(n_850),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1805),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1697),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1689),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1703),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1722),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1659),
.A2(n_611),
.B(n_610),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1755),
.B(n_10),
.Y(n_1892)
);

AO21x1_ASAP7_75t_L g1893 ( 
.A1(n_1643),
.A2(n_1664),
.B(n_1692),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1709),
.B(n_10),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1708),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1659),
.A2(n_614),
.B(n_11),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1738),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1717),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1652),
.A2(n_12),
.B(n_15),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1660),
.A2(n_15),
.B(n_16),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1653),
.B(n_16),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1669),
.A2(n_17),
.B(n_18),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1727),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1670),
.B(n_1785),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1715),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1788),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1808),
.B(n_19),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1739),
.Y(n_1908)
);

AOI33xp33_ASAP7_75t_L g1909 ( 
.A1(n_1665),
.A2(n_1747),
.A3(n_1711),
.B1(n_1772),
.B2(n_1810),
.B3(n_1752),
.Y(n_1909)
);

O2A1O1Ixp5_ASAP7_75t_L g1910 ( 
.A1(n_1758),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1701),
.B(n_22),
.Y(n_1911)
);

INVx3_ASAP7_75t_SL g1912 ( 
.A(n_1816),
.Y(n_1912)
);

AOI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1744),
.A2(n_23),
.B(n_24),
.Y(n_1913)
);

OAI22x1_ASAP7_75t_L g1914 ( 
.A1(n_1798),
.A2(n_555),
.B1(n_545),
.B2(n_27),
.Y(n_1914)
);

A2O1A1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1757),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1915)
);

O2A1O1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1763),
.A2(n_548),
.B(n_549),
.C(n_547),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1769),
.A2(n_25),
.B(n_26),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1759),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1770),
.A2(n_28),
.B(n_29),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1762),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1755),
.B(n_31),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1811),
.B(n_32),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1812),
.B(n_33),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1672),
.B(n_35),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1799),
.B(n_36),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1666),
.A2(n_37),
.B(n_38),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1644),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1799),
.B(n_39),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1666),
.A2(n_39),
.B(n_40),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1778),
.B(n_40),
.Y(n_1930)
);

AND2x6_ASAP7_75t_L g1931 ( 
.A(n_1771),
.B(n_41),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1675),
.A2(n_41),
.B(n_42),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1694),
.A2(n_42),
.B(n_43),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1815),
.B(n_44),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1760),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1740),
.B(n_45),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1794),
.B(n_45),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1676),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1787),
.B(n_46),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1757),
.B(n_47),
.C(n_48),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1794),
.B(n_47),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1742),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1802),
.B(n_49),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1779),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1714),
.A2(n_49),
.B(n_50),
.Y(n_1945)
);

NAND3xp33_ASAP7_75t_L g1946 ( 
.A(n_1678),
.B(n_50),
.C(n_51),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1821),
.B(n_51),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1667),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1714),
.A2(n_557),
.B(n_52),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1798),
.B(n_52),
.Y(n_1950)
);

INVx4_ASAP7_75t_L g1951 ( 
.A(n_1787),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1819),
.B(n_53),
.Y(n_1952)
);

O2A1O1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1803),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1953)
);

INVxp67_ASAP7_75t_SL g1954 ( 
.A(n_1765),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1776),
.B(n_55),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1784),
.Y(n_1956)
);

O2A1O1Ixp33_ASAP7_75t_L g1957 ( 
.A1(n_1681),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_R g1958 ( 
.A(n_1667),
.B(n_56),
.Y(n_1958)
);

NOR2xp67_ASAP7_75t_SL g1959 ( 
.A(n_1787),
.B(n_57),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1800),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1815),
.B(n_58),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1807),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1712),
.B(n_1743),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1775),
.B(n_1796),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1771),
.B(n_59),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1795),
.B(n_59),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1746),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1773),
.B(n_60),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1667),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1761),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1721),
.A2(n_61),
.B(n_62),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1792),
.A2(n_63),
.B(n_65),
.Y(n_1972)
);

OR2x6_ASAP7_75t_L g1973 ( 
.A(n_1793),
.B(n_65),
.Y(n_1973)
);

O2A1O1Ixp5_ASAP7_75t_L g1974 ( 
.A1(n_1814),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1809),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1806),
.A2(n_557),
.B(n_69),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1795),
.B(n_70),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1756),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1751),
.Y(n_1979)
);

OR2x6_ASAP7_75t_L g1980 ( 
.A(n_1797),
.B(n_72),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1718),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1774),
.B(n_74),
.Y(n_1982)
);

OR2x2_ASAP7_75t_SL g1983 ( 
.A(n_1753),
.B(n_75),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1753),
.Y(n_1984)
);

INVx4_ASAP7_75t_L g1985 ( 
.A(n_1753),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1768),
.B(n_76),
.Y(n_1986)
);

CKINVDCx16_ASAP7_75t_R g1987 ( 
.A(n_1786),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1732),
.A2(n_1698),
.B1(n_1791),
.B2(n_1662),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1822),
.A2(n_77),
.B(n_78),
.Y(n_1989)
);

OA22x2_ASAP7_75t_L g1990 ( 
.A1(n_1791),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_1990)
);

O2A1O1Ixp5_ASAP7_75t_SL g1991 ( 
.A1(n_1668),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1698),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1786),
.Y(n_1993)
);

OA22x2_ASAP7_75t_L g1994 ( 
.A1(n_1836),
.A2(n_1823),
.B1(n_1731),
.B2(n_1725),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_SL g1995 ( 
.A1(n_1825),
.A2(n_1801),
.B(n_1783),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1870),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1872),
.Y(n_1997)
);

NOR4xp25_ASAP7_75t_L g1998 ( 
.A(n_1940),
.B(n_1668),
.C(n_86),
.D(n_84),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_1866),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1987),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1967),
.B(n_1786),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1883),
.B(n_1710),
.Y(n_2002)
);

OAI21x1_ASAP7_75t_L g2003 ( 
.A1(n_1861),
.A2(n_1828),
.B(n_1831),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1978),
.B(n_1713),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1839),
.A2(n_1748),
.B(n_1691),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1835),
.B(n_1834),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_SL g2007 ( 
.A(n_1940),
.B(n_1777),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1833),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1830),
.B(n_1716),
.Y(n_2009)
);

BUFx3_ASAP7_75t_L g2010 ( 
.A(n_1979),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1934),
.B(n_1750),
.Y(n_2011)
);

AOI21xp33_ASAP7_75t_L g2012 ( 
.A1(n_1838),
.A2(n_1764),
.B(n_1734),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1905),
.Y(n_2013)
);

AO31x2_ASAP7_75t_L g2014 ( 
.A1(n_1893),
.A2(n_1884),
.A3(n_1840),
.B(n_1860),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1956),
.B(n_1701),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1836),
.A2(n_1724),
.B1(n_1749),
.B2(n_1729),
.Y(n_2016)
);

OAI21x1_ASAP7_75t_L g2017 ( 
.A1(n_1824),
.A2(n_1733),
.B(n_85),
.Y(n_2017)
);

OAI21x1_ASAP7_75t_L g2018 ( 
.A1(n_1868),
.A2(n_87),
.B(n_88),
.Y(n_2018)
);

NOR3xp33_ASAP7_75t_L g2019 ( 
.A(n_1909),
.B(n_87),
.C(n_88),
.Y(n_2019)
);

AOI211x1_ASAP7_75t_L g2020 ( 
.A1(n_1945),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_2020)
);

NOR2xp67_ASAP7_75t_L g2021 ( 
.A(n_1933),
.B(n_89),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_SL g2022 ( 
.A1(n_1915),
.A2(n_91),
.B(n_92),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_L g2023 ( 
.A1(n_1862),
.A2(n_92),
.B(n_93),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1961),
.B(n_93),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_1948),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1848),
.B(n_94),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_1938),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_2027)
);

BUFx10_ASAP7_75t_L g2028 ( 
.A(n_1905),
.Y(n_2028)
);

OAI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1891),
.A2(n_95),
.B(n_96),
.Y(n_2029)
);

OAI21x1_ASAP7_75t_L g2030 ( 
.A1(n_1849),
.A2(n_97),
.B(n_98),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1954),
.B(n_97),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1865),
.B(n_99),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1896),
.A2(n_100),
.B(n_101),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1879),
.A2(n_1913),
.B(n_1932),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1976),
.A2(n_100),
.B(n_101),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_SL g2036 ( 
.A1(n_1926),
.A2(n_102),
.B(n_103),
.Y(n_2036)
);

OAI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1917),
.A2(n_102),
.B(n_103),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1850),
.B(n_104),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1930),
.B(n_104),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1924),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_2040)
);

CKINVDCx11_ASAP7_75t_R g2041 ( 
.A(n_1829),
.Y(n_2041)
);

AO31x2_ASAP7_75t_L g2042 ( 
.A1(n_1929),
.A2(n_107),
.A3(n_105),
.B(n_106),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_1905),
.Y(n_2043)
);

A2O1A1Ixp33_ASAP7_75t_L g2044 ( 
.A1(n_1853),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_2044)
);

INVxp67_ASAP7_75t_L g2045 ( 
.A(n_1846),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1844),
.B(n_555),
.Y(n_2046)
);

AOI21x1_ASAP7_75t_L g2047 ( 
.A1(n_1949),
.A2(n_108),
.B(n_109),
.Y(n_2047)
);

OAI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1971),
.A2(n_1972),
.B(n_1827),
.Y(n_2048)
);

AOI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1937),
.A2(n_111),
.B(n_112),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1863),
.B(n_111),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1919),
.A2(n_112),
.B(n_113),
.Y(n_2051)
);

OAI21x1_ASAP7_75t_L g2052 ( 
.A1(n_1989),
.A2(n_113),
.B(n_114),
.Y(n_2052)
);

BUFx4f_ASAP7_75t_SL g2053 ( 
.A(n_1944),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1859),
.A2(n_114),
.B(n_115),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1941),
.B(n_115),
.Y(n_2055)
);

INVx4_ASAP7_75t_L g2056 ( 
.A(n_1826),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1936),
.B(n_554),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1963),
.B(n_1854),
.Y(n_2058)
);

OAI21x1_ASAP7_75t_L g2059 ( 
.A1(n_1902),
.A2(n_116),
.B(n_117),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1855),
.B(n_1871),
.Y(n_2060)
);

OAI21xp33_ASAP7_75t_L g2061 ( 
.A1(n_1982),
.A2(n_554),
.B(n_116),
.Y(n_2061)
);

AO21x1_ASAP7_75t_L g2062 ( 
.A1(n_1957),
.A2(n_1953),
.B(n_1916),
.Y(n_2062)
);

A2O1A1Ixp33_ASAP7_75t_L g2063 ( 
.A1(n_1874),
.A2(n_120),
.B(n_117),
.C(n_119),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1877),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_2064)
);

OR2x6_ASAP7_75t_L g2065 ( 
.A(n_1973),
.B(n_1980),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1857),
.A2(n_121),
.B(n_122),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1845),
.A2(n_123),
.B(n_124),
.Y(n_2067)
);

AO31x2_ASAP7_75t_L g2068 ( 
.A1(n_1988),
.A2(n_125),
.A3(n_123),
.B(n_124),
.Y(n_2068)
);

AO31x2_ASAP7_75t_L g2069 ( 
.A1(n_1837),
.A2(n_127),
.A3(n_125),
.B(n_126),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_1858),
.B(n_126),
.Y(n_2070)
);

OR2x6_ASAP7_75t_L g2071 ( 
.A(n_1973),
.B(n_127),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1875),
.B(n_553),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1895),
.B(n_553),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1898),
.B(n_128),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1903),
.B(n_128),
.Y(n_2075)
);

OAI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1946),
.A2(n_129),
.B(n_130),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1918),
.B(n_1935),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1880),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1852),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1912),
.Y(n_2080)
);

OAI21x1_ASAP7_75t_L g2081 ( 
.A1(n_1991),
.A2(n_129),
.B(n_130),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1904),
.B(n_131),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1927),
.B(n_132),
.Y(n_2083)
);

O2A1O1Ixp33_ASAP7_75t_SL g2084 ( 
.A1(n_1925),
.A2(n_137),
.B(n_133),
.C(n_136),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_1851),
.A2(n_136),
.B(n_137),
.Y(n_2085)
);

OAI21x1_ASAP7_75t_L g2086 ( 
.A1(n_1887),
.A2(n_138),
.B(n_139),
.Y(n_2086)
);

AND3x1_ASAP7_75t_L g2087 ( 
.A(n_1886),
.B(n_140),
.C(n_141),
.Y(n_2087)
);

OAI21x1_ASAP7_75t_L g2088 ( 
.A1(n_1889),
.A2(n_140),
.B(n_141),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1907),
.B(n_1922),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1890),
.A2(n_142),
.B(n_143),
.Y(n_2090)
);

A2O1A1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1946),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1892),
.B(n_144),
.Y(n_2092)
);

OAI21x1_ASAP7_75t_L g2093 ( 
.A1(n_1897),
.A2(n_145),
.B(n_146),
.Y(n_2093)
);

AOI21x1_ASAP7_75t_L g2094 ( 
.A1(n_1959),
.A2(n_145),
.B(n_147),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_1958),
.Y(n_2095)
);

OAI21x1_ASAP7_75t_SL g2096 ( 
.A1(n_1899),
.A2(n_147),
.B(n_148),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1921),
.B(n_148),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_1908),
.A2(n_149),
.B(n_150),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1942),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_L g2100 ( 
.A1(n_1964),
.A2(n_150),
.B(n_151),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1993),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1910),
.A2(n_152),
.B(n_153),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1974),
.A2(n_152),
.B(n_153),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1960),
.B(n_154),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1842),
.A2(n_155),
.B(n_156),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_1900),
.A2(n_1856),
.B(n_1847),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1985),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1962),
.B(n_552),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_1832),
.A2(n_155),
.B(n_156),
.Y(n_2109)
);

NAND2x1p5_ASAP7_75t_L g2110 ( 
.A(n_1826),
.B(n_157),
.Y(n_2110)
);

INVx2_ASAP7_75t_SL g2111 ( 
.A(n_1985),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2048),
.A2(n_1980),
.B(n_1973),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2087),
.A2(n_1983),
.B1(n_1886),
.B2(n_1975),
.Y(n_2113)
);

INVx1_ASAP7_75t_SL g2114 ( 
.A(n_1996),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1999),
.B(n_1969),
.Y(n_2115)
);

INVx3_ASAP7_75t_SL g2116 ( 
.A(n_2095),
.Y(n_2116)
);

INVx1_ASAP7_75t_SL g2117 ( 
.A(n_1996),
.Y(n_2117)
);

HB1xp67_ASAP7_75t_L g2118 ( 
.A(n_1999),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2025),
.B(n_2000),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1997),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2106),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_2013),
.Y(n_2122)
);

AOI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_2019),
.A2(n_2070),
.B1(n_2061),
.B2(n_2087),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_2078),
.Y(n_2124)
);

AOI21xp33_ASAP7_75t_L g2125 ( 
.A1(n_2033),
.A2(n_1986),
.B(n_1952),
.Y(n_2125)
);

O2A1O1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_2033),
.A2(n_1928),
.B(n_1977),
.C(n_1966),
.Y(n_2126)
);

AOI221x1_ASAP7_75t_L g2127 ( 
.A1(n_2061),
.A2(n_2036),
.B1(n_2022),
.B2(n_2076),
.C(n_2067),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2099),
.B(n_1947),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2001),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_2053),
.Y(n_2130)
);

AOI221xp5_ASAP7_75t_L g2131 ( 
.A1(n_1998),
.A2(n_1906),
.B1(n_1920),
.B2(n_1888),
.C(n_1970),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_2028),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2065),
.Y(n_2133)
);

BUFx2_ASAP7_75t_L g2134 ( 
.A(n_2008),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2043),
.B(n_1969),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_2065),
.B(n_1911),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_2065),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2060),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_2008),
.B(n_1911),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2024),
.B(n_1984),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_2013),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2077),
.Y(n_2142)
);

CKINVDCx6p67_ASAP7_75t_R g2143 ( 
.A(n_2010),
.Y(n_2143)
);

BUFx10_ASAP7_75t_L g2144 ( 
.A(n_2079),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2031),
.B(n_1923),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2040),
.A2(n_1990),
.B1(n_1981),
.B2(n_1968),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2058),
.Y(n_2147)
);

AND2x2_ASAP7_75t_SL g2148 ( 
.A(n_1998),
.B(n_1951),
.Y(n_2148)
);

A2O1A1Ixp33_ASAP7_75t_L g2149 ( 
.A1(n_2076),
.A2(n_1869),
.B(n_1864),
.C(n_1965),
.Y(n_2149)
);

AOI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_2003),
.A2(n_1980),
.B(n_1943),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2069),
.Y(n_2151)
);

AO32x1_ASAP7_75t_L g2152 ( 
.A1(n_2027),
.A2(n_1992),
.A3(n_1867),
.B1(n_1873),
.B2(n_1841),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2069),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2006),
.B(n_1876),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2015),
.B(n_1833),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_2013),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2069),
.B(n_1894),
.Y(n_2157)
);

INVx5_ASAP7_75t_L g2158 ( 
.A(n_2071),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_2079),
.Y(n_2159)
);

CKINVDCx6p67_ASAP7_75t_R g2160 ( 
.A(n_2080),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2071),
.B(n_1943),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2092),
.B(n_1914),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2071),
.B(n_1943),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2002),
.Y(n_2164)
);

BUFx10_ASAP7_75t_L g2165 ( 
.A(n_2079),
.Y(n_2165)
);

INVxp67_ASAP7_75t_SL g2166 ( 
.A(n_2004),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2068),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2009),
.B(n_1955),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2097),
.B(n_1885),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_SL g2170 ( 
.A1(n_2105),
.A2(n_1931),
.B1(n_1939),
.B2(n_1878),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2089),
.B(n_1864),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2014),
.B(n_1931),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2014),
.B(n_1931),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_2107),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2068),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2014),
.B(n_2048),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_2111),
.B(n_1931),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2045),
.B(n_2032),
.Y(n_2178)
);

OAI21x1_ASAP7_75t_SL g2179 ( 
.A1(n_2105),
.A2(n_1843),
.B(n_1882),
.Y(n_2179)
);

BUFx3_ASAP7_75t_L g2180 ( 
.A(n_2028),
.Y(n_2180)
);

INVx5_ASAP7_75t_L g2181 ( 
.A(n_2056),
.Y(n_2181)
);

INVx2_ASAP7_75t_SL g2182 ( 
.A(n_2107),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_2107),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2056),
.B(n_1901),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2068),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2049),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_2082),
.B(n_2083),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2101),
.Y(n_2188)
);

AOI22xp33_ASAP7_75t_L g2189 ( 
.A1(n_2170),
.A2(n_2062),
.B1(n_2040),
.B2(n_2007),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2123),
.A2(n_2007),
.B1(n_2091),
.B2(n_2044),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2166),
.B(n_2042),
.Y(n_2191)
);

OAI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_2127),
.A2(n_2055),
.B1(n_2066),
.B2(n_2021),
.Y(n_2192)
);

BUFx3_ASAP7_75t_L g2193 ( 
.A(n_2130),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2124),
.Y(n_2194)
);

INVx4_ASAP7_75t_L g2195 ( 
.A(n_2183),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_2113),
.A2(n_2096),
.B1(n_2011),
.B2(n_2021),
.Y(n_2196)
);

BUFx4f_ASAP7_75t_L g2197 ( 
.A(n_2160),
.Y(n_2197)
);

AOI22xp33_ASAP7_75t_L g2198 ( 
.A1(n_2113),
.A2(n_2131),
.B1(n_2125),
.B2(n_2146),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2120),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_2183),
.Y(n_2200)
);

BUFx10_ASAP7_75t_L g2201 ( 
.A(n_2183),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_SL g2202 ( 
.A1(n_2112),
.A2(n_2063),
.B(n_2110),
.Y(n_2202)
);

CKINVDCx11_ASAP7_75t_R g2203 ( 
.A(n_2116),
.Y(n_2203)
);

INVx2_ASAP7_75t_SL g2204 ( 
.A(n_2144),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_2159),
.Y(n_2205)
);

AOI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_2150),
.A2(n_1995),
.B(n_2005),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_SL g2207 ( 
.A1(n_2146),
.A2(n_2029),
.B1(n_2023),
.B2(n_2054),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2118),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_2159),
.Y(n_2209)
);

AOI22xp33_ASAP7_75t_L g2210 ( 
.A1(n_2131),
.A2(n_1869),
.B1(n_2041),
.B2(n_1994),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2133),
.Y(n_2211)
);

CKINVDCx6p67_ASAP7_75t_R g2212 ( 
.A(n_2143),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_2159),
.Y(n_2213)
);

INVx6_ASAP7_75t_L g2214 ( 
.A(n_2144),
.Y(n_2214)
);

CKINVDCx11_ASAP7_75t_R g2215 ( 
.A(n_2165),
.Y(n_2215)
);

INVx6_ASAP7_75t_L g2216 ( 
.A(n_2165),
.Y(n_2216)
);

HB1xp67_ASAP7_75t_L g2217 ( 
.A(n_2164),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2164),
.B(n_2147),
.Y(n_2218)
);

AOI22xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2158),
.A2(n_2030),
.B1(n_2064),
.B2(n_2085),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2114),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_SL g2221 ( 
.A1(n_2158),
.A2(n_2052),
.B1(n_2035),
.B2(n_2051),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2137),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_2186),
.Y(n_2223)
);

BUFx4_ASAP7_75t_SL g2224 ( 
.A(n_2180),
.Y(n_2224)
);

BUFx12f_ASAP7_75t_L g2225 ( 
.A(n_2132),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2114),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_2119),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_2122),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_2134),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2151),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2153),
.Y(n_2231)
);

INVx4_ASAP7_75t_L g2232 ( 
.A(n_2181),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2149),
.A2(n_2020),
.B1(n_2057),
.B2(n_2047),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_2115),
.Y(n_2234)
);

CKINVDCx6p67_ASAP7_75t_R g2235 ( 
.A(n_2156),
.Y(n_2235)
);

INVx6_ASAP7_75t_L g2236 ( 
.A(n_2122),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2167),
.Y(n_2237)
);

INVx6_ASAP7_75t_L g2238 ( 
.A(n_2122),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2175),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_SL g2240 ( 
.A1(n_2233),
.A2(n_2163),
.B(n_2161),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2217),
.B(n_2117),
.Y(n_2241)
);

AND2x4_ASAP7_75t_L g2242 ( 
.A(n_2211),
.B(n_2117),
.Y(n_2242)
);

BUFx2_ASAP7_75t_SL g2243 ( 
.A(n_2193),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2230),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2222),
.B(n_2223),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2198),
.A2(n_2158),
.B1(n_2020),
.B2(n_2161),
.Y(n_2246)
);

NAND2xp33_ASAP7_75t_SL g2247 ( 
.A(n_2189),
.B(n_2163),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2218),
.B(n_2129),
.Y(n_2248)
);

A2O1A1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2202),
.A2(n_2126),
.B(n_2125),
.C(n_2187),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2218),
.B(n_2129),
.Y(n_2250)
);

O2A1O1Ixp5_ASAP7_75t_L g2251 ( 
.A1(n_2233),
.A2(n_2176),
.B(n_2157),
.C(n_2150),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_SL g2252 ( 
.A1(n_2192),
.A2(n_2173),
.B(n_2172),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_2194),
.Y(n_2253)
);

OAI22xp5_ASAP7_75t_L g2254 ( 
.A1(n_2190),
.A2(n_2158),
.B1(n_2148),
.B2(n_2136),
.Y(n_2254)
);

INVx2_ASAP7_75t_SL g2255 ( 
.A(n_2229),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2220),
.B(n_2157),
.Y(n_2256)
);

O2A1O1Ixp33_ASAP7_75t_L g2257 ( 
.A1(n_2202),
.A2(n_2171),
.B(n_2084),
.C(n_2176),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2234),
.B(n_2185),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2226),
.B(n_2128),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_SL g2260 ( 
.A1(n_2190),
.A2(n_2206),
.B(n_2173),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2208),
.B(n_2172),
.Y(n_2261)
);

OAI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_2210),
.A2(n_2196),
.B1(n_2207),
.B2(n_2219),
.Y(n_2262)
);

O2A1O1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_2206),
.A2(n_2171),
.B(n_2179),
.C(n_2154),
.Y(n_2263)
);

INVx3_ASAP7_75t_SL g2264 ( 
.A(n_2212),
.Y(n_2264)
);

OA21x2_ASAP7_75t_L g2265 ( 
.A1(n_2191),
.A2(n_2121),
.B(n_2034),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2227),
.B(n_2178),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2244),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2253),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_R g2269 ( 
.A(n_2242),
.B(n_2169),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2245),
.Y(n_2270)
);

OAI21xp33_ASAP7_75t_L g2271 ( 
.A1(n_2262),
.A2(n_2207),
.B(n_2191),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2243),
.Y(n_2272)
);

OR2x6_ASAP7_75t_L g2273 ( 
.A(n_2260),
.B(n_2232),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_2241),
.B(n_2223),
.Y(n_2274)
);

OR2x2_ASAP7_75t_SL g2275 ( 
.A(n_2261),
.B(n_2214),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2245),
.Y(n_2276)
);

NAND2xp33_ASAP7_75t_R g2277 ( 
.A(n_2265),
.B(n_2154),
.Y(n_2277)
);

AO21x2_ASAP7_75t_L g2278 ( 
.A1(n_2271),
.A2(n_2252),
.B(n_2240),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2267),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2268),
.B(n_2245),
.Y(n_2280)
);

AOI21x1_ASAP7_75t_L g2281 ( 
.A1(n_2273),
.A2(n_2254),
.B(n_2256),
.Y(n_2281)
);

AOI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_2270),
.A2(n_2249),
.B1(n_2251),
.B2(n_2263),
.C(n_2247),
.Y(n_2282)
);

OA21x2_ASAP7_75t_L g2283 ( 
.A1(n_2276),
.A2(n_2249),
.B(n_2237),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2274),
.Y(n_2284)
);

AO21x2_ASAP7_75t_L g2285 ( 
.A1(n_2277),
.A2(n_2246),
.B(n_2239),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2273),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2278),
.B(n_2273),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2282),
.B(n_2242),
.Y(n_2288)
);

OR2x2_ASAP7_75t_L g2289 ( 
.A(n_2284),
.B(n_2275),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2279),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2283),
.Y(n_2291)
);

NAND2x1p5_ASAP7_75t_SL g2292 ( 
.A(n_2286),
.B(n_2204),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2279),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2278),
.B(n_2286),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2284),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2280),
.B(n_2242),
.Y(n_2296)
);

OAI221xp5_ASAP7_75t_L g2297 ( 
.A1(n_2288),
.A2(n_2247),
.B1(n_2286),
.B2(n_2281),
.C(n_2277),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2291),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2287),
.A2(n_2278),
.B1(n_2285),
.B2(n_2289),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2291),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2290),
.Y(n_2301)
);

BUFx3_ASAP7_75t_L g2302 ( 
.A(n_2294),
.Y(n_2302)
);

AOI31xp33_ASAP7_75t_L g2303 ( 
.A1(n_2287),
.A2(n_2272),
.A3(n_2269),
.B(n_2278),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2294),
.B(n_2283),
.Y(n_2304)
);

AOI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2295),
.A2(n_2285),
.B1(n_2283),
.B2(n_2219),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2293),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_2296),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_2292),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2298),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2308),
.B(n_2283),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2306),
.B(n_2292),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2302),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2302),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2300),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2307),
.B(n_2264),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_2302),
.B(n_2280),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2300),
.B(n_2281),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2312),
.B(n_2301),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2315),
.B(n_2311),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2309),
.B(n_2301),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2314),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2319),
.B(n_2312),
.Y(n_2322)
);

AOI22xp5_ASAP7_75t_L g2323 ( 
.A1(n_2318),
.A2(n_2297),
.B1(n_2285),
.B2(n_2305),
.Y(n_2323)
);

OR2x6_ASAP7_75t_L g2324 ( 
.A(n_2320),
.B(n_2313),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2318),
.B(n_2313),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2322),
.B(n_2310),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2324),
.Y(n_2327)
);

NOR2x1p5_ASAP7_75t_SL g2328 ( 
.A(n_2324),
.B(n_2300),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2325),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2323),
.B(n_2321),
.Y(n_2330)
);

INVxp67_ASAP7_75t_L g2331 ( 
.A(n_2325),
.Y(n_2331)
);

INVx5_ASAP7_75t_L g2332 ( 
.A(n_2326),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2329),
.Y(n_2333)
);

AND3x1_ASAP7_75t_L g2334 ( 
.A(n_2327),
.B(n_2320),
.C(n_2310),
.Y(n_2334)
);

AND2x4_ASAP7_75t_L g2335 ( 
.A(n_2331),
.B(n_2316),
.Y(n_2335)
);

AOI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2330),
.A2(n_2299),
.B1(n_2305),
.B2(n_2285),
.Y(n_2336)
);

INVxp67_ASAP7_75t_SL g2337 ( 
.A(n_2330),
.Y(n_2337)
);

OAI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2328),
.A2(n_2303),
.B1(n_2317),
.B2(n_2264),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2328),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2328),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2328),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2339),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2338),
.A2(n_2317),
.B(n_2304),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2340),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2341),
.Y(n_2345)
);

INVxp67_ASAP7_75t_L g2346 ( 
.A(n_2334),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_2332),
.B(n_2304),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2333),
.Y(n_2348)
);

AOI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_2337),
.A2(n_2257),
.B1(n_1881),
.B2(n_2039),
.C(n_2197),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2332),
.B(n_2203),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2335),
.B(n_2255),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2336),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2332),
.Y(n_2353)
);

OAI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2336),
.A2(n_2197),
.B1(n_1950),
.B2(n_2216),
.C(n_2214),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2347),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2353),
.Y(n_2356)
);

AOI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2350),
.A2(n_2225),
.B1(n_2215),
.B2(n_2216),
.Y(n_2357)
);

O2A1O1Ixp33_ASAP7_75t_SL g2358 ( 
.A1(n_2346),
.A2(n_2224),
.B(n_2046),
.C(n_2026),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2351),
.A2(n_2255),
.B1(n_2235),
.B2(n_2250),
.Y(n_2359)
);

A2O1A1Ixp33_ASAP7_75t_L g2360 ( 
.A1(n_2343),
.A2(n_2145),
.B(n_2100),
.C(n_2162),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2348),
.B(n_2266),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2348),
.B(n_2140),
.Y(n_2362)
);

O2A1O1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2352),
.A2(n_2342),
.B(n_2345),
.C(n_2344),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2354),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_SL g2365 ( 
.A(n_2349),
.B(n_1939),
.C(n_2038),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2347),
.B(n_2248),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2347),
.B(n_2258),
.Y(n_2367)
);

OAI322xp33_ASAP7_75t_L g2368 ( 
.A1(n_2346),
.A2(n_2075),
.A3(n_2073),
.B1(n_2104),
.B2(n_2108),
.C1(n_2074),
.C2(n_2072),
.Y(n_2368)
);

AOI221x1_ASAP7_75t_L g2369 ( 
.A1(n_2342),
.A2(n_2184),
.B1(n_159),
.B2(n_157),
.C(n_158),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2355),
.B(n_2265),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2361),
.B(n_2258),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2362),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2356),
.B(n_2265),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2357),
.B(n_2259),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2367),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2364),
.B(n_2195),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2369),
.B(n_2184),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2366),
.B(n_158),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2359),
.Y(n_2379)
);

OAI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2363),
.A2(n_2238),
.B1(n_2236),
.B2(n_2195),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2358),
.Y(n_2381)
);

NAND2xp33_ASAP7_75t_L g2382 ( 
.A(n_2360),
.B(n_2141),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2365),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2377),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2376),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2371),
.B(n_2368),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2381),
.B(n_2136),
.Y(n_2387)
);

OAI21xp33_ASAP7_75t_L g2388 ( 
.A1(n_2379),
.A2(n_2050),
.B(n_2182),
.Y(n_2388)
);

OAI21xp33_ASAP7_75t_L g2389 ( 
.A1(n_2374),
.A2(n_2050),
.B(n_2168),
.Y(n_2389)
);

NOR3xp33_ASAP7_75t_L g2390 ( 
.A(n_2375),
.B(n_2094),
.C(n_2168),
.Y(n_2390)
);

O2A1O1Ixp33_ASAP7_75t_SL g2391 ( 
.A1(n_2380),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2378),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2372),
.Y(n_2393)
);

AOI211xp5_ASAP7_75t_SL g2394 ( 
.A1(n_2383),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2380),
.B(n_162),
.Y(n_2395)
);

INVx1_ASAP7_75t_SL g2396 ( 
.A(n_2373),
.Y(n_2396)
);

AND3x1_ASAP7_75t_L g2397 ( 
.A(n_2370),
.B(n_163),
.C(n_164),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2382),
.A2(n_2152),
.B(n_2037),
.Y(n_2398)
);

AOI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2376),
.A2(n_2236),
.B1(n_2238),
.B2(n_2200),
.Y(n_2399)
);

NAND4xp25_ASAP7_75t_SL g2400 ( 
.A(n_2377),
.B(n_2221),
.C(n_2135),
.D(n_2188),
.Y(n_2400)
);

NAND4xp25_ASAP7_75t_L g2401 ( 
.A(n_2376),
.B(n_2232),
.C(n_2174),
.D(n_2177),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_2377),
.B(n_163),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2377),
.B(n_2141),
.Y(n_2403)
);

BUFx2_ASAP7_75t_L g2404 ( 
.A(n_2377),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2377),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2387),
.A2(n_2200),
.B1(n_2209),
.B2(n_2205),
.Y(n_2406)
);

AOI211x1_ASAP7_75t_L g2407 ( 
.A1(n_2403),
.A2(n_2231),
.B(n_167),
.C(n_165),
.Y(n_2407)
);

OAI21xp33_ASAP7_75t_L g2408 ( 
.A1(n_2388),
.A2(n_2200),
.B(n_2205),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2391),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2394),
.B(n_165),
.Y(n_2410)
);

OAI211xp5_ASAP7_75t_L g2411 ( 
.A1(n_2402),
.A2(n_169),
.B(n_166),
.C(n_168),
.Y(n_2411)
);

NOR2x1_ASAP7_75t_L g2412 ( 
.A(n_2404),
.B(n_166),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2395),
.B(n_168),
.Y(n_2413)
);

NOR2x1_ASAP7_75t_L g2414 ( 
.A(n_2384),
.B(n_2405),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2385),
.B(n_169),
.Y(n_2415)
);

AOI22xp33_ASAP7_75t_L g2416 ( 
.A1(n_2400),
.A2(n_2141),
.B1(n_2209),
.B2(n_2205),
.Y(n_2416)
);

AOI211xp5_ASAP7_75t_L g2417 ( 
.A1(n_2393),
.A2(n_173),
.B(n_170),
.C(n_171),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_SL g2418 ( 
.A(n_2396),
.B(n_170),
.C(n_171),
.Y(n_2418)
);

AOI21xp33_ASAP7_75t_SL g2419 ( 
.A1(n_2386),
.A2(n_173),
.B(n_174),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2397),
.Y(n_2420)
);

OAI21xp33_ASAP7_75t_SL g2421 ( 
.A1(n_2401),
.A2(n_2088),
.B(n_2086),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2392),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2389),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2399),
.B(n_174),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2390),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_2398),
.Y(n_2426)
);

AOI211xp5_ASAP7_75t_L g2427 ( 
.A1(n_2391),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_2427)
);

OAI321xp33_ASAP7_75t_L g2428 ( 
.A1(n_2384),
.A2(n_2213),
.A3(n_2209),
.B1(n_2228),
.B2(n_178),
.C(n_180),
.Y(n_2428)
);

NOR2xp67_ASAP7_75t_L g2429 ( 
.A(n_2384),
.B(n_176),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_L g2430 ( 
.A(n_2384),
.B(n_2093),
.C(n_2090),
.Y(n_2430)
);

OAI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2399),
.A2(n_2181),
.B1(n_2213),
.B2(n_2228),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2394),
.B(n_177),
.Y(n_2432)
);

NAND4xp25_ASAP7_75t_L g2433 ( 
.A(n_2386),
.B(n_180),
.C(n_178),
.D(n_179),
.Y(n_2433)
);

OAI21xp33_ASAP7_75t_L g2434 ( 
.A1(n_2387),
.A2(n_2213),
.B(n_2228),
.Y(n_2434)
);

AOI221x1_ASAP7_75t_L g2435 ( 
.A1(n_2402),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_2435)
);

NOR2x1_ASAP7_75t_L g2436 ( 
.A(n_2404),
.B(n_182),
.Y(n_2436)
);

NAND3xp33_ASAP7_75t_SL g2437 ( 
.A(n_2394),
.B(n_183),
.C(n_184),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2404),
.Y(n_2438)
);

AOI211x1_ASAP7_75t_L g2439 ( 
.A1(n_2403),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2394),
.B(n_185),
.Y(n_2440)
);

AOI21xp5_ASAP7_75t_L g2441 ( 
.A1(n_2391),
.A2(n_2152),
.B(n_2098),
.Y(n_2441)
);

O2A1O1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_2391),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2429),
.B(n_2409),
.Y(n_2443)
);

OAI211xp5_ASAP7_75t_L g2444 ( 
.A1(n_2419),
.A2(n_2427),
.B(n_2433),
.C(n_2442),
.Y(n_2444)
);

OAI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2414),
.A2(n_2109),
.B(n_2059),
.Y(n_2445)
);

NOR3xp33_ASAP7_75t_L g2446 ( 
.A(n_2422),
.B(n_188),
.C(n_190),
.Y(n_2446)
);

NAND4xp75_ASAP7_75t_L g2447 ( 
.A(n_2412),
.B(n_192),
.C(n_190),
.D(n_191),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2437),
.B(n_191),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_SL g2449 ( 
.A(n_2420),
.B(n_2181),
.Y(n_2449)
);

AOI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2438),
.A2(n_2177),
.B1(n_2201),
.B2(n_2155),
.Y(n_2450)
);

NAND4xp25_ASAP7_75t_L g2451 ( 
.A(n_2439),
.B(n_195),
.C(n_192),
.D(n_194),
.Y(n_2451)
);

NAND4xp25_ASAP7_75t_L g2452 ( 
.A(n_2407),
.B(n_197),
.C(n_194),
.D(n_195),
.Y(n_2452)
);

NAND3xp33_ASAP7_75t_L g2453 ( 
.A(n_2436),
.B(n_2435),
.C(n_2432),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2416),
.A2(n_2181),
.B1(n_2221),
.B2(n_2155),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2410),
.B(n_2201),
.Y(n_2455)
);

NAND3xp33_ASAP7_75t_L g2456 ( 
.A(n_2440),
.B(n_197),
.C(n_198),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2418),
.B(n_2415),
.Y(n_2457)
);

OAI211xp5_ASAP7_75t_L g2458 ( 
.A1(n_2411),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_2458)
);

AOI221xp5_ASAP7_75t_L g2459 ( 
.A1(n_2428),
.A2(n_202),
.B1(n_199),
.B2(n_201),
.C(n_203),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_L g2460 ( 
.A(n_2417),
.B(n_201),
.C(n_202),
.Y(n_2460)
);

NOR4xp25_ASAP7_75t_L g2461 ( 
.A(n_2426),
.B(n_205),
.C(n_203),
.D(n_204),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2413),
.Y(n_2462)
);

OAI221xp5_ASAP7_75t_L g2463 ( 
.A1(n_2434),
.A2(n_2408),
.B1(n_2424),
.B2(n_2423),
.C(n_2425),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2406),
.Y(n_2464)
);

NOR2x1_ASAP7_75t_L g2465 ( 
.A(n_2431),
.B(n_206),
.Y(n_2465)
);

NAND3xp33_ASAP7_75t_SL g2466 ( 
.A(n_2441),
.B(n_206),
.C(n_207),
.Y(n_2466)
);

OAI211xp5_ASAP7_75t_L g2467 ( 
.A1(n_2421),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2430),
.B(n_208),
.Y(n_2468)
);

OR3x1_ASAP7_75t_L g2469 ( 
.A(n_2428),
.B(n_209),
.C(n_210),
.Y(n_2469)
);

AND4x1_ASAP7_75t_L g2470 ( 
.A(n_2414),
.B(n_213),
.C(n_211),
.D(n_212),
.Y(n_2470)
);

NAND4xp25_ASAP7_75t_SL g2471 ( 
.A(n_2427),
.B(n_213),
.C(n_211),
.D(n_212),
.Y(n_2471)
);

NAND3xp33_ASAP7_75t_SL g2472 ( 
.A(n_2427),
.B(n_214),
.C(n_216),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_L g2473 ( 
.A(n_2427),
.B(n_216),
.C(n_217),
.Y(n_2473)
);

NAND3xp33_ASAP7_75t_L g2474 ( 
.A(n_2427),
.B(n_218),
.C(n_219),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_2433),
.B(n_218),
.C(n_219),
.Y(n_2475)
);

OAI211xp5_ASAP7_75t_L g2476 ( 
.A1(n_2419),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_2476)
);

NAND3xp33_ASAP7_75t_L g2477 ( 
.A(n_2427),
.B(n_221),
.C(n_222),
.Y(n_2477)
);

OAI21xp33_ASAP7_75t_L g2478 ( 
.A1(n_2434),
.A2(n_2115),
.B(n_2012),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2410),
.Y(n_2479)
);

OAI221xp5_ASAP7_75t_L g2480 ( 
.A1(n_2433),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.C(n_226),
.Y(n_2480)
);

NOR3x1_ASAP7_75t_L g2481 ( 
.A(n_2480),
.B(n_2453),
.C(n_2473),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2470),
.Y(n_2482)
);

NAND4xp25_ASAP7_75t_L g2483 ( 
.A(n_2459),
.B(n_226),
.C(n_223),
.D(n_224),
.Y(n_2483)
);

NOR2xp67_ASAP7_75t_L g2484 ( 
.A(n_2451),
.B(n_2452),
.Y(n_2484)
);

NOR3xp33_ASAP7_75t_L g2485 ( 
.A(n_2463),
.B(n_227),
.C(n_228),
.Y(n_2485)
);

NOR2xp67_ASAP7_75t_L g2486 ( 
.A(n_2471),
.B(n_227),
.Y(n_2486)
);

OAI211xp5_ASAP7_75t_SL g2487 ( 
.A1(n_2443),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2461),
.B(n_230),
.Y(n_2488)
);

NOR3xp33_ASAP7_75t_L g2489 ( 
.A(n_2456),
.B(n_231),
.C(n_232),
.Y(n_2489)
);

NAND4xp25_ASAP7_75t_L g2490 ( 
.A(n_2475),
.B(n_233),
.C(n_231),
.D(n_232),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2447),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2446),
.B(n_233),
.Y(n_2492)
);

NOR3xp33_ASAP7_75t_SL g2493 ( 
.A(n_2472),
.B(n_234),
.C(n_235),
.Y(n_2493)
);

NOR3xp33_ASAP7_75t_L g2494 ( 
.A(n_2448),
.B(n_234),
.C(n_236),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_SL g2495 ( 
.A(n_2474),
.B(n_237),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2455),
.B(n_237),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2469),
.Y(n_2497)
);

AOI211xp5_ASAP7_75t_L g2498 ( 
.A1(n_2458),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2498)
);

AOI211xp5_ASAP7_75t_L g2499 ( 
.A1(n_2476),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_2444),
.B(n_241),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2449),
.B(n_242),
.Y(n_2501)
);

OAI221xp5_ASAP7_75t_SL g2502 ( 
.A1(n_2467),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_2502)
);

NOR2x1_ASAP7_75t_L g2503 ( 
.A(n_2457),
.B(n_243),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2479),
.B(n_245),
.Y(n_2504)
);

NOR3xp33_ASAP7_75t_L g2505 ( 
.A(n_2464),
.B(n_247),
.C(n_248),
.Y(n_2505)
);

AOI221xp5_ASAP7_75t_L g2506 ( 
.A1(n_2466),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.C(n_250),
.Y(n_2506)
);

OAI322xp33_ASAP7_75t_L g2507 ( 
.A1(n_2468),
.A2(n_2462),
.A3(n_2477),
.B1(n_2460),
.B2(n_2454),
.C1(n_2465),
.C2(n_2450),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2478),
.B(n_249),
.Y(n_2508)
);

NAND4xp25_ASAP7_75t_L g2509 ( 
.A(n_2445),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2509)
);

OAI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2443),
.A2(n_2102),
.B(n_2103),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2470),
.Y(n_2511)
);

NOR3x1_ASAP7_75t_L g2512 ( 
.A(n_2480),
.B(n_253),
.C(n_254),
.Y(n_2512)
);

OAI321xp33_ASAP7_75t_L g2513 ( 
.A1(n_2463),
.A2(n_256),
.A3(n_259),
.B1(n_254),
.B2(n_255),
.C(n_257),
.Y(n_2513)
);

AND4x1_ASAP7_75t_L g2514 ( 
.A(n_2453),
.B(n_259),
.C(n_255),
.D(n_257),
.Y(n_2514)
);

OAI22xp33_ASAP7_75t_L g2515 ( 
.A1(n_2449),
.A2(n_2199),
.B1(n_2138),
.B2(n_2016),
.Y(n_2515)
);

NAND3xp33_ASAP7_75t_SL g2516 ( 
.A(n_2461),
.B(n_260),
.C(n_261),
.Y(n_2516)
);

AOI221xp5_ASAP7_75t_L g2517 ( 
.A1(n_2461),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2470),
.Y(n_2518)
);

NOR2x1_ASAP7_75t_L g2519 ( 
.A(n_2447),
.B(n_262),
.Y(n_2519)
);

OAI211xp5_ASAP7_75t_L g2520 ( 
.A1(n_2459),
.A2(n_266),
.B(n_263),
.C(n_265),
.Y(n_2520)
);

NAND4xp25_ASAP7_75t_L g2521 ( 
.A(n_2459),
.B(n_268),
.C(n_266),
.D(n_267),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_2443),
.A2(n_2152),
.B(n_268),
.Y(n_2522)
);

AOI221x1_ASAP7_75t_L g2523 ( 
.A1(n_2443),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_272),
.Y(n_2523)
);

AOI221xp5_ASAP7_75t_L g2524 ( 
.A1(n_2461),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.C(n_273),
.Y(n_2524)
);

NAND3xp33_ASAP7_75t_L g2525 ( 
.A(n_2470),
.B(n_273),
.C(n_274),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2470),
.B(n_275),
.Y(n_2526)
);

NAND4xp25_ASAP7_75t_L g2527 ( 
.A(n_2459),
.B(n_277),
.C(n_275),
.D(n_276),
.Y(n_2527)
);

NAND3x1_ASAP7_75t_L g2528 ( 
.A(n_2470),
.B(n_276),
.C(n_277),
.Y(n_2528)
);

OAI211xp5_ASAP7_75t_L g2529 ( 
.A1(n_2459),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2529)
);

O2A1O1Ixp33_ASAP7_75t_L g2530 ( 
.A1(n_2443),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2530)
);

NAND4xp25_ASAP7_75t_L g2531 ( 
.A(n_2459),
.B(n_283),
.C(n_281),
.D(n_282),
.Y(n_2531)
);

NOR3x1_ASAP7_75t_L g2532 ( 
.A(n_2480),
.B(n_282),
.C(n_283),
.Y(n_2532)
);

AND4x2_ASAP7_75t_L g2533 ( 
.A(n_2465),
.B(n_286),
.C(n_284),
.D(n_285),
.Y(n_2533)
);

NOR3xp33_ASAP7_75t_L g2534 ( 
.A(n_2463),
.B(n_284),
.C(n_285),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_SL g2535 ( 
.A(n_2447),
.B(n_287),
.Y(n_2535)
);

NOR3xp33_ASAP7_75t_L g2536 ( 
.A(n_2463),
.B(n_288),
.C(n_289),
.Y(n_2536)
);

OAI211xp5_ASAP7_75t_SL g2537 ( 
.A1(n_2463),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_2537)
);

NAND3x1_ASAP7_75t_L g2538 ( 
.A(n_2470),
.B(n_290),
.C(n_291),
.Y(n_2538)
);

NAND5xp2_ASAP7_75t_L g2539 ( 
.A(n_2449),
.B(n_294),
.C(n_292),
.D(n_293),
.E(n_295),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2470),
.B(n_292),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2455),
.B(n_2139),
.Y(n_2541)
);

NAND3xp33_ASAP7_75t_SL g2542 ( 
.A(n_2461),
.B(n_293),
.C(n_294),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_R g2543 ( 
.A(n_2516),
.B(n_295),
.Y(n_2543)
);

OAI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2535),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2482),
.B(n_2139),
.Y(n_2545)
);

NAND2xp33_ASAP7_75t_SL g2546 ( 
.A(n_2493),
.B(n_296),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2514),
.B(n_297),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2533),
.Y(n_2548)
);

AOI22xp33_ASAP7_75t_SL g2549 ( 
.A1(n_2500),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2511),
.B(n_299),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2503),
.Y(n_2551)
);

AOI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2484),
.A2(n_2018),
.B1(n_2081),
.B2(n_2142),
.Y(n_2552)
);

BUFx3_ASAP7_75t_L g2553 ( 
.A(n_2518),
.Y(n_2553)
);

AOI221xp5_ASAP7_75t_L g2554 ( 
.A1(n_2507),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.C(n_303),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2489),
.A2(n_2017),
.B1(n_305),
.B2(n_302),
.Y(n_2555)
);

INVxp67_ASAP7_75t_L g2556 ( 
.A(n_2539),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2505),
.B(n_304),
.Y(n_2557)
);

OAI211xp5_ASAP7_75t_L g2558 ( 
.A1(n_2506),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_2558)
);

AOI211xp5_ASAP7_75t_L g2559 ( 
.A1(n_2502),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_2559)
);

AOI22x1_ASAP7_75t_L g2560 ( 
.A1(n_2497),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_2560)
);

NAND2xp33_ASAP7_75t_L g2561 ( 
.A(n_2528),
.B(n_309),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2485),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_2562)
);

AOI322xp5_ASAP7_75t_L g2563 ( 
.A1(n_2491),
.A2(n_311),
.A3(n_312),
.B1(n_313),
.B2(n_314),
.C1(n_315),
.C2(n_316),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2526),
.A2(n_2540),
.B(n_2488),
.Y(n_2564)
);

BUFx2_ASAP7_75t_L g2565 ( 
.A(n_2538),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2537),
.B(n_313),
.Y(n_2566)
);

OAI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2525),
.A2(n_316),
.B(n_317),
.Y(n_2567)
);

NOR2x1_ASAP7_75t_L g2568 ( 
.A(n_2542),
.B(n_318),
.Y(n_2568)
);

NOR2x1_ASAP7_75t_L g2569 ( 
.A(n_2519),
.B(n_318),
.Y(n_2569)
);

OAI332xp33_ASAP7_75t_L g2570 ( 
.A1(n_2495),
.A2(n_319),
.A3(n_320),
.B1(n_321),
.B2(n_322),
.B3(n_323),
.C1(n_324),
.C2(n_325),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2512),
.Y(n_2571)
);

O2A1O1Ixp33_ASAP7_75t_L g2572 ( 
.A1(n_2530),
.A2(n_322),
.B(n_319),
.C(n_321),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2486),
.B(n_324),
.Y(n_2573)
);

O2A1O1Ixp33_ASAP7_75t_L g2574 ( 
.A1(n_2501),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_2574)
);

INVxp67_ASAP7_75t_L g2575 ( 
.A(n_2504),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_2534),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2541),
.B(n_328),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2496),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2517),
.B(n_329),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2492),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2508),
.A2(n_330),
.B(n_331),
.Y(n_2581)
);

OAI211xp5_ASAP7_75t_L g2582 ( 
.A1(n_2498),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_2582)
);

NAND4xp25_ASAP7_75t_L g2583 ( 
.A(n_2481),
.B(n_334),
.C(n_332),
.D(n_333),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_R g2584 ( 
.A(n_2487),
.B(n_334),
.Y(n_2584)
);

AOI21xp33_ASAP7_75t_L g2585 ( 
.A1(n_2520),
.A2(n_335),
.B(n_336),
.Y(n_2585)
);

NOR2x1_ASAP7_75t_L g2586 ( 
.A(n_2490),
.B(n_336),
.Y(n_2586)
);

O2A1O1Ixp33_ASAP7_75t_L g2587 ( 
.A1(n_2536),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_2587)
);

INVx2_ASAP7_75t_SL g2588 ( 
.A(n_2523),
.Y(n_2588)
);

OAI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2529),
.A2(n_339),
.B(n_341),
.Y(n_2589)
);

AOI221xp5_ASAP7_75t_L g2590 ( 
.A1(n_2524),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.C(n_344),
.Y(n_2590)
);

OAI21xp5_ASAP7_75t_SL g2591 ( 
.A1(n_2483),
.A2(n_342),
.B(n_345),
.Y(n_2591)
);

NOR2xp67_ASAP7_75t_L g2592 ( 
.A(n_2513),
.B(n_345),
.Y(n_2592)
);

HB1xp67_ASAP7_75t_L g2593 ( 
.A(n_2532),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2499),
.B(n_346),
.Y(n_2594)
);

NAND4xp25_ASAP7_75t_L g2595 ( 
.A(n_2521),
.B(n_348),
.C(n_346),
.D(n_347),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2494),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2509),
.B(n_347),
.Y(n_2597)
);

NOR3xp33_ASAP7_75t_L g2598 ( 
.A(n_2527),
.B(n_348),
.C(n_349),
.Y(n_2598)
);

AOI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2531),
.A2(n_351),
.B(n_352),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2509),
.B(n_351),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2515),
.Y(n_2601)
);

OR2x2_ASAP7_75t_L g2602 ( 
.A(n_2522),
.B(n_352),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2510),
.Y(n_2603)
);

AOI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2500),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.C(n_356),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2533),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_R g2606 ( 
.A(n_2516),
.B(n_355),
.Y(n_2606)
);

NAND3xp33_ASAP7_75t_L g2607 ( 
.A(n_2485),
.B(n_357),
.C(n_359),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2497),
.Y(n_2608)
);

NOR3xp33_ASAP7_75t_L g2609 ( 
.A(n_2500),
.B(n_361),
.C(n_362),
.Y(n_2609)
);

XOR2xp5_ASAP7_75t_L g2610 ( 
.A(n_2608),
.B(n_361),
.Y(n_2610)
);

NAND4xp75_ASAP7_75t_L g2611 ( 
.A(n_2569),
.B(n_364),
.C(n_362),
.D(n_363),
.Y(n_2611)
);

NAND4xp75_ASAP7_75t_L g2612 ( 
.A(n_2550),
.B(n_2568),
.C(n_2564),
.D(n_2573),
.Y(n_2612)
);

NAND2x1p5_ASAP7_75t_L g2613 ( 
.A(n_2551),
.B(n_2565),
.Y(n_2613)
);

NAND3x1_ASAP7_75t_L g2614 ( 
.A(n_2609),
.B(n_364),
.C(n_365),
.Y(n_2614)
);

NAND2x1p5_ASAP7_75t_L g2615 ( 
.A(n_2588),
.B(n_365),
.Y(n_2615)
);

XOR2xp5_ASAP7_75t_L g2616 ( 
.A(n_2583),
.B(n_2595),
.Y(n_2616)
);

CKINVDCx20_ASAP7_75t_R g2617 ( 
.A(n_2546),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2547),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2598),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2560),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2597),
.Y(n_2621)
);

NAND4xp75_ASAP7_75t_L g2622 ( 
.A(n_2586),
.B(n_2592),
.C(n_2557),
.D(n_2600),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_2570),
.B(n_368),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2577),
.Y(n_2624)
);

NAND4xp75_ASAP7_75t_L g2625 ( 
.A(n_2567),
.B(n_371),
.C(n_369),
.D(n_370),
.Y(n_2625)
);

NOR3xp33_ASAP7_75t_L g2626 ( 
.A(n_2571),
.B(n_370),
.C(n_371),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_L g2627 ( 
.A(n_2556),
.B(n_372),
.C(n_373),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2599),
.Y(n_2628)
);

XNOR2xp5_ASAP7_75t_L g2629 ( 
.A(n_2559),
.B(n_372),
.Y(n_2629)
);

XNOR2xp5_ASAP7_75t_L g2630 ( 
.A(n_2593),
.B(n_373),
.Y(n_2630)
);

AOI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2566),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2554),
.B(n_375),
.Y(n_2632)
);

NAND4xp75_ASAP7_75t_L g2633 ( 
.A(n_2594),
.B(n_378),
.C(n_376),
.D(n_377),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2561),
.Y(n_2634)
);

INVxp33_ASAP7_75t_L g2635 ( 
.A(n_2543),
.Y(n_2635)
);

XOR2xp5_ASAP7_75t_L g2636 ( 
.A(n_2578),
.B(n_377),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2549),
.B(n_378),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2545),
.Y(n_2638)
);

AND2x4_ASAP7_75t_L g2639 ( 
.A(n_2553),
.B(n_379),
.Y(n_2639)
);

NAND2x1p5_ASAP7_75t_SL g2640 ( 
.A(n_2606),
.B(n_379),
.Y(n_2640)
);

NAND4xp75_ASAP7_75t_L g2641 ( 
.A(n_2548),
.B(n_382),
.C(n_380),
.D(n_381),
.Y(n_2641)
);

NAND4xp75_ASAP7_75t_L g2642 ( 
.A(n_2605),
.B(n_382),
.C(n_380),
.D(n_381),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2602),
.Y(n_2643)
);

BUFx12f_ASAP7_75t_L g2644 ( 
.A(n_2596),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2587),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2579),
.Y(n_2646)
);

NAND2xp33_ASAP7_75t_L g2647 ( 
.A(n_2584),
.B(n_383),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2589),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2596),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2607),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2544),
.B(n_383),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2581),
.B(n_384),
.Y(n_2652)
);

XNOR2xp5_ASAP7_75t_L g2653 ( 
.A(n_2562),
.B(n_384),
.Y(n_2653)
);

AND2x2_ASAP7_75t_SL g2654 ( 
.A(n_2576),
.B(n_385),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2604),
.B(n_385),
.Y(n_2655)
);

CKINVDCx16_ASAP7_75t_R g2656 ( 
.A(n_2596),
.Y(n_2656)
);

NOR2x1_ASAP7_75t_L g2657 ( 
.A(n_2582),
.B(n_386),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2572),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2601),
.B(n_386),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2591),
.A2(n_2558),
.B1(n_2590),
.B2(n_2575),
.Y(n_2660)
);

NOR2xp67_ASAP7_75t_L g2661 ( 
.A(n_2603),
.B(n_387),
.Y(n_2661)
);

XNOR2xp5_ASAP7_75t_L g2662 ( 
.A(n_2580),
.B(n_387),
.Y(n_2662)
);

XOR2xp5_ASAP7_75t_L g2663 ( 
.A(n_2555),
.B(n_388),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2574),
.B(n_388),
.Y(n_2664)
);

NAND2xp33_ASAP7_75t_L g2665 ( 
.A(n_2585),
.B(n_389),
.Y(n_2665)
);

AND3x4_ASAP7_75t_L g2666 ( 
.A(n_2563),
.B(n_389),
.C(n_390),
.Y(n_2666)
);

AND2x2_ASAP7_75t_SL g2667 ( 
.A(n_2552),
.B(n_390),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2547),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2547),
.Y(n_2669)
);

XNOR2xp5_ASAP7_75t_L g2670 ( 
.A(n_2608),
.B(n_391),
.Y(n_2670)
);

XNOR2xp5_ASAP7_75t_L g2671 ( 
.A(n_2608),
.B(n_392),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2630),
.B(n_393),
.Y(n_2672)
);

NAND4xp75_ASAP7_75t_L g2673 ( 
.A(n_2659),
.B(n_2661),
.C(n_2657),
.D(n_2634),
.Y(n_2673)
);

AOI221xp5_ASAP7_75t_L g2674 ( 
.A1(n_2623),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.C(n_396),
.Y(n_2674)
);

NOR4xp75_ASAP7_75t_L g2675 ( 
.A(n_2612),
.B(n_394),
.C(n_396),
.D(n_397),
.Y(n_2675)
);

BUFx2_ASAP7_75t_L g2676 ( 
.A(n_2615),
.Y(n_2676)
);

AND2x4_ASAP7_75t_L g2677 ( 
.A(n_2624),
.B(n_397),
.Y(n_2677)
);

NOR3xp33_ASAP7_75t_SL g2678 ( 
.A(n_2656),
.B(n_398),
.C(n_400),
.Y(n_2678)
);

NOR4xp75_ASAP7_75t_SL g2679 ( 
.A(n_2614),
.B(n_398),
.C(n_400),
.D(n_401),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2610),
.Y(n_2680)
);

NOR3xp33_ASAP7_75t_L g2681 ( 
.A(n_2638),
.B(n_401),
.C(n_402),
.Y(n_2681)
);

NOR3xp33_ASAP7_75t_L g2682 ( 
.A(n_2647),
.B(n_402),
.C(n_403),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2670),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2671),
.Y(n_2684)
);

NOR5xp2_ASAP7_75t_L g2685 ( 
.A(n_2648),
.B(n_404),
.C(n_405),
.D(n_406),
.E(n_407),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_L g2686 ( 
.A(n_2660),
.B(n_2619),
.C(n_2637),
.D(n_2651),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2636),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2620),
.B(n_404),
.Y(n_2688)
);

AO211x2_ASAP7_75t_L g2689 ( 
.A1(n_2658),
.A2(n_405),
.B(n_406),
.C(n_407),
.Y(n_2689)
);

NAND4xp25_ASAP7_75t_L g2690 ( 
.A(n_2631),
.B(n_408),
.C(n_409),
.D(n_410),
.Y(n_2690)
);

NAND4xp25_ASAP7_75t_L g2691 ( 
.A(n_2649),
.B(n_408),
.C(n_411),
.D(n_412),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2611),
.Y(n_2692)
);

NOR2xp67_ASAP7_75t_L g2693 ( 
.A(n_2628),
.B(n_411),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2633),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2652),
.B(n_413),
.Y(n_2695)
);

NOR4xp25_ASAP7_75t_L g2696 ( 
.A(n_2665),
.B(n_414),
.C(n_415),
.D(n_416),
.Y(n_2696)
);

NOR4xp25_ASAP7_75t_L g2697 ( 
.A(n_2645),
.B(n_414),
.C(n_415),
.D(n_416),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2625),
.B(n_417),
.Y(n_2698)
);

AOI211xp5_ASAP7_75t_L g2699 ( 
.A1(n_2635),
.A2(n_417),
.B(n_418),
.C(n_419),
.Y(n_2699)
);

NAND5xp2_ASAP7_75t_L g2700 ( 
.A(n_2613),
.B(n_420),
.C(n_421),
.D(n_422),
.E(n_423),
.Y(n_2700)
);

AOI211xp5_ASAP7_75t_SL g2701 ( 
.A1(n_2650),
.A2(n_2617),
.B(n_2668),
.C(n_2669),
.Y(n_2701)
);

NOR3xp33_ASAP7_75t_SL g2702 ( 
.A(n_2622),
.B(n_420),
.C(n_422),
.Y(n_2702)
);

NOR4xp25_ASAP7_75t_L g2703 ( 
.A(n_2632),
.B(n_423),
.C(n_424),
.D(n_425),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2662),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2639),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2627),
.B(n_424),
.Y(n_2706)
);

NOR4xp25_ASAP7_75t_L g2707 ( 
.A(n_2618),
.B(n_425),
.C(n_426),
.D(n_427),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2626),
.B(n_426),
.Y(n_2708)
);

NOR3xp33_ASAP7_75t_L g2709 ( 
.A(n_2646),
.B(n_427),
.C(n_428),
.Y(n_2709)
);

NOR4xp75_ASAP7_75t_L g2710 ( 
.A(n_2655),
.B(n_2664),
.C(n_2641),
.D(n_2642),
.Y(n_2710)
);

XNOR2xp5_ASAP7_75t_L g2711 ( 
.A(n_2616),
.B(n_429),
.Y(n_2711)
);

XNOR2x1_ASAP7_75t_L g2712 ( 
.A(n_2666),
.B(n_430),
.Y(n_2712)
);

NAND3xp33_ASAP7_75t_SL g2713 ( 
.A(n_2643),
.B(n_430),
.C(n_431),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2640),
.B(n_432),
.Y(n_2714)
);

OR3x1_ASAP7_75t_L g2715 ( 
.A(n_2621),
.B(n_2629),
.C(n_2653),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2676),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2700),
.B(n_2652),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2687),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2693),
.B(n_2654),
.Y(n_2719)
);

OAI322xp33_ASAP7_75t_L g2720 ( 
.A1(n_2714),
.A2(n_2663),
.A3(n_2667),
.B1(n_2644),
.B2(n_2639),
.C1(n_438),
.C2(n_439),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2680),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2683),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2684),
.Y(n_2723)
);

BUFx4f_ASAP7_75t_SL g2724 ( 
.A(n_2704),
.Y(n_2724)
);

INVx1_ASAP7_75t_SL g2725 ( 
.A(n_2675),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2697),
.B(n_432),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2705),
.Y(n_2727)
);

INVx1_ASAP7_75t_SL g2728 ( 
.A(n_2677),
.Y(n_2728)
);

INVxp67_ASAP7_75t_L g2729 ( 
.A(n_2698),
.Y(n_2729)
);

CKINVDCx16_ASAP7_75t_R g2730 ( 
.A(n_2695),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2692),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2695),
.B(n_433),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2694),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_2678),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2672),
.Y(n_2735)
);

OAI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2712),
.A2(n_434),
.B(n_437),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2677),
.Y(n_2737)
);

INVx1_ASAP7_75t_SL g2738 ( 
.A(n_2688),
.Y(n_2738)
);

NAND2x1p5_ASAP7_75t_L g2739 ( 
.A(n_2688),
.B(n_434),
.Y(n_2739)
);

CKINVDCx16_ASAP7_75t_R g2740 ( 
.A(n_2696),
.Y(n_2740)
);

AOI221x1_ASAP7_75t_L g2741 ( 
.A1(n_2686),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.C(n_440),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2702),
.Y(n_2742)
);

HB1xp67_ASAP7_75t_L g2743 ( 
.A(n_2689),
.Y(n_2743)
);

INVx1_ASAP7_75t_SL g2744 ( 
.A(n_2711),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2706),
.Y(n_2745)
);

INVx1_ASAP7_75t_SL g2746 ( 
.A(n_2673),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2707),
.Y(n_2747)
);

OAI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2674),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_2748)
);

BUFx2_ASAP7_75t_L g2749 ( 
.A(n_2691),
.Y(n_2749)
);

AOI22x1_ASAP7_75t_L g2750 ( 
.A1(n_2701),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_2750)
);

AOI32xp33_ASAP7_75t_L g2751 ( 
.A1(n_2746),
.A2(n_2682),
.A3(n_2708),
.B1(n_2681),
.B2(n_2709),
.Y(n_2751)
);

AOI322xp5_ASAP7_75t_L g2752 ( 
.A1(n_2725),
.A2(n_2713),
.A3(n_2679),
.B1(n_2710),
.B2(n_2703),
.C1(n_2715),
.C2(n_2685),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2730),
.B(n_2699),
.Y(n_2753)
);

OAI211xp5_ASAP7_75t_L g2754 ( 
.A1(n_2736),
.A2(n_2690),
.B(n_445),
.C(n_446),
.Y(n_2754)
);

INVx1_ASAP7_75t_SL g2755 ( 
.A(n_2726),
.Y(n_2755)
);

OAI221xp5_ASAP7_75t_L g2756 ( 
.A1(n_2750),
.A2(n_444),
.B1(n_445),
.B2(n_447),
.C(n_448),
.Y(n_2756)
);

OAI221xp5_ASAP7_75t_L g2757 ( 
.A1(n_2748),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.C(n_450),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2743),
.B(n_2042),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2739),
.Y(n_2759)
);

OAI221xp5_ASAP7_75t_L g2760 ( 
.A1(n_2747),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.C(n_452),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2732),
.B(n_453),
.Y(n_2761)
);

A2O1A1Ixp33_ASAP7_75t_SL g2762 ( 
.A1(n_2729),
.A2(n_453),
.B(n_454),
.C(n_455),
.Y(n_2762)
);

OAI221xp5_ASAP7_75t_L g2763 ( 
.A1(n_2738),
.A2(n_454),
.B1(n_456),
.B2(n_457),
.C(n_458),
.Y(n_2763)
);

AOI322xp5_ASAP7_75t_L g2764 ( 
.A1(n_2744),
.A2(n_456),
.A3(n_457),
.B1(n_458),
.B2(n_459),
.C1(n_460),
.C2(n_461),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2740),
.B(n_2042),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2717),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2716),
.A2(n_461),
.B1(n_463),
.B2(n_465),
.Y(n_2767)
);

AOI32xp33_ASAP7_75t_L g2768 ( 
.A1(n_2728),
.A2(n_463),
.A3(n_466),
.B1(n_467),
.B2(n_468),
.Y(n_2768)
);

AOI322xp5_ASAP7_75t_L g2769 ( 
.A1(n_2734),
.A2(n_467),
.A3(n_468),
.B1(n_469),
.B2(n_470),
.C1(n_472),
.C2(n_473),
.Y(n_2769)
);

AOI322xp5_ASAP7_75t_L g2770 ( 
.A1(n_2719),
.A2(n_469),
.A3(n_470),
.B1(n_472),
.B2(n_473),
.C1(n_474),
.C2(n_475),
.Y(n_2770)
);

OAI211xp5_ASAP7_75t_SL g2771 ( 
.A1(n_2737),
.A2(n_474),
.B(n_476),
.C(n_477),
.Y(n_2771)
);

NOR2x1p5_ASAP7_75t_L g2772 ( 
.A(n_2742),
.B(n_476),
.Y(n_2772)
);

AOI221x1_ASAP7_75t_L g2773 ( 
.A1(n_2733),
.A2(n_477),
.B1(n_479),
.B2(n_480),
.C(n_481),
.Y(n_2773)
);

A2O1A1Ixp33_ASAP7_75t_L g2774 ( 
.A1(n_2727),
.A2(n_479),
.B(n_480),
.C(n_482),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_2741),
.Y(n_2775)
);

AOI322xp5_ASAP7_75t_L g2776 ( 
.A1(n_2731),
.A2(n_483),
.A3(n_484),
.B1(n_485),
.B2(n_486),
.C1(n_487),
.C2(n_488),
.Y(n_2776)
);

AOI22xp33_ASAP7_75t_L g2777 ( 
.A1(n_2766),
.A2(n_2724),
.B1(n_2733),
.B2(n_2749),
.Y(n_2777)
);

AOI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2771),
.A2(n_2722),
.B1(n_2723),
.B2(n_2718),
.Y(n_2778)
);

AND4x2_ASAP7_75t_L g2779 ( 
.A(n_2752),
.B(n_2720),
.C(n_2721),
.D(n_2733),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2765),
.A2(n_2735),
.B1(n_2745),
.B2(n_487),
.Y(n_2780)
);

HB1xp67_ASAP7_75t_L g2781 ( 
.A(n_2772),
.Y(n_2781)
);

BUFx2_ASAP7_75t_L g2782 ( 
.A(n_2775),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_2753),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2761),
.Y(n_2784)
);

AO22x2_ASAP7_75t_L g2785 ( 
.A1(n_2759),
.A2(n_484),
.B1(n_485),
.B2(n_488),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2755),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2756),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2754),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2760),
.Y(n_2789)
);

OAI22x1_ASAP7_75t_L g2790 ( 
.A1(n_2767),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_2790)
);

NAND4xp25_ASAP7_75t_L g2791 ( 
.A(n_2751),
.B(n_492),
.C(n_493),
.D(n_494),
.Y(n_2791)
);

OR2x6_ASAP7_75t_L g2792 ( 
.A(n_2782),
.B(n_2774),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2781),
.B(n_2757),
.Y(n_2793)
);

OAI221xp5_ASAP7_75t_L g2794 ( 
.A1(n_2780),
.A2(n_2762),
.B1(n_2768),
.B2(n_2763),
.C(n_2758),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2783),
.A2(n_2773),
.B1(n_2764),
.B2(n_2769),
.Y(n_2795)
);

NAND3xp33_ASAP7_75t_SL g2796 ( 
.A(n_2777),
.B(n_2776),
.C(n_2770),
.Y(n_2796)
);

OAI221xp5_ASAP7_75t_L g2797 ( 
.A1(n_2778),
.A2(n_494),
.B1(n_495),
.B2(n_496),
.C(n_497),
.Y(n_2797)
);

NAND3xp33_ASAP7_75t_L g2798 ( 
.A(n_2788),
.B(n_495),
.C(n_497),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2790),
.B(n_498),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2787),
.A2(n_499),
.B1(n_501),
.B2(n_502),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2779),
.Y(n_2801)
);

OAI22x1_ASAP7_75t_L g2802 ( 
.A1(n_2795),
.A2(n_2801),
.B1(n_2789),
.B2(n_2784),
.Y(n_2802)
);

NAND4xp75_ASAP7_75t_L g2803 ( 
.A(n_2793),
.B(n_2786),
.C(n_2791),
.D(n_2785),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2799),
.B(n_2785),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2798),
.B(n_499),
.Y(n_2805)
);

OA21x2_ASAP7_75t_L g2806 ( 
.A1(n_2794),
.A2(n_501),
.B(n_502),
.Y(n_2806)
);

XOR2xp5_ASAP7_75t_L g2807 ( 
.A(n_2796),
.B(n_503),
.Y(n_2807)
);

AO22x2_ASAP7_75t_L g2808 ( 
.A1(n_2792),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2800),
.B(n_504),
.Y(n_2809)
);

AOI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2807),
.A2(n_2797),
.B1(n_506),
.B2(n_507),
.Y(n_2810)
);

OAI22x1_ASAP7_75t_L g2811 ( 
.A1(n_2806),
.A2(n_505),
.B1(n_507),
.B2(n_508),
.Y(n_2811)
);

OAI22x1_ASAP7_75t_SL g2812 ( 
.A1(n_2802),
.A2(n_2803),
.B1(n_2804),
.B2(n_2805),
.Y(n_2812)
);

OAI31xp33_ASAP7_75t_SL g2813 ( 
.A1(n_2809),
.A2(n_508),
.A3(n_510),
.B(n_511),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_SL g2814 ( 
.A1(n_2808),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_2814)
);

OAI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2807),
.A2(n_512),
.B(n_513),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2807),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2813),
.B(n_515),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2815),
.B(n_2811),
.Y(n_2818)
);

OAI21x1_ASAP7_75t_L g2819 ( 
.A1(n_2816),
.A2(n_515),
.B(n_516),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2817),
.B(n_2810),
.Y(n_2820)
);

AOI22xp33_ASAP7_75t_L g2821 ( 
.A1(n_2818),
.A2(n_2814),
.B1(n_2812),
.B2(n_519),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2819),
.Y(n_2822)
);

AOI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2818),
.A2(n_516),
.B(n_518),
.Y(n_2823)
);

AOI22x1_ASAP7_75t_L g2824 ( 
.A1(n_2822),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.Y(n_2824)
);

OAI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2821),
.A2(n_520),
.B1(n_523),
.B2(n_524),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_SL g2826 ( 
.A(n_2825),
.B(n_2820),
.Y(n_2826)
);

OAI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2824),
.A2(n_2823),
.B(n_527),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_2826),
.Y(n_2828)
);

AOI221xp5_ASAP7_75t_L g2829 ( 
.A1(n_2828),
.A2(n_2827),
.B1(n_527),
.B2(n_528),
.C(n_529),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2829),
.A2(n_526),
.B(n_528),
.Y(n_2830)
);

AOI211xp5_ASAP7_75t_L g2831 ( 
.A1(n_2830),
.A2(n_530),
.B(n_531),
.C(n_532),
.Y(n_2831)
);


endmodule