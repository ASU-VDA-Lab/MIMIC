module fake_jpeg_10639_n_191 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx8_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_30),
.B1(n_32),
.B2(n_29),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_41),
.B1(n_33),
.B2(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_19),
.B1(n_18),
.B2(n_12),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_12),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_24),
.B(n_21),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_16),
.B1(n_15),
.B2(n_22),
.Y(n_48)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_43),
.B1(n_63),
.B2(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_17),
.B1(n_14),
.B2(n_3),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_44),
.C(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_52),
.B1(n_42),
.B2(n_45),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_43),
.C(n_42),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_55),
.C(n_53),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_58),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_61),
.B1(n_38),
.B2(n_49),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_60),
.B1(n_45),
.B2(n_48),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_48),
.B(n_41),
.C(n_37),
.D(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_87),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_52),
.B(n_48),
.C(n_51),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_96),
.B1(n_65),
.B2(n_75),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_70),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_60),
.B1(n_48),
.B2(n_42),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_81),
.B(n_74),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_98),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_36),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_36),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_82),
.B(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_89),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_86),
.C(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_122),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_96),
.B1(n_97),
.B2(n_93),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_116),
.B1(n_125),
.B2(n_129),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_89),
.B(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_104),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_17),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_127),
.C(n_106),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_1),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_112),
.B1(n_99),
.B2(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_111),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_119),
.B1(n_122),
.B2(n_102),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_121),
.C(n_127),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_153),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_137),
.B(n_142),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.C(n_5),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_140),
.B1(n_149),
.B2(n_148),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_147),
.C(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_1),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_3),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_161),
.B(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_4),
.B(n_7),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_4),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_167),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_182),
.B(n_176),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_8),
.C(n_9),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_8),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_184),
.B(n_185),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_178),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_186),
.C(n_174),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_8),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_189),
.A2(n_9),
.B(n_10),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_10),
.C(n_11),
.Y(n_191)
);


endmodule