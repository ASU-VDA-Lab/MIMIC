module fake_jpeg_21032_n_358 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_45),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_62),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_51),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_17),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_2),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_27),
.Y(n_112)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_85),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_35),
.B1(n_26),
.B2(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_91),
.Y(n_138)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_78),
.A2(n_110),
.B1(n_7),
.B2(n_8),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_82),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_22),
.B(n_39),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_35),
.B1(n_41),
.B2(n_24),
.Y(n_84)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_113),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_35),
.B1(n_41),
.B2(n_24),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_20),
.B1(n_39),
.B2(n_33),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_151)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_25),
.B1(n_36),
.B2(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_46),
.B(n_19),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_40),
.B1(n_19),
.B2(n_29),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_112),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_27),
.B1(n_38),
.B2(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_43),
.B(n_27),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_7),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_7),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_53),
.B1(n_38),
.B2(n_9),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_136),
.Y(n_158)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_63),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_139),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_58),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_149),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_78),
.A2(n_63),
.B(n_8),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_112),
.B(n_88),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_77),
.B(n_71),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_88),
.Y(n_161)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_71),
.B(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_153),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_16),
.B1(n_11),
.B2(n_12),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_15),
.B(n_16),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_70),
.B1(n_117),
.B2(n_75),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_68),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_78),
.B(n_14),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_161),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_144),
.B(n_124),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_166),
.B(n_161),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_110),
.B(n_86),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_76),
.B1(n_85),
.B2(n_103),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_172),
.B1(n_176),
.B2(n_179),
.Y(n_205)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_103),
.B1(n_76),
.B2(n_93),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_110),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_117),
.B1(n_70),
.B2(n_68),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_119),
.A2(n_69),
.B1(n_72),
.B2(n_89),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_72),
.B1(n_97),
.B2(n_82),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_138),
.B1(n_149),
.B2(n_132),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_97),
.B1(n_79),
.B2(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_118),
.B(n_101),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_193),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_131),
.A2(n_106),
.B1(n_81),
.B2(n_101),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_189),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_106),
.B1(n_15),
.B2(n_16),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_145),
.A2(n_15),
.B1(n_140),
.B2(n_136),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_135),
.A2(n_118),
.B1(n_153),
.B2(n_134),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_200),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_215),
.B(n_224),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_152),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_165),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_150),
.C(n_122),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_223),
.C(n_187),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_158),
.B(n_144),
.Y(n_208)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_123),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_156),
.B(n_160),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_220),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_218),
.B1(n_204),
.B2(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_123),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_120),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_124),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_184),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_193),
.Y(n_247)
);

BUFx12f_ASAP7_75t_SL g226 ( 
.A(n_164),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_227),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_142),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_246),
.B1(n_255),
.B2(n_213),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_162),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_244),
.Y(n_258)
);

OAI211xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_174),
.B(n_163),
.C(n_161),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_241),
.B(n_224),
.Y(n_270)
);

XOR2x2_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_191),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_243),
.B(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_162),
.B1(n_173),
.B2(n_190),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_173),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_204),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_181),
.C(n_183),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_199),
.C(n_228),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_220),
.B(n_147),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_195),
.A2(n_186),
.B1(n_177),
.B2(n_154),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_272),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_235),
.A2(n_224),
.B(n_196),
.C(n_201),
.Y(n_261)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_197),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_263),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_202),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_198),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_199),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_270),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_206),
.B(n_217),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_280),
.B(n_239),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_213),
.B(n_205),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_279),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_250),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_237),
.A2(n_216),
.B1(n_221),
.B2(n_219),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_240),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_239),
.A2(n_155),
.B(n_222),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_285),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_239),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_282),
.A2(n_293),
.B(n_209),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_274),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_249),
.C(n_254),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_294),
.C(n_298),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_297),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_252),
.B1(n_221),
.B2(n_194),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_296),
.B(n_261),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_233),
.C(n_244),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_253),
.C(n_232),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_230),
.C(n_251),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_280),
.C(n_272),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_278),
.B1(n_242),
.B2(n_266),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_306),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_265),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_313),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_314),
.B(n_289),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_261),
.B(n_270),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_291),
.B(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_309),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_275),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_311),
.C(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_259),
.C(n_257),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_276),
.B1(n_230),
.B2(n_245),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_285),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_271),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_242),
.B(n_252),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_315),
.A2(n_282),
.B1(n_284),
.B2(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_316),
.B(n_319),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_286),
.C(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_324),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_288),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_327),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_284),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_315),
.B(n_310),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_335),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_334),
.A2(n_336),
.B(n_337),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_313),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_303),
.B(n_312),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_286),
.C(n_302),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_331),
.B(n_316),
.Y(n_339)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_337),
.B(n_318),
.CI(n_317),
.CON(n_340),
.SN(n_340)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_341),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_188),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_330),
.A2(n_325),
.B1(n_318),
.B2(n_303),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_345),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_147),
.C(n_129),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_329),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_346),
.A2(n_194),
.B(n_125),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_129),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_347),
.B(n_345),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_344),
.C(n_349),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_350),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_352),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_354),
.A2(n_355),
.B(n_353),
.C(n_351),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_356),
.Y(n_358)
);


endmodule