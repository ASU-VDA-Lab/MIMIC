module fake_aes_1040_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_22;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_7), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_0), .Y(n_13) );
CKINVDCx14_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .B1(n_12), .B2(n_11), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_1), .Y(n_18) );
XOR2xp5_ASAP7_75t_L g19 ( .A(n_18), .B(n_2), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_10), .B1(n_4), .B2(n_6), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
endmodule