module fake_jpeg_15829_n_24 (n_3, n_2, n_1, n_0, n_4, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_1),
.C(n_4),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_0),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_0),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_2),
.B1(n_10),
.B2(n_8),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_16),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_12),
.C(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_9),
.B1(n_11),
.B2(n_19),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_21),
.C(n_22),
.Y(n_24)
);


endmodule