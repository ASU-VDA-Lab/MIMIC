module real_jpeg_26662_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_56),
.Y(n_93)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_1),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_1),
.A2(n_29),
.B(n_33),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_1),
.B(n_31),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_62),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_62),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_76),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_1),
.A2(n_92),
.B1(n_96),
.B2(n_258),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_1),
.A2(n_32),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_104),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_104),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_104),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_5),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_135),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_135),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_135),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_9),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_9),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_10),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_177),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_177),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_177),
.Y(n_258)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_11),
.A2(n_57),
.A3(n_62),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_12),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_166),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_166),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_166),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_13),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_102),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_102),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_102),
.Y(n_247)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_16),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_16),
.A2(n_27),
.B1(n_62),
.B2(n_63),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_16),
.A2(n_27),
.B1(n_56),
.B2(n_57),
.Y(n_127)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_22),
.B(n_43),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_24),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_26),
.A2(n_35),
.B(n_175),
.C(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_28),
.A2(n_31),
.B1(n_101),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_28),
.A2(n_31),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_28),
.A2(n_31),
.B1(n_134),
.B2(n_206),
.Y(n_220)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_31),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_32),
.A2(n_70),
.B(n_72),
.C(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_70),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_32),
.A2(n_63),
.A3(n_70),
.B1(n_275),
.B2(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_33),
.B(n_175),
.Y(n_275)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_84),
.B(n_338),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_77),
.C(n_79),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_44),
.A2(n_45),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_66),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_46),
.B(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_48),
.A2(n_81),
.B1(n_83),
.B2(n_103),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_52),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_52),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_52),
.A2(n_66),
.B1(n_144),
.B2(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_60),
.B(n_65),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_53),
.A2(n_60),
.B1(n_65),
.B2(n_113),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_60),
.B1(n_110),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_53),
.A2(n_60),
.B1(n_130),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_53),
.A2(n_60),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_53),
.A2(n_60),
.B1(n_233),
.B2(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_53),
.B(n_175),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_53),
.A2(n_60),
.B1(n_171),
.B2(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_55),
.B(n_56),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_56),
.B(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_62),
.B(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_66),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_75),
.B2(n_76),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_67),
.A2(n_68),
.B1(n_76),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_76),
.B1(n_119),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_68),
.A2(n_76),
.B1(n_165),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_68),
.A2(n_76),
.B1(n_132),
.B2(n_209),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_73),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_69),
.A2(n_73),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_69),
.A2(n_73),
.B1(n_164),
.B2(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_69),
.A2(n_73),
.B1(n_167),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_69),
.A2(n_73),
.B1(n_189),
.B2(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_70),
.Y(n_284)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_77),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_83),
.B1(n_100),
.B2(n_103),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_81),
.A2(n_83),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_331),
.B(n_337),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_147),
.A3(n_156),
.B1(n_329),
.B2(n_330),
.C(n_342),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_136),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_87),
.B(n_136),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_116),
.C(n_123),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_88),
.B(n_116),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_105),
.B1(n_106),
.B2(n_115),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_98),
.B2(n_99),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_90),
.A2(n_99),
.B(n_105),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_90),
.A2(n_91),
.B1(n_107),
.B2(n_108),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_97),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_97),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_92),
.A2(n_127),
.B1(n_128),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_92),
.A2(n_94),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_92),
.A2(n_94),
.B1(n_252),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_92),
.A2(n_128),
.B1(n_247),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_93),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_93),
.A2(n_95),
.B1(n_182),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_93),
.A2(n_95),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

INVx5_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_114),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_111),
.A2(n_114),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B(n_122),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_121),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_137),
.CI(n_146),
.CON(n_136),
.SN(n_136)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_137),
.C(n_146),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_123),
.A2(n_124),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.C(n_133),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_125),
.B(n_131),
.CI(n_133),
.CON(n_312),
.SN(n_312)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_126),
.B(n_129),
.Y(n_216)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_136),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_145),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_139),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_141),
.C(n_144),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_139),
.B(n_154),
.C(n_155),
.Y(n_332)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_148),
.B(n_149),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

AOI321xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_310),
.A3(n_318),
.B1(n_323),
.B2(n_328),
.C(n_343),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_211),
.C(n_223),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_193),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_159),
.B(n_193),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_178),
.C(n_185),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_160),
.B(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_173),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_169),
.C(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_175),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_178),
.A2(n_185),
.B1(n_186),
.B2(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_178),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_181),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_187),
.B(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_190),
.B(n_192),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_191),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_200),
.C(n_201),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_210),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_207),
.C(n_210),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_212),
.A2(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_213),
.B(n_214),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_216),
.B(n_217),
.C(n_222),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_218),
.B(n_220),
.C(n_221),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_304),
.B(n_309),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_290),
.B(n_303),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_268),
.B(n_289),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_248),
.B(n_267),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_228),
.B(n_238),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_230),
.B1(n_234),
.B2(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_243),
.C(n_245),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_244),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_246),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_255),
.B(n_266),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_265),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_270),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_281),
.B1(n_287),
.B2(n_288),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_280),
.C(n_288),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_278),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_281),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_299),
.C(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.C(n_314),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_312),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_324),
.B(n_327),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule