module fake_jpeg_24942_n_307 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_1),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_2),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_29),
.B1(n_18),
.B2(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_21),
.B1(n_33),
.B2(n_32),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_38),
.B1(n_36),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_72),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_36),
.B1(n_38),
.B2(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_24),
.C(n_35),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_37),
.C(n_21),
.Y(n_87)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_28),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_37),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_37),
.B(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_30),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_111)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_94),
.B(n_112),
.Y(n_131)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_82),
.B(n_115),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_84),
.B(n_89),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_98),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_37),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_52),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_50),
.B1(n_66),
.B2(n_8),
.Y(n_140)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_73),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_46),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_21),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_111),
.A2(n_61),
.B1(n_63),
.B2(n_56),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_57),
.A2(n_20),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_16),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_3),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_62),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_57),
.B(n_4),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_66),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_120),
.B(n_115),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_70),
.B1(n_77),
.B2(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_149),
.Y(n_159)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_56),
.B1(n_51),
.B2(n_50),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_128),
.A2(n_143),
.B1(n_100),
.B2(n_105),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_133),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_5),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_95),
.Y(n_165)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_134),
.Y(n_163)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_105),
.B1(n_96),
.B2(n_99),
.Y(n_181)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

AO22x2_ASAP7_75t_SL g143 ( 
.A1(n_80),
.A2(n_50),
.B1(n_66),
.B2(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_6),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_82),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_161),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_98),
.B(n_90),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_177),
.B(n_179),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_84),
.B(n_102),
.C(n_94),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_157),
.B(n_158),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_87),
.B(n_91),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_92),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_141),
.C(n_129),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_169),
.C(n_124),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_167),
.B(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_89),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_85),
.C(n_86),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_136),
.Y(n_184)
);

AO21x1_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_137),
.B(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_180),
.B1(n_181),
.B2(n_123),
.Y(n_198)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_85),
.B(n_86),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_83),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_124),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_183),
.C(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_184),
.B(n_186),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_121),
.C(n_135),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_135),
.Y(n_190)
);

NAND2xp33_ASAP7_75t_R g212 ( 
.A(n_190),
.B(n_193),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_121),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_206),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_127),
.B(n_99),
.Y(n_193)
);

NOR2x1_ASAP7_75t_R g197 ( 
.A(n_180),
.B(n_127),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_200),
.B(n_209),
.C(n_164),
.D(n_153),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_207),
.B1(n_175),
.B2(n_176),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_122),
.B(n_133),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_204),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_6),
.C(n_7),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_208),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_168),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_96),
.B1(n_97),
.B2(n_107),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_138),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_6),
.B(n_8),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_220),
.Y(n_245)
);

BUFx12_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_177),
.B1(n_181),
.B2(n_172),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_218),
.B1(n_222),
.B2(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

AO22x1_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_155),
.B1(n_178),
.B2(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_225),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_228),
.B(n_230),
.Y(n_237)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_167),
.B1(n_161),
.B2(n_150),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_229),
.A2(n_231),
.B1(n_198),
.B2(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_183),
.C(n_182),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_244),
.C(n_221),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_206),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_248),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_186),
.A3(n_196),
.B1(n_189),
.B2(n_209),
.C1(n_203),
.C2(n_208),
.Y(n_238)
);

OAI322xp33_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_219),
.A3(n_213),
.B1(n_223),
.B2(n_229),
.C1(n_228),
.C2(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_165),
.B1(n_191),
.B2(n_154),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_246),
.B1(n_222),
.B2(n_220),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_154),
.C(n_162),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_134),
.B1(n_126),
.B2(n_162),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_212),
.B(n_217),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_163),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_235),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_163),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_244),
.C(n_234),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_266),
.B1(n_247),
.B2(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_228),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_263),
.B(n_237),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_163),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

XOR2x2_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_227),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_11),
.B(n_12),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_242),
.B1(n_251),
.B2(n_15),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_276),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_272),
.B(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_273),
.C(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_267),
.B1(n_260),
.B2(n_265),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_13),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_284),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_286),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_268),
.B(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_253),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_259),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_291),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_274),
.B(n_14),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_16),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_13),
.B(n_14),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_15),
.B(n_16),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_292),
.C(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_286),
.C(n_302),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_299),
.B(n_297),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_303),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_305),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_304),
.Y(n_307)
);


endmodule