module real_aes_14152_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_924, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_924;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_905;
wire n_635;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g273 ( .A(n_0), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_1), .Y(n_205) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_2), .A2(n_48), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g219 ( .A(n_2), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_3), .B(n_155), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_4), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_5), .B(n_634), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_6), .B(n_312), .Y(n_587) );
AND2x2_ASAP7_75t_L g163 ( .A(n_7), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_8), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_9), .B(n_250), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_10), .B(n_250), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_11), .B(n_600), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_12), .B(n_144), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_13), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_14), .B(n_272), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_15), .Y(n_608) );
BUFx3_ASAP7_75t_L g140 ( .A(n_16), .Y(n_140) );
INVx1_ASAP7_75t_L g146 ( .A(n_16), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_17), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_18), .B(n_138), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_19), .Y(n_582) );
BUFx10_ASAP7_75t_L g559 ( .A(n_20), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_21), .B(n_226), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_22), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_23), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_24), .B(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_25), .B(n_201), .C(n_290), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_26), .B(n_226), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_27), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_28), .B(n_138), .Y(n_651) );
NAND2xp33_ASAP7_75t_L g665 ( .A(n_29), .B(n_139), .Y(n_665) );
AND2x2_ASAP7_75t_L g908 ( .A(n_30), .B(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g190 ( .A(n_31), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_32), .A2(n_142), .B(n_210), .C(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_33), .A2(n_99), .B1(n_564), .B2(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_33), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_34), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_35), .B(n_207), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_36), .B(n_155), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_37), .B(n_179), .Y(n_639) );
INVx1_ASAP7_75t_L g111 ( .A(n_38), .Y(n_111) );
AND3x2_ASAP7_75t_L g912 ( .A(n_38), .B(n_905), .C(n_906), .Y(n_912) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_39), .B(n_252), .Y(n_251) );
AO221x1_ASAP7_75t_L g688 ( .A1(n_40), .A2(n_81), .B1(n_178), .B2(n_226), .C(n_264), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_41), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_42), .B(n_209), .Y(n_208) );
AND2x4_ASAP7_75t_L g189 ( .A(n_43), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_44), .B(n_192), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_45), .B(n_132), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_46), .B(n_209), .C(n_210), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_47), .B(n_192), .Y(n_306) );
INVx1_ASAP7_75t_L g220 ( .A(n_48), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_49), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_50), .A2(n_154), .B(n_271), .C(n_274), .Y(n_270) );
INVx1_ASAP7_75t_L g134 ( .A(n_51), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_52), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g613 ( .A1(n_53), .A2(n_614), .B(n_615), .C(n_617), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_54), .B(n_192), .Y(n_213) );
INVx2_ASAP7_75t_L g616 ( .A(n_55), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_56), .B(n_132), .Y(n_589) );
AND2x4_ASAP7_75t_L g919 ( .A(n_57), .B(n_920), .Y(n_919) );
INVx3_ASAP7_75t_L g239 ( .A(n_58), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_59), .B(n_72), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_60), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g920 ( .A(n_61), .Y(n_920) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_62), .B(n_235), .Y(n_317) );
INVx1_ASAP7_75t_L g177 ( .A(n_63), .Y(n_177) );
AND2x2_ASAP7_75t_L g641 ( .A(n_64), .B(n_132), .Y(n_641) );
INVx1_ASAP7_75t_L g693 ( .A(n_65), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_66), .A2(n_94), .B1(n_119), .B2(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_66), .Y(n_119) );
INVx2_ASAP7_75t_L g109 ( .A(n_67), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_68), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_69), .B(n_203), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_70), .B(n_201), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_71), .A2(n_74), .B1(n_600), .B2(n_634), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_73), .B(n_210), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_75), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g265 ( .A(n_76), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_77), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_78), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_79), .B(n_290), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_80), .Y(n_113) );
AND2x2_ASAP7_75t_L g623 ( .A(n_82), .B(n_164), .Y(n_623) );
INVx1_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
INVx1_ASAP7_75t_L g161 ( .A(n_83), .Y(n_161) );
BUFx3_ASAP7_75t_L g174 ( .A(n_83), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_84), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g237 ( .A(n_85), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_86), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_87), .B(n_276), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_88), .B(n_143), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_89), .B(n_164), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_90), .B(n_584), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_91), .B(n_132), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_92), .B(n_315), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_93), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_94), .Y(n_120) );
INVx1_ASAP7_75t_L g225 ( .A(n_95), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_96), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_97), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_98), .A2(n_102), .B1(n_913), .B2(n_921), .Y(n_101) );
INVx1_ASAP7_75t_L g564 ( .A(n_99), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_100), .B(n_235), .Y(n_309) );
OR2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_114), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_103), .A2(n_116), .B(n_553), .Y(n_115) );
NOR2x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_113), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g556 ( .A(n_107), .Y(n_556) );
NOR2x1p5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g906 ( .A(n_109), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
BUFx2_ASAP7_75t_L g570 ( .A(n_111), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g917 ( .A(n_111), .B(n_906), .C(n_918), .Y(n_917) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_112), .Y(n_905) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_557), .B(n_560), .Y(n_114) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
XOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
AO22x2_ASAP7_75t_L g566 ( .A1(n_121), .A2(n_567), .B1(n_568), .B2(n_571), .Y(n_566) );
NAND4xp75_ASAP7_75t_L g121 ( .A(n_122), .B(n_399), .C(n_464), .D(n_512), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_357), .C(n_369), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_334), .C(n_341), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_243), .B1(n_294), .B2(n_300), .C(n_322), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_127), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_193), .Y(n_127) );
INVx1_ASAP7_75t_L g295 ( .A(n_128), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_128), .B(n_415), .Y(n_495) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_166), .Y(n_128) );
INVx1_ASAP7_75t_L g333 ( .A(n_129), .Y(n_333) );
AND2x2_ASAP7_75t_L g336 ( .A(n_129), .B(n_196), .Y(n_336) );
AND2x4_ASAP7_75t_L g392 ( .A(n_129), .B(n_195), .Y(n_392) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_135), .B(n_162), .Y(n_129) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_130), .A2(n_247), .B(n_258), .Y(n_246) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_130), .A2(n_247), .B(n_258), .Y(n_385) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2x1_ASAP7_75t_SL g319 ( .A(n_131), .B(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g356 ( .A(n_132), .Y(n_356) );
INVx2_ASAP7_75t_L g631 ( .A(n_132), .Y(n_631) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_132), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_132), .B(n_228), .Y(n_685) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
BUFx2_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
INVx1_ASAP7_75t_L g221 ( .A(n_134), .Y(n_221) );
INVx2_ASAP7_75t_L g345 ( .A(n_135), .Y(n_345) );
AOI22x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_148), .B1(n_150), .B2(n_158), .Y(n_135) );
OAI22x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B1(n_142), .B2(n_147), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
INVx2_ASAP7_75t_L g203 ( .A(n_139), .Y(n_203) );
INVx2_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
INVx2_ASAP7_75t_L g250 ( .A(n_139), .Y(n_250) );
INVx3_ASAP7_75t_L g264 ( .A(n_139), .Y(n_264) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g252 ( .A(n_144), .Y(n_252) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_144), .Y(n_267) );
INVx2_ASAP7_75t_L g287 ( .A(n_144), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_144), .B(n_608), .Y(n_607) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_145), .Y(n_226) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
INVx1_ASAP7_75t_L g274 ( .A(n_148), .Y(n_274) );
AOI21x1_ASAP7_75t_L g284 ( .A1(n_148), .A2(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_SL g632 ( .A1(n_148), .A2(n_633), .B(n_635), .Y(n_632) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B1(n_154), .B2(n_157), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVxp67_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
INVx2_ASAP7_75t_L g312 ( .A(n_156), .Y(n_312) );
INVx1_ASAP7_75t_L g316 ( .A(n_156), .Y(n_316) );
INVx1_ASAP7_75t_L g606 ( .A(n_156), .Y(n_606) );
AOI21x1_ASAP7_75t_SL g262 ( .A1(n_158), .A2(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_159), .A2(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_159), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_160), .A2(n_661), .B(n_662), .Y(n_660) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g253 ( .A(n_161), .Y(n_253) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AO31x2_ASAP7_75t_L g344 ( .A1(n_163), .A2(n_345), .A3(n_346), .B(n_347), .Y(n_344) );
AO31x2_ASAP7_75t_L g379 ( .A1(n_163), .A2(n_345), .A3(n_346), .B(n_347), .Y(n_379) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g326 ( .A(n_166), .Y(n_326) );
AND2x2_ASAP7_75t_L g337 ( .A(n_166), .B(n_215), .Y(n_337) );
INVx1_ASAP7_75t_L g376 ( .A(n_166), .Y(n_376) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_166), .Y(n_413) );
INVx3_ASAP7_75t_L g460 ( .A(n_166), .Y(n_460) );
INVx2_ASAP7_75t_L g473 ( .A(n_166), .Y(n_473) );
AND2x2_ASAP7_75t_L g511 ( .A(n_166), .B(n_214), .Y(n_511) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_191), .Y(n_167) );
OAI21x1_ASAP7_75t_L g197 ( .A1(n_168), .A2(n_198), .B(n_213), .Y(n_197) );
OAI21x1_ASAP7_75t_L g579 ( .A1(n_168), .A2(n_580), .B(n_589), .Y(n_579) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVxp67_ASAP7_75t_L g625 ( .A(n_169), .Y(n_625) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_181), .B(n_188), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_175), .Y(n_171) );
INVx2_ASAP7_75t_L g178 ( .A(n_174), .Y(n_178) );
INVx2_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_174), .B(n_228), .Y(n_227) );
NOR3xp33_ASAP7_75t_L g236 ( .A(n_174), .B(n_228), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g585 ( .A(n_174), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_179), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g609 ( .A(n_178), .Y(n_609) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g201 ( .A(n_180), .Y(n_201) );
INVx2_ASAP7_75t_L g584 ( .A(n_180), .Y(n_584) );
INVx2_ASAP7_75t_L g634 ( .A(n_180), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_186), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
INVx2_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
INVx2_ASAP7_75t_L g600 ( .A(n_185), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_186), .A2(n_200), .B(n_202), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_255), .B(n_256), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_186), .A2(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g622 ( .A(n_186), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_186), .A2(n_639), .B(n_640), .Y(n_638) );
BUFx10_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_188), .A2(n_248), .B(n_254), .Y(n_247) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_188), .A2(n_581), .B(n_586), .Y(n_580) );
BUFx6f_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g212 ( .A(n_189), .Y(n_212) );
INVx3_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
INVx1_ASAP7_75t_L g278 ( .A(n_189), .Y(n_278) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_192), .Y(n_282) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_214), .Y(n_194) );
OR2x2_ASAP7_75t_L g429 ( .A(n_195), .B(n_379), .Y(n_429) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g297 ( .A(n_196), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g327 ( .A(n_196), .Y(n_327) );
INVx2_ASAP7_75t_L g350 ( .A(n_196), .Y(n_350) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_204), .B(n_211), .Y(n_198) );
O2A1O1Ixp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_208), .C(n_210), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_206), .A2(n_653), .B(n_654), .Y(n_652) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_211), .A2(n_284), .B(n_288), .Y(n_283) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_SL g321 ( .A(n_212), .Y(n_321) );
BUFx2_ASAP7_75t_L g330 ( .A(n_214), .Y(n_330) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_214), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_214), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g427 ( .A(n_214), .Y(n_427) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_241), .Y(n_215) );
AO21x1_ASAP7_75t_L g299 ( .A1(n_216), .A2(n_222), .B(n_241), .Y(n_299) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_217), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_217), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_R g691 ( .A(n_218), .B(n_228), .Y(n_691) );
AOI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_227), .B1(n_229), .B2(n_232), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g240 ( .A(n_226), .Y(n_240) );
INVx2_ASAP7_75t_L g257 ( .A(n_226), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_228), .B(n_233), .Y(n_232) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_228), .B(n_233), .C(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g626 ( .A(n_228), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g235 ( .A(n_231), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B1(n_238), .B2(n_240), .Y(n_234) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_259), .Y(n_243) );
OR2x2_ASAP7_75t_L g339 ( .A(n_244), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g358 ( .A(n_244), .B(n_304), .Y(n_358) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_245), .B(n_383), .Y(n_389) );
BUFx3_ASAP7_75t_L g395 ( .A(n_245), .Y(n_395) );
AND2x4_ASAP7_75t_L g441 ( .A(n_245), .B(n_390), .Y(n_441) );
AND2x2_ASAP7_75t_L g504 ( .A(n_245), .B(n_398), .Y(n_504) );
AND2x2_ASAP7_75t_L g552 ( .A(n_245), .B(n_302), .Y(n_552) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_246), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_251), .B(n_253), .Y(n_248) );
INVx2_ASAP7_75t_L g318 ( .A(n_253), .Y(n_318) );
INVx1_ASAP7_75t_L g617 ( .A(n_253), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_253), .A2(n_664), .B(n_665), .Y(n_663) );
INVxp67_ASAP7_75t_L g291 ( .A(n_257), .Y(n_291) );
OR2x2_ASAP7_75t_L g434 ( .A(n_259), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g549 ( .A(n_259), .B(n_303), .Y(n_549) );
OR2x6_ASAP7_75t_L g259 ( .A(n_260), .B(n_279), .Y(n_259) );
OR2x2_ASAP7_75t_SL g353 ( .A(n_260), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g390 ( .A(n_260), .Y(n_390) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_268), .B(n_275), .Y(n_261) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OAI21xp33_ASAP7_75t_L g275 ( .A1(n_269), .A2(n_276), .B(n_278), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVxp67_ASAP7_75t_L g346 ( .A(n_276), .Y(n_346) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_277), .B(n_321), .Y(n_596) );
INVx1_ASAP7_75t_L g348 ( .A(n_278), .Y(n_348) );
AND2x2_ASAP7_75t_L g408 ( .A(n_279), .B(n_385), .Y(n_408) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_280), .Y(n_397) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_293), .Y(n_281) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_283), .A2(n_293), .B(n_355), .Y(n_354) );
O2A1O1Ixp5_ASAP7_75t_L g581 ( .A1(n_287), .A2(n_582), .B(n_583), .C(n_585), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_292), .Y(n_288) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_295), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_445) );
OR2x2_ASAP7_75t_L g458 ( .A(n_296), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g367 ( .A(n_297), .Y(n_367) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_297), .Y(n_480) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_299), .B(n_333), .Y(n_417) );
AND2x2_ASAP7_75t_L g472 ( .A(n_299), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g329 ( .A(n_302), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_302), .B(n_332), .Y(n_340) );
AND2x2_ASAP7_75t_L g360 ( .A(n_302), .B(n_354), .Y(n_360) );
AND2x4_ASAP7_75t_L g384 ( .A(n_302), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g476 ( .A(n_303), .Y(n_476) );
AND2x2_ASAP7_75t_L g508 ( .A(n_303), .B(n_390), .Y(n_508) );
NOR2xp67_ASAP7_75t_R g522 ( .A(n_303), .B(n_328), .Y(n_522) );
OR2x2_ASAP7_75t_L g528 ( .A(n_303), .B(n_326), .Y(n_528) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g325 ( .A(n_304), .Y(n_325) );
INVx2_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
BUFx2_ASAP7_75t_L g435 ( .A(n_304), .Y(n_435) );
AND2x2_ASAP7_75t_L g442 ( .A(n_304), .B(n_354), .Y(n_442) );
AND2x4_ASAP7_75t_L g456 ( .A(n_304), .B(n_332), .Y(n_456) );
OR2x2_ASAP7_75t_L g538 ( .A(n_304), .B(n_397), .Y(n_538) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2x1_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OAI21x1_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_313), .B(n_319), .Y(n_307) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
NOR5xp2_ASAP7_75t_L g323 ( .A(n_324), .B(n_328), .C(n_330), .D(n_331), .E(n_333), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .C(n_327), .Y(n_324) );
INVx2_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx2_ASAP7_75t_L g364 ( .A(n_326), .Y(n_364) );
AND2x2_ASAP7_75t_L g493 ( .A(n_326), .B(n_377), .Y(n_493) );
AND2x2_ASAP7_75t_L g377 ( .A(n_327), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g452 ( .A(n_327), .Y(n_452) );
AND2x2_ASAP7_75t_L g517 ( .A(n_327), .B(n_427), .Y(n_517) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g438 ( .A(n_329), .B(n_408), .Y(n_438) );
AND2x2_ASAP7_75t_L g469 ( .A(n_330), .B(n_392), .Y(n_469) );
AOI32xp33_ASAP7_75t_L g542 ( .A1(n_330), .A2(n_543), .A3(n_545), .B1(n_546), .B2(n_547), .Y(n_542) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g383 ( .A(n_332), .Y(n_383) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g471 ( .A(n_336), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g391 ( .A(n_337), .B(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_337), .Y(n_524) );
AND2x2_ASAP7_75t_L g547 ( .A(n_337), .B(n_343), .Y(n_547) );
AO21x1_ASAP7_75t_L g513 ( .A1(n_338), .A2(n_514), .B(n_518), .Y(n_513) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_351), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_349), .Y(n_342) );
INVx1_ASAP7_75t_L g545 ( .A(n_343), .Y(n_545) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g368 ( .A(n_344), .Y(n_368) );
BUFx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_349), .B(n_412), .Y(n_444) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_349), .Y(n_506) );
INVx1_ASAP7_75t_L g415 ( .A(n_350), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_350), .B(n_460), .Y(n_532) );
NOR2xp67_ASAP7_75t_L g535 ( .A(n_350), .B(n_459), .Y(n_535) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g359 ( .A(n_352), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
OR2x2_ASAP7_75t_L g482 ( .A(n_353), .B(n_385), .Y(n_482) );
OA21x2_ASAP7_75t_L g658 ( .A1(n_355), .A2(n_659), .B(n_666), .Y(n_658) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OAI21xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B(n_361), .Y(n_357) );
INVx2_ASAP7_75t_L g509 ( .A(n_359), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_360), .B(n_395), .Y(n_446) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_363), .A2(n_488), .B(n_549), .C(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2x1p5_ASAP7_75t_L g428 ( .A(n_364), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g479 ( .A(n_364), .B(n_480), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_364), .B(n_395), .C(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g380 ( .A(n_366), .Y(n_380) );
INVx3_ASAP7_75t_L g478 ( .A(n_366), .Y(n_478) );
OR2x6_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_368), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_386), .Y(n_369) );
AOI22x1_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B1(n_380), .B2(n_381), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g475 ( .A(n_372), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_372), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g540 ( .A(n_373), .Y(n_540) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g453 ( .A(n_374), .Y(n_453) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g499 ( .A(n_379), .B(n_460), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_380), .A2(n_387), .B1(n_391), .B2(n_393), .Y(n_386) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_382), .B(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g403 ( .A(n_384), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_384), .B(n_423), .Y(n_492) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_384), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g546 ( .A(n_384), .B(n_442), .Y(n_546) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
OR2x2_ASAP7_75t_L g501 ( .A(n_389), .B(n_423), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_392), .B(n_412), .Y(n_447) );
INVx2_ASAP7_75t_L g488 ( .A(n_392), .Y(n_488) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
OR2x2_ASAP7_75t_L g433 ( .A(n_395), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_395), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g463 ( .A(n_395), .Y(n_463) );
BUFx3_ASAP7_75t_L g489 ( .A(n_396), .Y(n_489) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
BUFx2_ASAP7_75t_L g404 ( .A(n_398), .Y(n_404) );
INVx1_ASAP7_75t_L g423 ( .A(n_398), .Y(n_423) );
AND4x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_418), .C(n_436), .D(n_449), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI31xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .A3(n_409), .B(n_411), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g533 ( .A(n_410), .B(n_504), .Y(n_533) );
OR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_414), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g531 ( .A(n_417), .B(n_532), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_424), .B1(n_430), .B2(n_432), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
OR2x2_ASAP7_75t_L g519 ( .A(n_420), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_428), .A2(n_497), .B1(n_500), .B2(n_502), .C(n_505), .Y(n_496) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_434), .B(n_462), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_440), .B2(n_443), .C(n_445), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g448 ( .A(n_438), .Y(n_448) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx3_ASAP7_75t_R g490 ( .A(n_441), .Y(n_490) );
INVx2_ASAP7_75t_L g520 ( .A(n_442), .Y(n_520) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_454), .B1(n_457), .B2(n_461), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g518 ( .A1(n_452), .A2(n_519), .B(n_521), .C(n_523), .Y(n_518) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g544 ( .A(n_456), .Y(n_544) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g536 ( .A(n_463), .B(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_520), .Y(n_541) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_483), .Y(n_464) );
OAI21xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_474), .B(n_477), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g539 ( .A1(n_470), .A2(n_501), .B1(n_540), .B2(n_541), .C(n_542), .Y(n_539) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g487 ( .A(n_472), .Y(n_487) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_481), .Y(n_477) );
NAND2x1_ASAP7_75t_L g526 ( .A(n_478), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g497 ( .A(n_480), .B(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
AOI322xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_489), .A3(n_490), .B1(n_491), .B2(n_493), .C1(n_494), .C2(n_924), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_526), .B(n_529), .Y(n_525) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g516 ( .A(n_498), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_509), .B2(n_510), .Y(n_505) );
NOR4xp75_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .C(n_539), .D(n_548), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVxp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_533), .B1(n_534), .B2(n_536), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g550 ( .A(n_538), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
CKINVDCx11_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g907 ( .A(n_559), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_559), .B(n_912), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_902), .B(n_908), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_566), .B2(n_901), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_SL g901 ( .A(n_566), .Y(n_901) );
INVx11_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx8_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_816), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_725), .C(n_775), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_697), .Y(n_573) );
OAI21xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_642), .B(n_667), .Y(n_574) );
NAND2x1_ASAP7_75t_SL g575 ( .A(n_576), .B(n_590), .Y(n_575) );
INVx1_ASAP7_75t_L g706 ( .A(n_576), .Y(n_706) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_SL g694 ( .A(n_577), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_577), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g774 ( .A(n_577), .B(n_728), .Y(n_774) );
INVx2_ASAP7_75t_L g859 ( .A(n_577), .Y(n_859) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g756 ( .A(n_578), .Y(n_756) );
INVx1_ASAP7_75t_L g810 ( .A(n_578), .Y(n_810) );
AND2x2_ASAP7_75t_L g885 ( .A(n_578), .B(n_628), .Y(n_885) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g714 ( .A(n_579), .B(n_628), .Y(n_714) );
INVxp33_ASAP7_75t_L g761 ( .A(n_579), .Y(n_761) );
INVx2_ASAP7_75t_SL g636 ( .A(n_584), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_585), .A2(n_650), .B(n_651), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_585), .A2(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g796 ( .A(n_590), .Y(n_796) );
OAI21xp33_ASAP7_75t_L g856 ( .A1(n_590), .A2(n_780), .B(n_857), .Y(n_856) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_611), .Y(n_590) );
OR2x2_ASAP7_75t_L g727 ( .A(n_591), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g716 ( .A(n_593), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g723 ( .A(n_593), .B(n_612), .Y(n_723) );
AND2x2_ASAP7_75t_L g760 ( .A(n_593), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g795 ( .A(n_593), .B(n_717), .Y(n_795) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_594), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g778 ( .A(n_594), .B(n_756), .Y(n_778) );
AO21x2_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_602), .Y(n_594) );
AO21x1_ASAP7_75t_SL g710 ( .A1(n_595), .A2(n_597), .B(n_602), .Y(n_710) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OAI21x1_ASAP7_75t_SL g602 ( .A1(n_596), .A2(n_603), .B(n_610), .Y(n_602) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B(n_609), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g614 ( .A(n_606), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_609), .A2(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g808 ( .A(n_611), .B(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g890 ( .A(n_611), .B(n_709), .Y(n_890) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_627), .Y(n_611) );
OR2x2_ASAP7_75t_L g696 ( .A(n_612), .B(n_628), .Y(n_696) );
INVx2_ASAP7_75t_L g717 ( .A(n_612), .Y(n_717) );
INVx1_ASAP7_75t_L g730 ( .A(n_612), .Y(n_730) );
INVx1_ASAP7_75t_L g746 ( .A(n_612), .Y(n_746) );
AND2x2_ASAP7_75t_L g843 ( .A(n_612), .B(n_729), .Y(n_843) );
AO21x2_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_618), .B(n_624), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g615 ( .A(n_614), .B(n_616), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_623), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_623), .A2(n_625), .B(n_626), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_625), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g630 ( .A(n_626), .B(n_631), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_626), .A2(n_660), .B(n_663), .Y(n_659) );
INVx2_ASAP7_75t_L g729 ( .A(n_627), .Y(n_729) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g788 ( .A(n_628), .Y(n_788) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_629), .B(n_637), .Y(n_628) );
NAND2x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AOI21x1_ASAP7_75t_L g637 ( .A1(n_630), .A2(n_638), .B(n_641), .Y(n_637) );
O2A1O1Ixp5_ASAP7_75t_L g648 ( .A1(n_630), .A2(n_649), .B(n_652), .C(n_655), .Y(n_648) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x6_ASAP7_75t_L g803 ( .A(n_644), .B(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_L g878 ( .A(n_644), .B(n_879), .Y(n_878) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_657), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_645), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g719 ( .A(n_645), .Y(n_719) );
AND2x2_ASAP7_75t_L g779 ( .A(n_645), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_646), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g769 ( .A(n_646), .B(n_687), .Y(n_769) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_SL g703 ( .A(n_647), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_647), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_647), .B(n_658), .Y(n_739) );
INVx1_ASAP7_75t_L g748 ( .A(n_647), .Y(n_748) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g854 ( .A(n_657), .B(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g670 ( .A(n_658), .Y(n_670) );
INVx1_ASAP7_75t_L g705 ( .A(n_658), .Y(n_705) );
INVx1_ASAP7_75t_L g737 ( .A(n_658), .Y(n_737) );
AND2x2_ASAP7_75t_L g752 ( .A(n_658), .B(n_674), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_658), .B(n_674), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_686), .B(n_694), .Y(n_667) );
AND2x4_ASAP7_75t_L g828 ( .A(n_668), .B(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_668), .B(n_829), .Y(n_870) );
AND2x4_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g827 ( .A(n_669), .Y(n_827) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_670), .B(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g762 ( .A(n_672), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g701 ( .A(n_673), .Y(n_701) );
AND2x2_ASAP7_75t_L g721 ( .A(n_673), .B(n_687), .Y(n_721) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_674), .Y(n_734) );
OR2x2_ASAP7_75t_L g741 ( .A(n_674), .B(n_687), .Y(n_741) );
AND2x2_ASAP7_75t_L g771 ( .A(n_674), .B(n_705), .Y(n_771) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B(n_685), .Y(n_678) );
AND2x4_ASAP7_75t_L g770 ( .A(n_686), .B(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_L g704 ( .A(n_687), .B(n_705), .Y(n_704) );
BUFx3_ASAP7_75t_L g754 ( .A(n_687), .Y(n_754) );
INVx2_ASAP7_75t_SL g764 ( .A(n_687), .Y(n_764) );
AND2x2_ASAP7_75t_L g892 ( .A(n_687), .B(n_701), .Y(n_892) );
AO31x2_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .A3(n_691), .B(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g759 ( .A(n_696), .Y(n_759) );
OR2x2_ASAP7_75t_L g815 ( .A(n_696), .B(n_810), .Y(n_815) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_706), .A3(n_707), .B1(n_711), .B2(n_718), .C1(n_722), .C2(n_724), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g866 ( .A(n_700), .B(n_739), .Y(n_866) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g805 ( .A(n_701), .B(n_764), .Y(n_805) );
INVx1_ASAP7_75t_L g855 ( .A(n_701), .Y(n_855) );
NOR2x1_ASAP7_75t_SL g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g751 ( .A(n_703), .B(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g847 ( .A(n_703), .B(n_704), .Y(n_847) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_704), .Y(n_724) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g849 ( .A(n_708), .B(n_850), .Y(n_849) );
AND2x4_ASAP7_75t_L g862 ( .A(n_708), .B(n_863), .Y(n_862) );
AND2x2_ASAP7_75t_L g865 ( .A(n_708), .B(n_759), .Y(n_865) );
NAND2x1_ASAP7_75t_L g869 ( .A(n_708), .B(n_712), .Y(n_869) );
INVx5_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g753 ( .A(n_709), .B(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_L g802 ( .A(n_709), .B(n_799), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_709), .B(n_820), .Y(n_819) );
AND2x4_ASAP7_75t_L g842 ( .A(n_709), .B(n_843), .Y(n_842) );
AND2x2_ASAP7_75t_L g880 ( .A(n_709), .B(n_712), .Y(n_880) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g786 ( .A(n_710), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
NAND2x1_ASAP7_75t_L g837 ( .A(n_712), .B(n_823), .Y(n_837) );
INVx6_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx4_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_714), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g882 ( .A(n_716), .B(n_883), .Y(n_882) );
OR2x2_ASAP7_75t_L g899 ( .A(n_716), .B(n_755), .Y(n_899) );
OR2x2_ASAP7_75t_L g799 ( .A(n_717), .B(n_756), .Y(n_799) );
INVx1_ASAP7_75t_L g823 ( .A(n_717), .Y(n_823) );
AND2x2_ASAP7_75t_L g863 ( .A(n_717), .B(n_761), .Y(n_863) );
OR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
AND2x2_ASAP7_75t_L g891 ( .A(n_719), .B(n_892), .Y(n_891) );
A2O1A1Ixp33_ASAP7_75t_L g818 ( .A1(n_720), .A2(n_819), .B(n_821), .C(n_824), .Y(n_818) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g773 ( .A(n_721), .B(n_739), .Y(n_773) );
AND2x2_ASAP7_75t_L g800 ( .A(n_721), .B(n_735), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_723), .B(n_885), .Y(n_884) );
AOI211xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_731), .B(n_742), .C(n_765), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g840 ( .A(n_728), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
OR2x2_ASAP7_75t_L g755 ( .A(n_729), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g833 ( .A(n_730), .B(n_756), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_738), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g749 ( .A(n_734), .Y(n_749) );
AND2x2_ASAP7_75t_L g876 ( .A(n_735), .B(n_764), .Y(n_876) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g791 ( .A(n_736), .B(n_741), .Y(n_791) );
BUFx2_ASAP7_75t_L g888 ( .A(n_736), .Y(n_888) );
OAI221xp5_ASAP7_75t_SL g881 ( .A1(n_738), .A2(n_882), .B1(n_884), .B2(n_886), .C(n_889), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_SL g898 ( .A(n_739), .Y(n_898) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI322xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_747), .A3(n_749), .B1(n_750), .B2(n_755), .C1(n_757), .C2(n_762), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g826 ( .A(n_745), .Y(n_826) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_751), .B(n_783), .Y(n_782) );
OAI21xp33_ASAP7_75t_L g811 ( .A1(n_751), .A2(n_812), .B(n_814), .Y(n_811) );
INVx2_ASAP7_75t_L g838 ( .A(n_751), .Y(n_838) );
AND2x4_ASAP7_75t_SL g780 ( .A(n_752), .B(n_764), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_752), .B(n_754), .Y(n_813) );
BUFx2_ASAP7_75t_L g896 ( .A(n_752), .Y(n_896) );
INVx1_ASAP7_75t_L g784 ( .A(n_754), .Y(n_784) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_754), .Y(n_829) );
INVx1_ASAP7_75t_L g852 ( .A(n_754), .Y(n_852) );
AOI32xp33_ASAP7_75t_L g889 ( .A1(n_754), .A2(n_842), .A3(n_887), .B1(n_890), .B2(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g793 ( .A(n_755), .Y(n_793) );
INVx1_ASAP7_75t_L g850 ( .A(n_755), .Y(n_850) );
INVx2_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_L g835 ( .A(n_759), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_760), .B(n_840), .Y(n_846) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_772), .B(n_774), .Y(n_765) );
NOR2x1_ASAP7_75t_R g766 ( .A(n_767), .B(n_770), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AND2x2_ASAP7_75t_L g895 ( .A(n_769), .B(n_896), .Y(n_895) );
INVx3_ASAP7_75t_L g806 ( .A(n_770), .Y(n_806) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI211xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_779), .B(n_781), .C(n_801), .Y(n_775) );
INVxp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g822 ( .A(n_778), .B(n_823), .Y(n_822) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_779), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_785), .B(n_789), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g897 ( .A(n_784), .B(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_784), .B(n_854), .Y(n_900) );
NAND2x1p5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
INVx1_ASAP7_75t_L g798 ( .A(n_787), .Y(n_798) );
INVx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_792), .B1(n_797), .B2(n_800), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OAI21xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B(n_796), .Y(n_792) );
OAI222xp33_ASAP7_75t_L g893 ( .A1(n_794), .A2(n_802), .B1(n_894), .B2(n_897), .C1(n_899), .C2(n_900), .Y(n_893) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_798), .Y(n_820) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B1(n_806), .B2(n_807), .C(n_811), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_803), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_836) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_805), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g825 ( .A(n_809), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g883 ( .A(n_809), .Y(n_883) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_841), .C(n_867), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_827), .B1(n_828), .B2(n_830), .C(n_836), .Y(n_817) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g858 ( .A(n_823), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_834), .Y(n_830) );
INVxp67_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
BUFx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI21xp33_ASAP7_75t_L g860 ( .A1(n_838), .A2(n_861), .B(n_864), .Y(n_860) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI211xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .B(n_845), .C(n_860), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_843), .B(n_859), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B1(n_848), .B2(n_851), .C(n_856), .Y(n_845) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
OR2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
INVxp67_ASAP7_75t_L g879 ( .A(n_852), .Y(n_879) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NOR2xp33_ASAP7_75t_SL g857 ( .A(n_858), .B(n_859), .Y(n_857) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
NOR3xp33_ASAP7_75t_L g867 ( .A(n_868), .B(n_881), .C(n_893), .Y(n_867) );
OAI21xp33_ASAP7_75t_SL g868 ( .A1(n_869), .A2(n_870), .B(n_871), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_874), .B1(n_877), .B2(n_880), .Y(n_871) );
INVx2_ASAP7_75t_SL g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx6_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
OR2x6_ASAP7_75t_L g903 ( .A(n_904), .B(n_907), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_905), .Y(n_916) );
INVx2_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
BUFx3_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
BUFx10_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
BUFx6f_ASAP7_75t_SL g914 ( .A(n_915), .Y(n_914) );
BUFx3_ASAP7_75t_L g922 ( .A(n_915), .Y(n_922) );
AND2x4_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
endmodule