module fake_jpeg_28463_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

AND2x4_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_18),
.Y(n_22)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_16),
.B1(n_13),
.B2(n_9),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B1(n_27),
.B2(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_21),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_31),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_32),
.C(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_12),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_25),
.B1(n_13),
.B2(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.C(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_45),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_41),
.B(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_46),
.C(n_5),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B(n_47),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_5),
.C(n_6),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_6),
.Y(n_53)
);

AOI321xp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_7),
.C(n_35),
.Y(n_54)
);

BUFx24_ASAP7_75t_SL g55 ( 
.A(n_54),
.Y(n_55)
);


endmodule