module fake_jpeg_25642_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_12),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_26),
.B1(n_13),
.B2(n_15),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_22),
.B1(n_23),
.B2(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_26),
.B1(n_15),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_47),
.B1(n_18),
.B2(n_22),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_26),
.B1(n_35),
.B2(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_59),
.B1(n_42),
.B2(n_48),
.Y(n_82)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_48),
.B1(n_44),
.B2(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_63),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_36),
.B(n_28),
.C(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_29),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_48),
.B1(n_40),
.B2(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_70),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_53),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_82),
.B(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_40),
.B1(n_58),
.B2(n_39),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_44),
.B1(n_70),
.B2(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_89),
.Y(n_105)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_69),
.B1(n_64),
.B2(n_52),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_63),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_95),
.C(n_89),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_94),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_58),
.C(n_60),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_88),
.B1(n_75),
.B2(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_40),
.B1(n_68),
.B2(n_61),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_75),
.B1(n_87),
.B2(n_84),
.Y(n_126)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_103),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_109),
.B(n_76),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_59),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_85),
.B1(n_74),
.B2(n_80),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_78),
.B1(n_82),
.B2(n_73),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_130),
.B(n_105),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_18),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_124),
.B1(n_127),
.B2(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_126),
.B1(n_128),
.B2(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_65),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_73),
.B1(n_72),
.B2(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_73),
.B1(n_72),
.B2(n_47),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_55),
.B1(n_62),
.B2(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_99),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_71),
.B(n_18),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_62),
.B1(n_71),
.B2(n_51),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_104),
.B1(n_100),
.B2(n_97),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_148),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_138),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_139),
.B(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_143),
.B1(n_149),
.B2(n_151),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_95),
.B1(n_104),
.B2(n_102),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_129),
.C(n_114),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_117),
.B1(n_127),
.B2(n_128),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_130),
.B(n_132),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_118),
.B(n_124),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_103),
.B1(n_99),
.B2(n_62),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_33),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_127),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_115),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_169),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_131),
.B1(n_132),
.B2(n_116),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_167),
.B(n_175),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_121),
.C(n_131),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_125),
.B1(n_106),
.B2(n_14),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_19),
.B1(n_16),
.B2(n_14),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_106),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_179),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_137),
.B(n_140),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_137),
.B1(n_155),
.B2(n_106),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_27),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_27),
.B1(n_25),
.B2(n_33),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_140),
.B(n_135),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_147),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.C(n_151),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_33),
.C(n_32),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

BUFx12_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_197),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_160),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_142),
.C(n_154),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_193),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_165),
.B1(n_170),
.B2(n_175),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_196),
.B(n_199),
.Y(n_208)
);

XOR2x1_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_25),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_16),
.B1(n_19),
.B2(n_14),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_19),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_201),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_159),
.B(n_173),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_210),
.B(n_158),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_209),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_162),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_159),
.B(n_173),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_166),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_195),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_188),
.B1(n_200),
.B2(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_221),
.B1(n_234),
.B2(n_203),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_161),
.B1(n_190),
.B2(n_189),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_187),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_185),
.C(n_182),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_228),
.C(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_182),
.C(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_218),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_232),
.B(n_204),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_9),
.B(n_12),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_7),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_236),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_210),
.C(n_208),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_245),
.C(n_246),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_224),
.A2(n_32),
.B(n_19),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_241),
.A2(n_234),
.B(n_219),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_220),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_16),
.B1(n_17),
.B2(n_32),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_247),
.B1(n_6),
.B2(n_12),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_230),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_27),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_17),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_248),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_226),
.B1(n_222),
.B2(n_8),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_4),
.B1(n_11),
.B2(n_10),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_255),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_17),
.B(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_258),
.C(n_4),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_5),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_0),
.C(n_1),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_238),
.C(n_239),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_5),
.B(n_11),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_262),
.Y(n_272)
);

OAI321xp33_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_246),
.A3(n_239),
.B1(n_8),
.B2(n_3),
.C(n_4),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_267),
.B(n_3),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_251),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_4),
.B1(n_11),
.B2(n_10),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_265),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_3),
.C(n_10),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_268),
.B(n_269),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_256),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_259),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_276),
.B(n_273),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_272),
.C(n_266),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_278),
.B(n_267),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_12),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_0),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_282),
.A2(n_0),
.B(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_0),
.C(n_2),
.Y(n_284)
);


endmodule