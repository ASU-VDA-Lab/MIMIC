module fake_jpeg_16644_n_113 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_61),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_49),
.B1(n_55),
.B2(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_74),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_54),
.B1(n_57),
.B2(n_50),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_70),
.B1(n_77),
.B2(n_80),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_52),
.B1(n_48),
.B2(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_53),
.B1(n_56),
.B2(n_3),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_19),
.B1(n_39),
.B2(n_37),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_78),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_1),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_51),
.B(n_2),
.C(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_15),
.B1(n_36),
.B2(n_33),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_87),
.B(n_69),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_88),
.B1(n_73),
.B2(n_71),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_75),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_79),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_93),
.B(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_101),
.B1(n_82),
.B2(n_97),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_87),
.B1(n_98),
.B2(n_71),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_20),
.B(n_32),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_16),
.B1(n_27),
.B2(n_6),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_14),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_22),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_12),
.B(n_29),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_80),
.C(n_11),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_9),
.B(n_10),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_112),
.Y(n_113)
);


endmodule