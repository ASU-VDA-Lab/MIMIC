module fake_jpeg_13536_n_389 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_55),
.Y(n_117)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_13),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_0),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_81),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_78),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_10),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_2),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_22),
.B1(n_17),
.B2(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_86),
.A2(n_107),
.B1(n_115),
.B2(n_3),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_17),
.B(n_34),
.Y(n_87)
);

OR2x2_ASAP7_75t_SL g153 ( 
.A(n_87),
.B(n_127),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_22),
.B1(n_26),
.B2(n_15),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_48),
.A2(n_15),
.B1(n_26),
.B2(n_31),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_10),
.C(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_26),
.B1(n_37),
.B2(n_31),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_40),
.B1(n_37),
.B2(n_31),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_124),
.B1(n_40),
.B2(n_66),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_46),
.B(n_39),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_39),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_121),
.B(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_77),
.B(n_29),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_32),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_50),
.A2(n_40),
.B1(n_37),
.B2(n_33),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_29),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_20),
.C(n_24),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_132),
.B(n_134),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_21),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_21),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_139),
.B(n_140),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_33),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_99),
.C(n_96),
.Y(n_141)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_153),
.B(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_52),
.B1(n_58),
.B2(n_67),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_150),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_62),
.B1(n_60),
.B2(n_69),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_146),
.B(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_127),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_81),
.B1(n_80),
.B2(n_71),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_102),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_72),
.B1(n_56),
.B2(n_53),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_85),
.B1(n_120),
.B2(n_142),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_91),
.B(n_32),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_104),
.B(n_45),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_164),
.B(n_84),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_2),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_88),
.B(n_3),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_85),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_171),
.B1(n_175),
.B2(n_120),
.Y(n_210)
);

AO22x2_ASAP7_75t_L g167 ( 
.A1(n_98),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_131),
.B1(n_98),
.B2(n_103),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_84),
.B1(n_131),
.B2(n_97),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_93),
.A2(n_8),
.B1(n_10),
.B2(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_101),
.A2(n_129),
.B1(n_130),
.B2(n_97),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_126),
.C(n_108),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_108),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_171),
.B1(n_166),
.B2(n_148),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_150),
.B1(n_137),
.B2(n_167),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_138),
.A2(n_170),
.B(n_174),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_157),
.B(n_159),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_144),
.C(n_133),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_158),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_235),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_219),
.A2(n_222),
.B1(n_231),
.B2(n_220),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_187),
.B1(n_199),
.B2(n_207),
.Y(n_222)
);

AO21x2_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_167),
.B(n_143),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_224),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_176),
.B(n_135),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_248),
.B(n_193),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_233),
.C(n_236),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_180),
.B(n_191),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_140),
.B1(n_164),
.B2(n_163),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_151),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_167),
.B(n_147),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_167),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_238),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_172),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_246),
.Y(n_265)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_152),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_249),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_247),
.B1(n_195),
.B2(n_180),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_137),
.B1(n_191),
.B2(n_206),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_206),
.B(n_191),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_186),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_254),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_213),
.B(n_197),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_271),
.B(n_278),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_218),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_264),
.B1(n_268),
.B2(n_273),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_195),
.B1(n_177),
.B2(n_196),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_267),
.B1(n_243),
.B2(n_208),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_222),
.A2(n_178),
.B1(n_179),
.B2(n_196),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_245),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_186),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_232),
.A2(n_182),
.B(n_183),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_275),
.B(n_224),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_224),
.A2(n_244),
.B1(n_221),
.B2(n_218),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_232),
.A2(n_183),
.B(n_212),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_220),
.A2(n_188),
.B(n_184),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_240),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_220),
.B1(n_219),
.B2(n_231),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_294),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_234),
.B1(n_224),
.B2(n_221),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_217),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_224),
.B1(n_225),
.B2(n_230),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_226),
.B(n_238),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_252),
.B(n_226),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_299),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_224),
.B1(n_229),
.B2(n_243),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_229),
.C(n_208),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_300),
.C(n_278),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_297),
.A2(n_302),
.B(n_265),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_268),
.B1(n_270),
.B2(n_274),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_253),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_228),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_SL g302 ( 
.A(n_253),
.B(n_242),
.C(n_228),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_266),
.B1(n_276),
.B2(n_271),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_284),
.B1(n_294),
.B2(n_282),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_306),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_312),
.B1(n_322),
.B2(n_269),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_251),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_277),
.C(n_251),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_280),
.C(n_295),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_264),
.B1(n_258),
.B2(n_271),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_289),
.A2(n_267),
.B1(n_250),
.B2(n_257),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_284),
.B1(n_301),
.B2(n_283),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_279),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_319),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_300),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_198),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_318),
.A2(n_302),
.B1(n_272),
.B2(n_282),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_297),
.A2(n_265),
.B(n_275),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_290),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_321),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_286),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_260),
.B1(n_256),
.B2(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_312),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_306),
.B(n_291),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_339),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_326),
.A2(n_328),
.B1(n_313),
.B2(n_315),
.Y(n_351)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_301),
.C(n_285),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_285),
.C(n_256),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_269),
.C(n_228),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_340),
.Y(n_350)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_321),
.B1(n_320),
.B2(n_308),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

BUFx12_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_345),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_329),
.B(n_310),
.Y(n_347)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_347),
.Y(n_359)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_352),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_316),
.Y(n_352)
);

INVx13_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_320),
.B1(n_308),
.B2(n_305),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_342),
.C(n_329),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_355),
.B(n_362),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_335),
.C(n_334),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_332),
.C(n_325),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_311),
.C(n_348),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_341),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_367),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g365 ( 
.A1(n_356),
.A2(n_327),
.B(n_311),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_365),
.A2(n_361),
.B(n_352),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_351),
.B(n_326),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_366),
.B(n_368),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_337),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_349),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_372),
.C(n_354),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_352),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_376),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_361),
.B1(n_344),
.B2(n_349),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_378),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_369),
.A2(n_331),
.B1(n_303),
.B2(n_318),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_373),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_380),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_373),
.A2(n_370),
.B(n_374),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_382),
.B(n_350),
.Y(n_384)
);

OAI311xp33_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_381),
.A3(n_353),
.B1(n_372),
.C1(n_366),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_383),
.C(n_319),
.Y(n_386)
);

OAI21x1_ASAP7_75t_SL g387 ( 
.A1(n_386),
.A2(n_345),
.B(n_204),
.Y(n_387)
);

OAI211xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_198),
.B(n_345),
.C(n_379),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_388),
.Y(n_389)
);


endmodule