module real_aes_7610_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
INVx1_ASAP7_75t_L g495 ( .A(n_1), .Y(n_495) );
INVx1_ASAP7_75t_L g274 ( .A(n_2), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_3), .A2(n_36), .B1(n_193), .B2(n_523), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g181 ( .A1(n_4), .A2(n_182), .B(n_183), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_5), .B(n_180), .Y(n_472) );
AND2x6_ASAP7_75t_L g155 ( .A(n_6), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_7), .A2(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_8), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_8), .B(n_37), .Y(n_128) );
INVx1_ASAP7_75t_L g190 ( .A(n_9), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_10), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g152 ( .A(n_11), .Y(n_152) );
INVx1_ASAP7_75t_L g491 ( .A(n_12), .Y(n_491) );
INVx1_ASAP7_75t_L g256 ( .A(n_13), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_14), .B(n_158), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_15), .B(n_148), .Y(n_500) );
AO32x2_ASAP7_75t_L g520 ( .A1(n_16), .A2(n_147), .A3(n_180), .B1(n_483), .B2(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_17), .B(n_193), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_18), .B(n_201), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_19), .B(n_148), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_20), .A2(n_49), .B1(n_193), .B2(n_523), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_21), .B(n_182), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_22), .A2(n_75), .B1(n_158), .B2(n_193), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_23), .B(n_193), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_24), .B(n_178), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_25), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_26), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_27), .B(n_195), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_28), .B(n_188), .Y(n_275) );
INVx1_ASAP7_75t_L g166 ( .A(n_29), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_30), .B(n_195), .Y(n_517) );
INVx2_ASAP7_75t_L g160 ( .A(n_31), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_32), .B(n_193), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_33), .B(n_195), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_34), .A2(n_41), .B1(n_751), .B2(n_752), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_34), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_35), .A2(n_155), .B(n_167), .C(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g109 ( .A(n_37), .Y(n_109) );
INVx1_ASAP7_75t_L g164 ( .A(n_38), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_39), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_40), .B(n_188), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_41), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_42), .B(n_193), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_43), .A2(n_87), .B1(n_218), .B2(n_523), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_44), .B(n_193), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_45), .B(n_193), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_46), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_47), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_48), .B(n_182), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_50), .A2(n_59), .B1(n_158), .B2(n_193), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_51), .A2(n_158), .B1(n_161), .B2(n_167), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_52), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_53), .B(n_193), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_54), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_55), .B(n_193), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_56), .A2(n_187), .B(n_189), .C(n_192), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_57), .Y(n_231) );
INVx1_ASAP7_75t_L g184 ( .A(n_58), .Y(n_184) );
INVx1_ASAP7_75t_L g156 ( .A(n_60), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_61), .B(n_193), .Y(n_496) );
INVx1_ASAP7_75t_L g151 ( .A(n_62), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_63), .Y(n_121) );
AO32x2_ASAP7_75t_L g540 ( .A1(n_64), .A2(n_180), .A3(n_236), .B1(n_483), .B2(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g480 ( .A(n_65), .Y(n_480) );
INVx1_ASAP7_75t_L g512 ( .A(n_66), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_67), .A2(n_749), .B1(n_750), .B2(n_753), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_67), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_SL g200 ( .A1(n_68), .A2(n_192), .B(n_201), .C(n_202), .Y(n_200) );
INVxp67_ASAP7_75t_L g203 ( .A(n_69), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_70), .B(n_158), .Y(n_513) );
INVx1_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_72), .Y(n_175) );
INVx1_ASAP7_75t_L g224 ( .A(n_73), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_74), .A2(n_101), .B1(n_136), .B2(n_137), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_74), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_76), .A2(n_104), .B1(n_115), .B2(n_755), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_77), .A2(n_155), .B(n_167), .C(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_78), .B(n_523), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_79), .B(n_158), .Y(n_516) );
AOI222xp33_ASAP7_75t_SL g130 ( .A1(n_80), .A2(n_131), .B1(n_132), .B2(n_138), .C1(n_738), .C2(n_741), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_81), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_83), .B(n_201), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_84), .B(n_158), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_85), .A2(n_155), .B(n_167), .C(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
OR2x2_ASAP7_75t_L g124 ( .A(n_86), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g454 ( .A(n_86), .B(n_126), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_88), .A2(n_102), .B1(n_158), .B2(n_159), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_89), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_90), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_91), .A2(n_155), .B(n_167), .C(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_92), .Y(n_246) );
INVx1_ASAP7_75t_L g199 ( .A(n_93), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_94), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_95), .B(n_214), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_96), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_96), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_97), .B(n_158), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_98), .B(n_180), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_100), .A2(n_182), .B(n_198), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g137 ( .A(n_101), .Y(n_137) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g756 ( .A(n_107), .Y(n_756) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x2_ASAP7_75t_L g737 ( .A(n_111), .B(n_126), .Y(n_737) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_111), .B(n_125), .Y(n_743) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_130), .B1(n_744), .B2(n_745), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g744 ( .A(n_119), .Y(n_744) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_122), .A2(n_746), .B(n_754), .Y(n_745) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_129), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_124), .Y(n_754) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
CKINVDCx14_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_452), .B1(n_455), .B2(n_735), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_139), .A2(n_140), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_140), .A2(n_452), .B1(n_739), .B2(n_740), .Y(n_738) );
AND3x1_ASAP7_75t_L g140 ( .A(n_141), .B(n_377), .C(n_426), .Y(n_140) );
NOR3xp33_ASAP7_75t_SL g141 ( .A(n_142), .B(n_284), .C(n_322), .Y(n_141) );
OAI222xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_205), .B1(n_259), .B2(n_265), .C1(n_279), .C2(n_282), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_176), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_144), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_144), .B(n_327), .Y(n_418) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g295 ( .A(n_145), .B(n_196), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_145), .B(n_177), .Y(n_303) );
AND2x2_ASAP7_75t_L g338 ( .A(n_145), .B(n_315), .Y(n_338) );
OR2x2_ASAP7_75t_L g362 ( .A(n_145), .B(n_177), .Y(n_362) );
OR2x2_ASAP7_75t_L g370 ( .A(n_145), .B(n_269), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_145), .B(n_196), .Y(n_373) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g267 ( .A(n_146), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_146), .B(n_196), .Y(n_281) );
AND2x2_ASAP7_75t_L g331 ( .A(n_146), .B(n_269), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_146), .B(n_177), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_146), .B(n_430), .Y(n_451) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B(n_174), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_147), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g219 ( .A(n_147), .Y(n_219) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_147), .A2(n_270), .B(n_277), .Y(n_269) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_149), .B(n_150), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_157), .B1(n_170), .B2(n_171), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_154), .A2(n_184), .B(n_185), .C(n_186), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_185), .B(n_199), .C(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_154), .A2(n_185), .B(n_252), .C(n_253), .Y(n_251) );
INVx4_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_155), .B(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g182 ( .A(n_155), .B(n_172), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_155), .A2(n_464), .B(n_467), .Y(n_463) );
BUFx3_ASAP7_75t_L g483 ( .A(n_155), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_155), .A2(n_490), .B(n_494), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_155), .A2(n_511), .B(n_514), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_155), .A2(n_527), .B(n_531), .Y(n_526) );
INVx2_ASAP7_75t_L g276 ( .A(n_158), .Y(n_276) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
INVx1_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g161 ( .A1(n_162), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_161) );
INVx2_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
INVx4_ASAP7_75t_L g254 ( .A(n_162), .Y(n_254) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
AND2x2_ASAP7_75t_L g172 ( .A(n_163), .B(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
INVx3_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
INVx1_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
INVx5_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
AND2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_168), .Y(n_193) );
BUFx3_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVx1_ASAP7_75t_L g523 ( .A(n_168), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_171), .A2(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_171), .A2(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g470 ( .A(n_173), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_176), .A2(n_370), .B(n_371), .C(n_374), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_176), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_176), .B(n_314), .Y(n_436) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_196), .Y(n_176) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_177), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_177), .B(n_315), .Y(n_321) );
INVx1_ASAP7_75t_SL g329 ( .A(n_177), .Y(n_329) );
AND2x2_ASAP7_75t_L g352 ( .A(n_177), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g430 ( .A(n_177), .Y(n_430) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_181), .B(n_194), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_SL g220 ( .A(n_179), .B(n_221), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_179), .B(n_483), .C(n_502), .Y(n_501) );
AO21x1_ASAP7_75t_L g546 ( .A1(n_179), .A2(n_502), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_180), .A2(n_197), .B(n_204), .Y(n_196) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_180), .A2(n_463), .B(n_472), .Y(n_462) );
BUFx2_ASAP7_75t_L g250 ( .A(n_182), .Y(n_250) );
O2A1O1Ixp5_ASAP7_75t_L g479 ( .A1(n_187), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_187), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx4_ASAP7_75t_L g242 ( .A(n_188), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_188), .A2(n_471), .B1(n_503), .B2(n_504), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_188), .A2(n_471), .B1(n_522), .B2(n_524), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g541 ( .A1(n_188), .A2(n_191), .B1(n_542), .B2(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_191), .B(n_203), .Y(n_202) );
INVx5_ASAP7_75t_L g214 ( .A(n_191), .Y(n_214) );
O2A1O1Ixp5_ASAP7_75t_SL g511 ( .A1(n_192), .A2(n_214), .B(n_512), .C(n_513), .Y(n_511) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_193), .Y(n_243) );
INVx1_ASAP7_75t_L g232 ( .A(n_195), .Y(n_232) );
INVx2_ASAP7_75t_L g236 ( .A(n_195), .Y(n_236) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_195), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_195), .A2(n_510), .B(n_517), .Y(n_509) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_195), .A2(n_526), .B(n_534), .Y(n_525) );
BUFx2_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
INVx1_ASAP7_75t_L g328 ( .A(n_196), .Y(n_328) );
INVx3_ASAP7_75t_L g353 ( .A(n_196), .Y(n_353) );
INVx1_ASAP7_75t_L g530 ( .A(n_201), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_205), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_233), .Y(n_205) );
INVx1_ASAP7_75t_L g349 ( .A(n_206), .Y(n_349) );
OAI32xp33_ASAP7_75t_L g355 ( .A1(n_206), .A2(n_294), .A3(n_356), .B1(n_357), .B2(n_358), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_206), .A2(n_360), .B1(n_363), .B2(n_368), .Y(n_359) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g297 ( .A(n_207), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g375 ( .A(n_207), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g445 ( .A(n_207), .B(n_391), .Y(n_445) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g260 ( .A(n_208), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
INVx1_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
OR2x2_ASAP7_75t_L g317 ( .A(n_208), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g324 ( .A(n_208), .B(n_298), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_208), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_208), .B(n_263), .Y(n_345) );
INVx3_ASAP7_75t_L g367 ( .A(n_208), .Y(n_367) );
AND2x2_ASAP7_75t_L g392 ( .A(n_208), .B(n_264), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_208), .B(n_357), .Y(n_440) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_211), .B(n_219), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_215), .B(n_216), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_214), .A2(n_274), .B(n_275), .C(n_276), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_214), .A2(n_465), .B(n_466), .Y(n_464) );
INVx2_ASAP7_75t_L g471 ( .A(n_214), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_214), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
INVx1_ASAP7_75t_L g229 ( .A(n_219), .Y(n_229) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_219), .A2(n_475), .B(n_484), .Y(n_474) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_219), .A2(n_489), .B(n_497), .Y(n_488) );
INVx2_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
AND2x2_ASAP7_75t_L g396 ( .A(n_222), .B(n_234), .Y(n_396) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_230), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_232), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_232), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g438 ( .A(n_233), .Y(n_438) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_247), .Y(n_233) );
INVx1_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
AND2x2_ASAP7_75t_L g310 ( .A(n_234), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_234), .B(n_264), .Y(n_318) );
AND2x2_ASAP7_75t_L g376 ( .A(n_234), .B(n_299), .Y(n_376) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g262 ( .A(n_235), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_235), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g298 ( .A(n_235), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_235), .B(n_264), .Y(n_364) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_247), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_247), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_247), .B(n_264), .Y(n_357) );
AND2x2_ASAP7_75t_L g366 ( .A(n_247), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g391 ( .A(n_247), .Y(n_391) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g263 ( .A(n_248), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g299 ( .A(n_248), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g493 ( .A(n_254), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_254), .A2(n_515), .B(n_516), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_259), .A2(n_269), .B1(n_428), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OAI21xp5_ASAP7_75t_SL g450 ( .A1(n_261), .A2(n_372), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_262), .B(n_367), .Y(n_384) );
INVx1_ASAP7_75t_L g409 ( .A(n_262), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_263), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g336 ( .A(n_263), .B(n_289), .Y(n_336) );
INVx2_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
INVx1_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_265), .A2(n_417), .B1(n_434), .B2(n_437), .C(n_439), .Y(n_433) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_266), .B(n_315), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_267), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g358 ( .A(n_267), .B(n_304), .Y(n_358) );
INVx3_ASAP7_75t_SL g399 ( .A(n_267), .Y(n_399) );
AND2x2_ASAP7_75t_L g343 ( .A(n_268), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g372 ( .A(n_268), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_268), .B(n_281), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_268), .B(n_327), .Y(n_413) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g315 ( .A(n_269), .Y(n_315) );
OAI322xp33_ASAP7_75t_L g410 ( .A1(n_269), .A2(n_341), .A3(n_363), .B1(n_411), .B2(n_413), .C1(n_414), .C2(n_415), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_276), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_280), .A2(n_283), .B(n_435), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g360 ( .A(n_281), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g382 ( .A(n_281), .B(n_294), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_281), .B(n_321), .Y(n_397) );
INVxp67_ASAP7_75t_L g348 ( .A(n_283), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g354 ( .A1(n_283), .A2(n_355), .B(n_359), .C(n_369), .Y(n_354) );
OAI221xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_293), .B1(n_296), .B2(n_300), .C(n_305), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g425 ( .A(n_292), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_293), .A2(n_442), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_441) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_294), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g341 ( .A(n_294), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_294), .B(n_372), .Y(n_379) );
AND2x2_ASAP7_75t_L g421 ( .A(n_294), .B(n_399), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_295), .B(n_320), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_295), .A2(n_307), .B1(n_417), .B2(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g447 ( .A(n_295), .B(n_315), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g424 ( .A(n_298), .Y(n_424) );
AND2x2_ASAP7_75t_L g449 ( .A(n_298), .B(n_392), .Y(n_449) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_SL g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g313 ( .A(n_303), .B(n_314), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_316), .B2(n_319), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g380 ( .A(n_308), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_308), .B(n_348), .Y(n_415) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_310), .A2(n_340), .A3(n_342), .B1(n_343), .B2(n_345), .C1(n_346), .C2(n_350), .Y(n_339) );
INVxp67_ASAP7_75t_L g333 ( .A(n_311), .Y(n_333) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_313), .A2(n_318), .B1(n_335), .B2(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_314), .B(n_327), .Y(n_414) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_315), .B(n_353), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_315), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g411 ( .A(n_317), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND3xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_339), .C(n_354), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_330), .B2(n_332), .C(n_334), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_326), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g340 ( .A(n_331), .B(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_333), .Y(n_412) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_338), .B(n_352), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_341), .B(n_399), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_342), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g417 ( .A(n_345), .Y(n_417) );
AND2x2_ASAP7_75t_L g432 ( .A(n_345), .B(n_409), .Y(n_432) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_356), .A2(n_427), .B(n_433), .C(n_441), .Y(n_426) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g395 ( .A(n_366), .B(n_396), .Y(n_395) );
NAND2x1_ASAP7_75t_SL g437 ( .A(n_367), .B(n_438), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_370), .Y(n_407) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
AND2x2_ASAP7_75t_L g406 ( .A(n_376), .B(n_392), .Y(n_406) );
NOR5xp2_ASAP7_75t_L g377 ( .A(n_378), .B(n_393), .C(n_410), .D(n_416), .E(n_419), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_381), .B2(n_383), .C(n_385), .Y(n_378) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_382), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g408 ( .A(n_392), .B(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
AOI211xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B(n_424), .C(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx14_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g739 ( .A(n_455), .Y(n_739) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_456), .B(n_659), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_617), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_557), .C(n_593), .D(n_607), .Y(n_457) );
OAI221xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_505), .B1(n_535), .B2(n_544), .C(n_548), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_459), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_485), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
AND2x2_ASAP7_75t_L g554 ( .A(n_462), .B(n_474), .Y(n_554) );
INVx3_ASAP7_75t_L g562 ( .A(n_462), .Y(n_562) );
AND2x2_ASAP7_75t_L g616 ( .A(n_462), .B(n_488), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_462), .B(n_487), .Y(n_652) );
AND2x2_ASAP7_75t_L g710 ( .A(n_462), .B(n_572), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_471), .Y(n_467) );
INVx2_ASAP7_75t_L g481 ( .A(n_470), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_471), .A2(n_481), .B(n_495), .C(n_496), .Y(n_494) );
AND2x2_ASAP7_75t_L g545 ( .A(n_473), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g559 ( .A(n_473), .B(n_488), .Y(n_559) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_474), .B(n_488), .Y(n_574) );
AND2x2_ASAP7_75t_L g586 ( .A(n_474), .B(n_562), .Y(n_586) );
OR2x2_ASAP7_75t_L g588 ( .A(n_474), .B(n_546), .Y(n_588) );
AND2x2_ASAP7_75t_L g623 ( .A(n_474), .B(n_546), .Y(n_623) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_474), .Y(n_668) );
INVx1_ASAP7_75t_L g676 ( .A(n_474), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_483), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_485), .A2(n_594), .B1(n_598), .B2(n_602), .C(n_603), .Y(n_593) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
INVx2_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
AND2x2_ASAP7_75t_L g605 ( .A(n_487), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g624 ( .A(n_487), .B(n_562), .Y(n_624) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g687 ( .A(n_488), .B(n_562), .Y(n_687) );
AND2x2_ASAP7_75t_L g609 ( .A(n_498), .B(n_554), .Y(n_609) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_498), .A2(n_633), .A3(n_678), .B1(n_680), .B2(n_683), .C1(n_685), .C2(n_689), .Y(n_677) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_499), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g573 ( .A(n_499), .Y(n_573) );
AND2x2_ASAP7_75t_L g682 ( .A(n_499), .B(n_562), .Y(n_682) );
AND2x2_ASAP7_75t_L g714 ( .A(n_499), .B(n_586), .Y(n_714) );
OR2x2_ASAP7_75t_L g717 ( .A(n_499), .B(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g547 ( .A(n_500), .Y(n_547) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
INVx1_ASAP7_75t_L g730 ( .A(n_507), .Y(n_730) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g537 ( .A(n_508), .B(n_525), .Y(n_537) );
INVx2_ASAP7_75t_L g570 ( .A(n_508), .Y(n_570) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g592 ( .A(n_509), .Y(n_592) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_509), .Y(n_600) );
OR2x2_ASAP7_75t_L g724 ( .A(n_509), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g549 ( .A(n_518), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g589 ( .A(n_518), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g641 ( .A(n_518), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g538 ( .A(n_519), .B(n_539), .Y(n_538) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_519), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g650 ( .A(n_519), .B(n_540), .Y(n_650) );
OR2x2_ASAP7_75t_L g658 ( .A(n_519), .B(n_592), .Y(n_658) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_520), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g601 ( .A(n_520), .B(n_525), .Y(n_601) );
AND2x2_ASAP7_75t_L g665 ( .A(n_520), .B(n_540), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_525), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_525), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g578 ( .A(n_525), .Y(n_578) );
INVx1_ASAP7_75t_L g583 ( .A(n_525), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_525), .B(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_525), .Y(n_673) );
INVx1_ASAP7_75t_L g725 ( .A(n_525), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_530), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g702 ( .A(n_536), .B(n_611), .Y(n_702) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g629 ( .A(n_538), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g728 ( .A(n_538), .B(n_663), .Y(n_728) );
INVx1_ASAP7_75t_L g550 ( .A(n_539), .Y(n_550) );
AND2x2_ASAP7_75t_L g576 ( .A(n_539), .B(n_570), .Y(n_576) );
BUFx2_ASAP7_75t_L g635 ( .A(n_539), .Y(n_635) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_540), .Y(n_556) );
INVx1_ASAP7_75t_L g566 ( .A(n_540), .Y(n_566) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_544), .B(n_551), .Y(n_704) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI32xp33_ASAP7_75t_L g548 ( .A1(n_545), .A2(n_549), .A3(n_551), .B1(n_553), .B2(n_555), .Y(n_548) );
AND2x2_ASAP7_75t_L g688 ( .A(n_545), .B(n_561), .Y(n_688) );
AND2x2_ASAP7_75t_L g726 ( .A(n_545), .B(n_624), .Y(n_726) );
INVx1_ASAP7_75t_L g606 ( .A(n_546), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_550), .B(n_612), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_551), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_551), .B(n_554), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_551), .B(n_623), .Y(n_705) );
OR2x2_ASAP7_75t_L g719 ( .A(n_551), .B(n_588), .Y(n_719) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_554), .Y(n_646) );
OR2x2_ASAP7_75t_L g655 ( .A(n_552), .B(n_642), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_554), .B(n_605), .Y(n_627) );
INVx2_ASAP7_75t_L g642 ( .A(n_556), .Y(n_642) );
OR2x2_ASAP7_75t_L g657 ( .A(n_556), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g672 ( .A(n_556), .B(n_673), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_556), .A2(n_649), .B(n_730), .C(n_731), .Y(n_729) );
OAI321xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_563), .A3(n_568), .B1(n_571), .B2(n_575), .C(n_579), .Y(n_557) );
INVx1_ASAP7_75t_L g670 ( .A(n_558), .Y(n_670) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g681 ( .A(n_559), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_562), .B(n_676), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_563), .A2(n_701), .B1(n_703), .B2(n_705), .C(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x2_ASAP7_75t_L g638 ( .A(n_565), .B(n_612), .Y(n_638) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_566), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g611 ( .A(n_567), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_568), .A2(n_609), .B(n_654), .C(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g620 ( .A(n_570), .B(n_577), .Y(n_620) );
BUFx2_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
INVx1_ASAP7_75t_L g645 ( .A(n_570), .Y(n_645) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
OR2x2_ASAP7_75t_L g651 ( .A(n_573), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g734 ( .A(n_573), .Y(n_734) );
INVx1_ASAP7_75t_L g727 ( .A(n_574), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g580 ( .A(n_576), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g684 ( .A(n_576), .B(n_601), .Y(n_684) );
INVx1_ASAP7_75t_L g613 ( .A(n_577), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B1(n_587), .B2(n_589), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_581), .B(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g649 ( .A(n_582), .B(n_650), .Y(n_649) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_583), .B(n_592), .Y(n_612) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g604 ( .A(n_586), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g614 ( .A(n_588), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_591), .A2(n_709), .B1(n_711), .B2(n_712), .C(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g597 ( .A(n_592), .Y(n_597) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_592), .Y(n_663) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_595), .B(n_714), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_596), .A2(n_601), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_599), .B(n_609), .Y(n_706) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g675 ( .A(n_600), .Y(n_675) );
AND2x2_ASAP7_75t_L g634 ( .A(n_601), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g723 ( .A(n_601), .Y(n_723) );
INVx1_ASAP7_75t_L g639 ( .A(n_604), .Y(n_639) );
INVx1_ASAP7_75t_L g694 ( .A(n_605), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_613), .B2(n_614), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_611), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g679 ( .A(n_612), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_612), .B(n_650), .Y(n_716) );
OR2x2_ASAP7_75t_L g689 ( .A(n_613), .B(n_642), .Y(n_689) );
INVx1_ASAP7_75t_L g628 ( .A(n_614), .Y(n_628) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_616), .B(n_667), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_636), .C(n_647), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_625), .C(n_631), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_620), .A2(n_691), .B1(n_695), .B2(n_698), .C(n_700), .Y(n_690) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g632 ( .A(n_623), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g686 ( .A(n_623), .B(n_687), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g671 ( .A1(n_624), .A2(n_672), .B(n_674), .C(n_676), .Y(n_671) );
INVx2_ASAP7_75t_L g718 ( .A(n_624), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_628), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g697 ( .A(n_630), .B(n_650), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_639), .B(n_640), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_643), .B(n_646), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_641), .B(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_646), .B(n_733), .Y(n_732) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_653), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g674 ( .A(n_650), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND4x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_690), .C(n_707), .D(n_729), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_677), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_666), .B(n_669), .C(n_671), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_665), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_676), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g711 ( .A(n_686), .Y(n_711) );
INVx2_ASAP7_75t_SL g699 ( .A(n_687), .Y(n_699) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g712 ( .A(n_697), .Y(n_712) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_715), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
OAI221xp5_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g740 ( .A(n_736), .Y(n_740) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
endmodule