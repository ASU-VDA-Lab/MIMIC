module fake_netlist_6_2748_n_1671 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1671);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1671;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_102),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_24),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_34),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_48),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_38),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_6),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_6),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_38),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_85),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_42),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_45),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_26),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_41),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_74),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_28),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_103),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_44),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_4),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

INVxp33_ASAP7_75t_R g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_9),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_108),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_28),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_69),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_59),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_47),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_68),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_58),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_32),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_110),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_137),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_51),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_87),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_80),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_122),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_124),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_62),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_94),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_65),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_145),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_116),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_21),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_34),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_5),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_40),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_70),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_88),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_86),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_119),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_7),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_39),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_54),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_22),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_66),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_15),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_13),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_111),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_52),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_46),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_53),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_146),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_22),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_27),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_13),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_140),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_71),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_44),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_96),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_75),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_115),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_1),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_64),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_26),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_27),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_84),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_35),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_50),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_9),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_24),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_0),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_30),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_12),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_25),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_77),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_23),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_37),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_61),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_20),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_43),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_12),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_107),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_183),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_183),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_160),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_183),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_153),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_183),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_155),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_156),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_161),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_183),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_183),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_166),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_215),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_206),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_206),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_206),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_175),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_206),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_206),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_158),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_160),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_206),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_173),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_167),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_160),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_167),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_163),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_260),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_215),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_235),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_235),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_171),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_179),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_170),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_181),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_168),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_181),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_182),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_263),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_185),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_187),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_168),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_188),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_178),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_186),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_234),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_182),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_238),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_244),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_193),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_349),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_170),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_307),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_309),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_317),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_310),
.B(n_229),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_209),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_311),
.B(n_209),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_315),
.B(n_301),
.Y(n_389)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_302),
.A2(n_257),
.B(n_164),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_361),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_323),
.B(n_301),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_302),
.B(n_174),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_303),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_229),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_303),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_326),
.A2(n_217),
.B1(n_299),
.B2(n_267),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_306),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_358),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_306),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_312),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_312),
.A2(n_257),
.B(n_164),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_313),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_359),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_314),
.B(n_262),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_314),
.B(n_262),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_318),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_329),
.A2(n_290),
.B1(n_245),
.B2(n_296),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_298),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_319),
.A2(n_293),
.B(n_162),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_248),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_343),
.B(n_255),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_293),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_316),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_321),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_324),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g433 ( 
.A1(n_325),
.A2(n_165),
.B(n_159),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_339),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_328),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_328),
.B(n_169),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_331),
.B(n_172),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_385),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_386),
.B(n_341),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_387),
.B(n_367),
.Y(n_454)
);

BUFx6f_ASAP7_75t_SL g455 ( 
.A(n_393),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_378),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_426),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_406),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_331),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_336),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_437),
.A2(n_304),
.B1(n_353),
.B2(n_286),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_305),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g465 ( 
.A1(n_409),
.A2(n_189),
.B(n_180),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_332),
.C(n_327),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_428),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

OAI22xp33_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_251),
.B1(n_290),
.B2(n_231),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_375),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_389),
.B(n_345),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_378),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_428),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_396),
.B(n_333),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_430),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_410),
.Y(n_482)
);

AO22x2_ASAP7_75t_L g483 ( 
.A1(n_376),
.A2(n_274),
.B1(n_288),
.B2(n_294),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_407),
.Y(n_484)
);

BUFx6f_ASAP7_75t_SL g485 ( 
.A(n_393),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_SL g486 ( 
.A1(n_409),
.A2(n_338),
.B(n_333),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_431),
.B(n_364),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_418),
.A2(n_395),
.B1(n_438),
.B2(n_431),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_438),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_411),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_415),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_393),
.B(n_201),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_432),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_415),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_375),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_421),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_375),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_338),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_435),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_417),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_420),
.B(n_367),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_417),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_413),
.B(n_340),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_407),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_401),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_401),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_407),
.Y(n_527)
);

CKINVDCx11_ASAP7_75t_R g528 ( 
.A(n_405),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_417),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_413),
.B(n_340),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_401),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_372),
.Y(n_533)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_387),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_372),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_382),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_373),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_407),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_387),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_420),
.B(n_354),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_405),
.B(n_207),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_373),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_402),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_377),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_391),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_422),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_377),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_391),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_391),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_380),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_391),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_391),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_380),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_413),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_405),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_383),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_413),
.B(n_219),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_383),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_397),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_397),
.Y(n_564)
);

XOR2x2_ASAP7_75t_SL g565 ( 
.A(n_416),
.B(n_217),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_397),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_397),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_397),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_422),
.A2(n_211),
.B1(n_221),
.B2(n_157),
.Y(n_569)
);

AND3x2_ASAP7_75t_L g570 ( 
.A(n_414),
.B(n_232),
.C(n_191),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_414),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_387),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_397),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_437),
.B(n_207),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_404),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_437),
.B(n_184),
.C(n_176),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_404),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_404),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_414),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_398),
.B(n_174),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_419),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_439),
.A2(n_295),
.B1(n_174),
.B2(n_370),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_419),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_551),
.A2(n_439),
.B(n_390),
.Y(n_586)
);

NOR2xp67_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_414),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_558),
.B(n_439),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_578),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_441),
.B(n_439),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_558),
.B(n_404),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_571),
.B(n_404),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_433),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_450),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_551),
.A2(n_433),
.B1(n_390),
.B2(n_267),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_534),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_474),
.B(n_462),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_487),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_551),
.B(n_174),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_578),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_460),
.A2(n_241),
.B1(n_292),
.B2(n_224),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_459),
.B(n_224),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_548),
.B(n_347),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_464),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_433),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_461),
.B(n_561),
.C(n_487),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_514),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_454),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_580),
.B(n_478),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_466),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_514),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_559),
.B(n_242),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_454),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_493),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_458),
.B(n_390),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_458),
.B(n_390),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_523),
.B(n_364),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_467),
.B(n_398),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

INVx8_ASAP7_75t_L g623 ( 
.A(n_455),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_456),
.A2(n_241),
.B1(n_292),
.B2(n_355),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_467),
.B(n_398),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_521),
.A2(n_190),
.B(n_276),
.C(n_275),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_442),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_455),
.Y(n_628)
);

NAND2x1p5_ASAP7_75t_L g629 ( 
.A(n_456),
.B(n_192),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_488),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_470),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_468),
.B(n_398),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_572),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_442),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_468),
.B(n_398),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_530),
.B(n_194),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_444),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_582),
.B(n_210),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_507),
.B(n_213),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_477),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_483),
.A2(n_299),
.B1(n_230),
.B2(n_239),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_582),
.A2(n_226),
.B(n_268),
.C(n_270),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_479),
.B(n_398),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_455),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_479),
.B(n_240),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_SL g647 ( 
.A(n_485),
.B(n_368),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_480),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_541),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_444),
.A2(n_394),
.B(n_392),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_507),
.B(n_243),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_440),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_541),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_488),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_482),
.B(n_249),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_488),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_534),
.Y(n_657)
);

BUFx5_ASAP7_75t_L g658 ( 
.A(n_585),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_482),
.B(n_252),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_446),
.B(n_264),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_453),
.B(n_271),
.Y(n_661)
);

BUFx12f_ASAP7_75t_L g662 ( 
.A(n_536),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_534),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_510),
.B(n_197),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_451),
.B(n_365),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_489),
.B(n_392),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_576),
.B(n_476),
.C(n_491),
.Y(n_667)
);

OAI221xp5_ASAP7_75t_L g668 ( 
.A1(n_583),
.A2(n_365),
.B1(n_370),
.B2(n_369),
.C(n_366),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_574),
.B(n_154),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_570),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_540),
.A2(n_208),
.B1(n_297),
.B2(n_287),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_483),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_540),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_510),
.B(n_203),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_481),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_492),
.B(n_394),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_494),
.B(n_154),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_512),
.B(n_204),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_497),
.B(n_237),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_483),
.A2(n_298),
.B1(n_300),
.B2(n_273),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_483),
.Y(n_681)
);

BUFx5_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_569),
.B(n_237),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_500),
.B(n_247),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_451),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_502),
.B(n_205),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_508),
.B(n_212),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_511),
.B(n_247),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_513),
.B(n_214),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_516),
.B(n_216),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_572),
.B(n_218),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_517),
.B(n_220),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_540),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_536),
.B(n_273),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_512),
.B(n_222),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_572),
.B(n_223),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_522),
.B(n_225),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_465),
.A2(n_300),
.B1(n_369),
.B2(n_366),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_465),
.A2(n_266),
.B1(n_196),
.B2(n_198),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_543),
.B(n_195),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_536),
.B(n_256),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_227),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_518),
.B(n_228),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_498),
.B(n_354),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_465),
.A2(n_272),
.B1(n_202),
.B2(n_233),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_520),
.B(n_246),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_522),
.B(n_531),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_520),
.B(n_253),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_472),
.B(n_200),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_545),
.A2(n_278),
.B1(n_250),
.B2(n_258),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_524),
.B(n_236),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_524),
.B(n_279),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_531),
.B(n_254),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_525),
.B(n_526),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_445),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_525),
.B(n_269),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_526),
.B(n_259),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_495),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_533),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_445),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_545),
.A2(n_261),
.B1(n_282),
.B2(n_277),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_532),
.B(n_281),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_486),
.A2(n_283),
.B(n_285),
.C(n_357),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_447),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_485),
.Y(n_726)
);

INVx4_ASAP7_75t_SL g727 ( 
.A(n_485),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_533),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_447),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_532),
.B(n_291),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_542),
.B(n_362),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_448),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_448),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_449),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_535),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_469),
.B(n_362),
.C(n_360),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_449),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_484),
.A2(n_360),
.B1(n_357),
.B2(n_356),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_527),
.B(n_356),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_535),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_527),
.B(n_539),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_538),
.B(n_150),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_598),
.B(n_542),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_598),
.B(n_504),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_586),
.A2(n_503),
.B(n_501),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_622),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_622),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_633),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_731),
.B(n_542),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_593),
.A2(n_608),
.B(n_612),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_590),
.B(n_537),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_716),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_587),
.B(n_506),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_652),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_611),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_633),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_616),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_685),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_720),
.Y(n_759)
);

NOR2x1p5_ASAP7_75t_L g760 ( 
.A(n_662),
.B(n_528),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_728),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_603),
.B(n_498),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_539),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_735),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_603),
.B(n_498),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_740),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_633),
.B(n_565),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_614),
.B(n_498),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_627),
.Y(n_769)
);

BUFx2_ASAP7_75t_SL g770 ( 
.A(n_685),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_590),
.A2(n_550),
.B1(n_547),
.B2(n_553),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_633),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_597),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_617),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_642),
.A2(n_549),
.B1(n_537),
.B2(n_544),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_596),
.B(n_544),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_649),
.B(n_565),
.Y(n_777)
);

BUFx12f_ASAP7_75t_L g778 ( 
.A(n_705),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_716),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_653),
.B(n_538),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_701),
.A2(n_556),
.B1(n_563),
.B2(n_566),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_635),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_638),
.Y(n_783)
);

NOR2x1p5_ASAP7_75t_L g784 ( 
.A(n_630),
.B(n_528),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_721),
.Y(n_785)
);

NOR2x1_ASAP7_75t_R g786 ( 
.A(n_654),
.B(n_440),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_599),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_725),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_729),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_732),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_656),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_600),
.B(n_538),
.Y(n_792)
);

AND2x6_ASAP7_75t_L g793 ( 
.A(n_618),
.B(n_501),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_733),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_665),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_596),
.B(n_546),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_647),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_623),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_609),
.B(n_549),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_715),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_600),
.B(n_538),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_619),
.B(n_503),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_620),
.B(n_554),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_734),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_737),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_658),
.B(n_682),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_594),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_623),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_658),
.B(n_554),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_589),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_595),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_658),
.B(n_557),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_658),
.B(n_557),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_601),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_667),
.B(n_727),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_672),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_658),
.B(n_560),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_606),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_658),
.B(n_682),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_727),
.B(n_560),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_705),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_701),
.B(n_562),
.C(n_581),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_628),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_666),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_682),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_615),
.B(n_562),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_628),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_676),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_682),
.B(n_496),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_615),
.B(n_538),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_604),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_682),
.B(n_499),
.Y(n_832)
);

AND3x1_ASAP7_75t_L g833 ( 
.A(n_602),
.B(n_496),
.C(n_499),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_629),
.B(n_575),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_669),
.B(n_581),
.C(n_564),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_682),
.B(n_519),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_739),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_628),
.B(n_577),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_639),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_629),
.B(n_555),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_605),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_695),
.B(n_555),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_699),
.B(n_519),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_727),
.B(n_568),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_708),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_607),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_708),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_669),
.B(n_555),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_645),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_712),
.A2(n_568),
.B(n_567),
.C(n_577),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_645),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_722),
.B(n_573),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_724),
.A2(n_564),
.B(n_573),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_681),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_613),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_645),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_657),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_705),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_726),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_686),
.B(n_555),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_588),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_710),
.B(n_509),
.Y(n_862)
);

AND2x6_ASAP7_75t_SL g863 ( 
.A(n_710),
.B(n_677),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_687),
.B(n_689),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_670),
.B(n_567),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_624),
.B(n_509),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_717),
.A2(n_509),
.B1(n_519),
.B2(n_552),
.Y(n_867)
);

INVx5_ASAP7_75t_L g868 ( 
.A(n_639),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_700),
.B(n_443),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_683),
.B(n_490),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_730),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_700),
.B(n_443),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_726),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_664),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_690),
.B(n_579),
.Y(n_875)
);

CKINVDCx8_ASAP7_75t_R g876 ( 
.A(n_726),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_639),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_642),
.A2(n_552),
.B1(n_443),
.B2(n_452),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_722),
.B(n_452),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_631),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_706),
.B(n_452),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_663),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_634),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_717),
.A2(n_490),
.B1(n_584),
.B2(n_515),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_L g885 ( 
.A(n_711),
.B(n_584),
.C(n_490),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_706),
.B(n_473),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_641),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_591),
.A2(n_584),
.B(n_473),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_648),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_693),
.B(n_579),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_643),
.A2(n_475),
.B(n_473),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_646),
.B(n_475),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_675),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_660),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_696),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_655),
.B(n_475),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_741),
.B(n_529),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_659),
.B(n_475),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_673),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_711),
.B(n_677),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_637),
.A2(n_475),
.B(n_473),
.C(n_575),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_712),
.B(n_579),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_719),
.B(n_473),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_691),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_694),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_736),
.B(n_579),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_713),
.B(n_529),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_592),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_713),
.B(n_529),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_661),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_592),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_900),
.A2(n_688),
.B(n_684),
.C(n_679),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_791),
.B(n_697),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_744),
.B(n_824),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_825),
.A2(n_697),
.B(n_692),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_774),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_755),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_SL g918 ( 
.A1(n_754),
.A2(n_680),
.B1(n_668),
.B2(n_702),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_826),
.A2(n_718),
.B(n_679),
.C(n_684),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_744),
.B(n_718),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_SL g921 ( 
.A1(n_862),
.A2(n_799),
.B(n_870),
.C(n_826),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_749),
.B(n_688),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_825),
.A2(n_505),
.B(n_515),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_816),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_806),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_862),
.A2(n_703),
.B1(n_723),
.B2(n_704),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_776),
.A2(n_680),
.B1(n_637),
.B2(n_625),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_748),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_777),
.A2(n_674),
.B1(n_678),
.B2(n_664),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_R g930 ( 
.A(n_851),
.B(n_639),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_750),
.A2(n_644),
.B(n_621),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_828),
.B(n_674),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_776),
.A2(n_636),
.B1(n_632),
.B2(n_742),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_852),
.A2(n_678),
.B1(n_714),
.B2(n_698),
.Y(n_934)
);

BUFx12f_ASAP7_75t_L g935 ( 
.A(n_859),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_806),
.A2(n_505),
.B(n_515),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_796),
.A2(n_742),
.B1(n_698),
.B2(n_714),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_800),
.B(n_709),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_871),
.B(n_837),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_795),
.B(n_736),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_816),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_743),
.B(n_707),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_819),
.A2(n_505),
.B(n_529),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_819),
.A2(n_505),
.B(n_529),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_757),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_799),
.A2(n_650),
.B(n_671),
.C(n_651),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_746),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_854),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_866),
.A2(n_651),
.B(n_640),
.C(n_626),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_750),
.A2(n_515),
.B(n_505),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_866),
.A2(n_640),
.B(n_738),
.C(n_639),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_787),
.B(n_575),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_787),
.B(n_575),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_751),
.A2(n_141),
.B(n_138),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_L g955 ( 
.A1(n_848),
.A2(n_135),
.B(n_134),
.C(n_132),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_854),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_769),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_748),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_767),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_959)
);

NAND3xp33_ASAP7_75t_SL g960 ( 
.A(n_762),
.B(n_2),
.C(n_4),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_803),
.A2(n_8),
.B(n_10),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_894),
.B(n_15),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_910),
.B(n_17),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_902),
.A2(n_82),
.B(n_127),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_895),
.B(n_18),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_818),
.B(n_19),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_797),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_809),
.A2(n_89),
.B(n_114),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_748),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_782),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_747),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_756),
.B(n_772),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_861),
.A2(n_19),
.B(n_20),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_756),
.B(n_93),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_756),
.B(n_63),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_747),
.Y(n_976)
);

AND2x6_ASAP7_75t_L g977 ( 
.A(n_820),
.B(n_95),
.Y(n_977)
);

OAI22x1_ASAP7_75t_L g978 ( 
.A1(n_765),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_796),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_772),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_758),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_874),
.A2(n_31),
.B(n_35),
.C(n_36),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_879),
.A2(n_36),
.B(n_40),
.C(n_97),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_772),
.B(n_99),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_880),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_869),
.A2(n_100),
.B(n_101),
.C(n_104),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_768),
.B(n_763),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_758),
.B(n_105),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_770),
.B(n_783),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_863),
.B(n_753),
.Y(n_990)
);

OA22x2_ASAP7_75t_L g991 ( 
.A1(n_768),
.A2(n_821),
.B1(n_858),
.B2(n_814),
.Y(n_991)
);

BUFx2_ASAP7_75t_SL g992 ( 
.A(n_798),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_886),
.A2(n_864),
.B(n_881),
.C(n_869),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_872),
.A2(n_881),
.B(n_886),
.C(n_908),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_810),
.B(n_865),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_809),
.A2(n_812),
.B(n_817),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_872),
.A2(n_842),
.B(n_759),
.C(n_761),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_764),
.A2(n_766),
.B(n_843),
.C(n_830),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_839),
.Y(n_999)
);

INVx3_ASAP7_75t_SL g1000 ( 
.A(n_873),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_775),
.A2(n_843),
.B1(n_878),
.B2(n_833),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_812),
.A2(n_817),
.B(n_813),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_865),
.B(n_763),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_883),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_815),
.B(n_820),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_873),
.B(n_798),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_SL g1007 ( 
.A(n_904),
.B(n_834),
.C(n_840),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_813),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_853),
.A2(n_890),
.B(n_875),
.C(n_860),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_SL g1010 ( 
.A(n_822),
.B(n_876),
.C(n_885),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_775),
.B(n_845),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_850),
.A2(n_822),
.B(n_909),
.C(n_907),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_773),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_887),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_778),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_906),
.A2(n_815),
.B1(n_847),
.B2(n_911),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_878),
.A2(n_839),
.B1(n_877),
.B2(n_868),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_907),
.A2(n_909),
.B(n_885),
.C(n_835),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_808),
.B(n_823),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_752),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_785),
.B(n_788),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_829),
.A2(n_832),
.B(n_836),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_789),
.B(n_790),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_829),
.A2(n_832),
.B(n_836),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_745),
.A2(n_901),
.B(n_802),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_839),
.A2(n_868),
.B1(n_877),
.B2(n_801),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_786),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_857),
.B(n_899),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_794),
.B(n_804),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_901),
.A2(n_793),
.B(n_802),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_808),
.B(n_849),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_823),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_855),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_823),
.Y(n_1034)
);

BUFx4f_ASAP7_75t_L g1035 ( 
.A(n_827),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_889),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_792),
.A2(n_805),
.B(n_893),
.C(n_811),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_857),
.B(n_882),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_899),
.B(n_905),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_779),
.B(n_846),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_905),
.B(n_807),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_827),
.B(n_849),
.Y(n_1042)
);

BUFx4_ASAP7_75t_SL g1043 ( 
.A(n_838),
.Y(n_1043)
);

NAND2xp33_ASAP7_75t_SL g1044 ( 
.A(n_827),
.B(n_849),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_831),
.B(n_841),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_903),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_916),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_957),
.Y(n_1048)
);

OA22x2_ASAP7_75t_L g1049 ( 
.A1(n_978),
.A2(n_781),
.B1(n_838),
.B2(n_897),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_914),
.B(n_856),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_967),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_920),
.B(n_898),
.Y(n_1052)
);

NAND2x1p5_ASAP7_75t_L g1053 ( 
.A(n_1035),
.B(n_856),
.Y(n_1053)
);

AOI221xp5_ASAP7_75t_L g1054 ( 
.A1(n_918),
.A2(n_892),
.B1(n_896),
.B2(n_898),
.C(n_771),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_938),
.B(n_896),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_SL g1056 ( 
.A(n_919),
.B(n_892),
.C(n_884),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_947),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1018),
.A2(n_802),
.B(n_793),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_SL g1059 ( 
.A1(n_998),
.A2(n_891),
.B(n_888),
.Y(n_1059)
);

NAND2x1_ASAP7_75t_L g1060 ( 
.A(n_1013),
.B(n_773),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_SL g1061 ( 
.A1(n_959),
.A2(n_867),
.B(n_844),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_917),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_1035),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_1025),
.A2(n_888),
.B(n_903),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_945),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_970),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_R g1067 ( 
.A(n_930),
.B(n_844),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_939),
.B(n_802),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_912),
.A2(n_868),
.B(n_839),
.C(n_877),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_971),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_992),
.B(n_873),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_993),
.A2(n_793),
.B(n_802),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_926),
.A2(n_897),
.B(n_780),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_922),
.B(n_838),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_994),
.A2(n_793),
.A3(n_784),
.B(n_760),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_937),
.A2(n_793),
.B(n_932),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1016),
.A2(n_1008),
.B1(n_1017),
.B2(n_929),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_1001),
.A2(n_937),
.A3(n_927),
.B(n_973),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1017),
.A2(n_1039),
.B1(n_995),
.B2(n_1041),
.Y(n_1079)
);

AOI221x1_ASAP7_75t_L g1080 ( 
.A1(n_1010),
.A2(n_979),
.B1(n_1001),
.B2(n_983),
.C(n_1030),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_915),
.A2(n_950),
.B(n_996),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1003),
.B(n_942),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_940),
.B(n_966),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1034),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1012),
.A2(n_1009),
.B(n_1024),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_936),
.A2(n_943),
.B(n_944),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_976),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1019),
.B(n_1031),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_960),
.A2(n_961),
.B1(n_990),
.B2(n_965),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1002),
.A2(n_1025),
.B(n_921),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_999),
.A2(n_1022),
.B(n_946),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_931),
.A2(n_933),
.B(n_951),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_981),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_1015),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1046),
.B(n_1011),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_962),
.B(n_963),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1020),
.B(n_924),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_989),
.B(n_941),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_948),
.B(n_956),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1033),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_927),
.A2(n_949),
.A3(n_933),
.B(n_979),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_991),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_986),
.A2(n_923),
.A3(n_1026),
.B(n_982),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_954),
.A2(n_1028),
.A3(n_1038),
.B(n_968),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_987),
.B(n_1036),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1021),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_964),
.A2(n_997),
.B(n_1037),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_913),
.B(n_988),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_985),
.B(n_1004),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_969),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_999),
.A2(n_934),
.B(n_1013),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_SL g1113 ( 
.A1(n_1023),
.A2(n_1029),
.B1(n_1045),
.B2(n_1005),
.C(n_953),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_977),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_SL g1115 ( 
.A1(n_974),
.A2(n_984),
.B(n_975),
.C(n_928),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1014),
.B(n_952),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1007),
.A2(n_1040),
.B1(n_972),
.B2(n_958),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_969),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_955),
.A2(n_972),
.B(n_958),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1044),
.A2(n_1042),
.B(n_928),
.C(n_1032),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_SL g1121 ( 
.A(n_977),
.B(n_935),
.Y(n_1121)
);

AOI221x1_ASAP7_75t_L g1122 ( 
.A1(n_969),
.A2(n_980),
.B1(n_1043),
.B2(n_977),
.C(n_1027),
.Y(n_1122)
);

AO21x2_ASAP7_75t_L g1123 ( 
.A1(n_977),
.A2(n_980),
.B(n_1006),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_977),
.B(n_980),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1006),
.B(n_1000),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_920),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_920),
.B(n_598),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_947),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1018),
.A2(n_994),
.A3(n_1001),
.B(n_919),
.Y(n_1129)
);

AND2x6_ASAP7_75t_L g1130 ( 
.A(n_1013),
.B(n_820),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1131)
);

OA21x2_ASAP7_75t_L g1132 ( 
.A1(n_1025),
.A2(n_1030),
.B(n_1018),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1035),
.Y(n_1133)
);

AO32x2_ASAP7_75t_L g1134 ( 
.A1(n_1001),
.A2(n_979),
.A3(n_927),
.B1(n_937),
.B2(n_672),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1013),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1018),
.A2(n_994),
.A3(n_1001),
.B(n_919),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_919),
.A2(n_900),
.B(n_598),
.C(n_912),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1018),
.A2(n_825),
.B(n_819),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_SL g1140 ( 
.A(n_930),
.B(n_1000),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_920),
.B(n_598),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_L g1142 ( 
.A1(n_919),
.A2(n_598),
.B(n_900),
.C(n_912),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_947),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_967),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_957),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_947),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_919),
.A2(n_598),
.B(n_900),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_919),
.A2(n_900),
.B(n_598),
.C(n_912),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_916),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1018),
.A2(n_825),
.B(n_819),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_919),
.A2(n_900),
.B(n_598),
.C(n_912),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_1006),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_917),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_947),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1018),
.A2(n_919),
.B(n_993),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_919),
.B(n_598),
.C(n_602),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_947),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_919),
.A2(n_900),
.B(n_598),
.C(n_912),
.Y(n_1158)
);

OAI22x1_ASAP7_75t_L g1159 ( 
.A1(n_990),
.A2(n_900),
.B1(n_598),
.B2(n_602),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1017),
.A2(n_825),
.B(n_925),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_920),
.B(n_598),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1163)
);

OAI22x1_ASAP7_75t_L g1164 ( 
.A1(n_990),
.A2(n_900),
.B1(n_598),
.B2(n_602),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_947),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_920),
.B(n_598),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_940),
.B(n_749),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_950),
.A2(n_745),
.B(n_936),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_938),
.B(n_871),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1035),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_925),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1018),
.A2(n_825),
.B(n_819),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1019),
.B(n_1031),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_940),
.B(n_749),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_920),
.B(n_598),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_920),
.B(n_598),
.Y(n_1179)
);

AO32x2_ASAP7_75t_L g1180 ( 
.A1(n_1001),
.A2(n_979),
.A3(n_927),
.B1(n_937),
.B2(n_672),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1018),
.A2(n_825),
.B(n_819),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1159),
.A2(n_1164),
.B1(n_1147),
.B2(n_1156),
.C(n_1148),
.Y(n_1182)
);

NAND2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1152),
.B(n_1114),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1081),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1133),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1131),
.A2(n_1161),
.B(n_1138),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1048),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1066),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1145),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1133),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1163),
.A2(n_1166),
.B(n_1165),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1083),
.B(n_1170),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1123),
.B(n_1114),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1082),
.B(n_1096),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1127),
.A2(n_1141),
.B1(n_1178),
.B2(n_1179),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1133),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1123),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1169),
.A2(n_1171),
.B(n_1108),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1059),
.A2(n_1085),
.B(n_1090),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1167),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1100),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1085),
.A2(n_1072),
.B(n_1058),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1072),
.A2(n_1058),
.B(n_1139),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1177),
.B(n_1126),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1152),
.B(n_1063),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1092),
.A2(n_1155),
.B(n_1076),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1119),
.A2(n_1150),
.B(n_1175),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1142),
.A2(n_1113),
.B(n_1137),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1062),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1065),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1128),
.B(n_1097),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1181),
.A2(n_1112),
.B(n_1073),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1151),
.A2(n_1158),
.A3(n_1077),
.B(n_1069),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1153),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1152),
.B(n_1088),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1113),
.A2(n_1054),
.B(n_1068),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1162),
.A2(n_1168),
.B(n_1089),
.C(n_1174),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1088),
.B(n_1176),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1089),
.A2(n_1109),
.B1(n_1079),
.B2(n_1056),
.C(n_1098),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1110),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1157),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1176),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1173),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_1055),
.A2(n_1052),
.B(n_1074),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1064),
.A2(n_1115),
.B(n_1132),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1105),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1099),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1132),
.A2(n_1117),
.B(n_1049),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1124),
.A2(n_1060),
.B(n_1095),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1050),
.B(n_1154),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1107),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_1143),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1106),
.A2(n_1102),
.B1(n_1061),
.B2(n_1093),
.C(n_1087),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_SL g1234 ( 
.A1(n_1116),
.A2(n_1061),
.B(n_1122),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1051),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1130),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1135),
.B(n_1173),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1118),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1134),
.A2(n_1180),
.B(n_1078),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1172),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1172),
.A2(n_1120),
.B(n_1087),
.C(n_1094),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1121),
.A2(n_1130),
.B(n_1135),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1078),
.A2(n_1180),
.A3(n_1134),
.B(n_1101),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1130),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1053),
.A2(n_1125),
.B(n_1104),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1104),
.A2(n_1103),
.B(n_1129),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1173),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1121),
.A2(n_1101),
.B(n_1134),
.C(n_1180),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1070),
.B(n_1149),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1129),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1136),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1075),
.A2(n_1130),
.B(n_1067),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1075),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1111),
.A2(n_1144),
.B(n_1071),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1084),
.B(n_1111),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1140),
.A2(n_1071),
.B(n_1047),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1071),
.A2(n_1086),
.B(n_1091),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1048),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1147),
.A2(n_598),
.B(n_919),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1048),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1081),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1123),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1174),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1080),
.A2(n_1090),
.A3(n_1148),
.B(n_1137),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1051),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1146),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1147),
.A2(n_598),
.B(n_912),
.C(n_900),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1080),
.A2(n_1090),
.B(n_1092),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1133),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1152),
.B(n_1114),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1127),
.A2(n_598),
.B1(n_602),
.B2(n_900),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1123),
.B(n_1114),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1048),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1048),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1127),
.B(n_598),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1127),
.B(n_1141),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1048),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1091),
.A2(n_1160),
.B(n_825),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1127),
.B(n_1141),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1147),
.A2(n_598),
.B(n_912),
.C(n_900),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1081),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1127),
.B(n_1141),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1080),
.A2(n_1090),
.A3(n_1148),
.B(n_1137),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_1072),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1048),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1156),
.A2(n_900),
.B1(n_1147),
.B2(n_598),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1083),
.B(n_1170),
.Y(n_1287)
);

BUFx8_ASAP7_75t_L g1288 ( 
.A(n_1133),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1048),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1127),
.B(n_598),
.Y(n_1290)
);

CKINVDCx8_ASAP7_75t_R g1291 ( 
.A(n_1051),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1081),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1127),
.B(n_598),
.Y(n_1293)
);

BUFx8_ASAP7_75t_L g1294 ( 
.A(n_1133),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1048),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1156),
.A2(n_900),
.B1(n_1147),
.B2(n_598),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_1072),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1147),
.B(n_598),
.C(n_900),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1156),
.A2(n_900),
.B1(n_1147),
.B2(n_598),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1133),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1048),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1263),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1204),
.B(n_1211),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1192),
.B(n_1287),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_L g1305 ( 
.A(n_1240),
.B(n_1235),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1193),
.B(n_1272),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1222),
.B(n_1218),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1221),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1266),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1235),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1194),
.B(n_1195),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_L g1312 ( 
.A(n_1200),
.B(n_1249),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1286),
.A2(n_1296),
.B1(n_1299),
.B2(n_1290),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1201),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1267),
.A2(n_1280),
.B(n_1217),
.C(n_1286),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1273),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1220),
.B(n_1230),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1299),
.A2(n_1293),
.B1(n_1290),
.B2(n_1275),
.Y(n_1318)
);

AOI211xp5_ASAP7_75t_L g1319 ( 
.A1(n_1182),
.A2(n_1219),
.B(n_1275),
.C(n_1293),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1230),
.B(n_1227),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1215),
.B(n_1231),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1265),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1276),
.B(n_1279),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1282),
.A2(n_1217),
.B1(n_1233),
.B2(n_1241),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1215),
.B(n_1209),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1248),
.A2(n_1212),
.B(n_1203),
.C(n_1202),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1263),
.B(n_1273),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1242),
.A2(n_1205),
.B(n_1254),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1277),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1224),
.B(n_1234),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1209),
.B(n_1226),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1255),
.A2(n_1232),
.B(n_1248),
.C(n_1238),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1197),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1210),
.B(n_1214),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1225),
.A2(n_1199),
.B(n_1203),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1289),
.B(n_1295),
.Y(n_1336)
);

AOI221x1_ASAP7_75t_SL g1337 ( 
.A1(n_1232),
.A2(n_1260),
.B1(n_1258),
.B2(n_1274),
.C(n_1285),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1295),
.B(n_1301),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1223),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1288),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1225),
.A2(n_1184),
.B(n_1281),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1223),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1253),
.A2(n_1197),
.B(n_1262),
.C(n_1250),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1188),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1189),
.A2(n_1268),
.B(n_1206),
.C(n_1183),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1265),
.Y(n_1346)
);

OA22x2_ASAP7_75t_L g1347 ( 
.A1(n_1228),
.A2(n_1256),
.B1(n_1252),
.B2(n_1245),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1237),
.B(n_1256),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1237),
.B(n_1245),
.Y(n_1349)
);

O2A1O1Ixp5_ASAP7_75t_L g1350 ( 
.A1(n_1253),
.A2(n_1251),
.B(n_1236),
.C(n_1244),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1183),
.A2(n_1270),
.B(n_1185),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1246),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1264),
.B(n_1283),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1264),
.B(n_1283),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1185),
.B(n_1300),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1291),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1216),
.B(n_1213),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1288),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1190),
.B(n_1300),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1184),
.A2(n_1292),
.B(n_1281),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1190),
.B(n_1269),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1261),
.A2(n_1292),
.B(n_1207),
.Y(n_1362)
);

AOI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1284),
.A2(n_1297),
.B1(n_1247),
.B2(n_1269),
.C(n_1236),
.Y(n_1363)
);

INVxp33_ASAP7_75t_L g1364 ( 
.A(n_1229),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1246),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_SL g1366 ( 
.A1(n_1208),
.A2(n_1294),
.B(n_1288),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1270),
.A2(n_1244),
.B(n_1239),
.C(n_1213),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1196),
.A2(n_1239),
.B1(n_1294),
.B2(n_1243),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1257),
.A2(n_1186),
.B(n_1191),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1196),
.B(n_1294),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1198),
.A2(n_900),
.B(n_1147),
.C(n_598),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1239),
.A2(n_1278),
.B(n_1259),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1243),
.B(n_1192),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1243),
.A2(n_598),
.B(n_912),
.C(n_1271),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1243),
.B(n_1192),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1286),
.A2(n_598),
.B1(n_602),
.B2(n_900),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1187),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1204),
.B(n_1211),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1298),
.A2(n_900),
.B(n_1147),
.C(n_598),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1225),
.A2(n_1080),
.B(n_1199),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1328),
.B(n_1372),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1369),
.A2(n_1347),
.B(n_1343),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1373),
.B(n_1375),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1311),
.B(n_1302),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1302),
.B(n_1318),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1380),
.B(n_1353),
.Y(n_1386)
);

OAI21xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1330),
.A2(n_1324),
.B(n_1363),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1376),
.A2(n_1313),
.B1(n_1330),
.B2(n_1323),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1347),
.B(n_1326),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1345),
.B(n_1367),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1365),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1360),
.A2(n_1341),
.B(n_1362),
.Y(n_1392)
);

INVxp67_ASAP7_75t_R g1393 ( 
.A(n_1349),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1354),
.B(n_1357),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1352),
.Y(n_1395)
);

AND2x6_ASAP7_75t_SL g1396 ( 
.A(n_1370),
.B(n_1355),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1335),
.B(n_1306),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1348),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1371),
.A2(n_1379),
.B(n_1374),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1333),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1327),
.B(n_1364),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1368),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1314),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1319),
.B(n_1344),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1316),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1329),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1321),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1377),
.Y(n_1408)
);

OAI31xp33_ASAP7_75t_L g1409 ( 
.A1(n_1379),
.A2(n_1315),
.A3(n_1332),
.B(n_1308),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1336),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1331),
.Y(n_1412)
);

NAND2x1_ASAP7_75t_L g1413 ( 
.A(n_1351),
.B(n_1362),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1391),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1409),
.B(n_1312),
.C(n_1320),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1387),
.A2(n_1317),
.B1(n_1304),
.B2(n_1309),
.C(n_1378),
.Y(n_1416)
);

OAI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1409),
.A2(n_1305),
.B1(n_1303),
.B2(n_1346),
.C(n_1358),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1397),
.B(n_1325),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1391),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1391),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_L g1421 ( 
.A(n_1381),
.B(n_1334),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1397),
.B(n_1358),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1401),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1395),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1395),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1400),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1401),
.B(n_1307),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1383),
.B(n_1350),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1394),
.B(n_1359),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1383),
.B(n_1361),
.Y(n_1430)
);

NAND2x1_ASAP7_75t_L g1431 ( 
.A(n_1381),
.B(n_1339),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1381),
.B(n_1340),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1388),
.A2(n_1310),
.B1(n_1340),
.B2(n_1356),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1384),
.B(n_1342),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1388),
.B(n_1322),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1395),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1415),
.B(n_1404),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1431),
.A2(n_1392),
.B(n_1382),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1435),
.A2(n_1387),
.B1(n_1381),
.B2(n_1399),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1424),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1426),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_SL g1442 ( 
.A(n_1432),
.B(n_1389),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1414),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1414),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1428),
.B(n_1418),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1434),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1419),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1428),
.B(n_1393),
.Y(n_1448)
);

NAND4xp25_ASAP7_75t_L g1449 ( 
.A(n_1415),
.B(n_1404),
.C(n_1385),
.D(n_1411),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1433),
.B(n_1322),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1420),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1422),
.A2(n_1385),
.B1(n_1396),
.B2(n_1402),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_1416),
.B(n_1417),
.C(n_1411),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1416),
.B(n_1381),
.C(n_1390),
.Y(n_1454)
);

NOR2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1431),
.B(n_1413),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1434),
.B(n_1384),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1424),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1417),
.A2(n_1381),
.B1(n_1399),
.B2(n_1402),
.Y(n_1459)
);

OAI322xp33_ASAP7_75t_L g1460 ( 
.A1(n_1423),
.A2(n_1412),
.A3(n_1410),
.B1(n_1406),
.B2(n_1408),
.C1(n_1403),
.C2(n_1405),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1427),
.B(n_1407),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1418),
.B(n_1389),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1421),
.B(n_1389),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1418),
.B(n_1389),
.Y(n_1464)
);

OAI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1432),
.A2(n_1381),
.B1(n_1389),
.B2(n_1390),
.C(n_1398),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1423),
.B(n_1429),
.Y(n_1466)
);

NAND4xp25_ASAP7_75t_L g1467 ( 
.A(n_1429),
.B(n_1410),
.C(n_1386),
.D(n_1403),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1432),
.B(n_1390),
.C(n_1389),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1443),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1463),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1441),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1440),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1448),
.B(n_1445),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1443),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1452),
.Y(n_1475)
);

INVx4_ASAP7_75t_SL g1476 ( 
.A(n_1463),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1463),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1452),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1440),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1441),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1437),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1458),
.Y(n_1482)
);

INVx4_ASAP7_75t_SL g1483 ( 
.A(n_1463),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1425),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1449),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1447),
.Y(n_1486)
);

AND4x1_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_1356),
.C(n_1396),
.D(n_1366),
.Y(n_1487)
);

INVx4_ASAP7_75t_SL g1488 ( 
.A(n_1441),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1444),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1466),
.B(n_1436),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1457),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1453),
.B(n_1422),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1451),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1449),
.B(n_1310),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1466),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1469),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1469),
.Y(n_1499)
);

OAI211xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1485),
.A2(n_1439),
.B(n_1459),
.C(n_1454),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1489),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1491),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1481),
.B(n_1430),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1485),
.B(n_1430),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1478),
.B(n_1445),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1476),
.B(n_1448),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1474),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1474),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1467),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

OAI211xp5_ASAP7_75t_L g1511 ( 
.A1(n_1475),
.A2(n_1454),
.B(n_1468),
.C(n_1450),
.Y(n_1511)
);

NOR3xp33_ASAP7_75t_L g1512 ( 
.A(n_1495),
.B(n_1468),
.C(n_1465),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1493),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1472),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1476),
.B(n_1462),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1476),
.B(n_1462),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1476),
.B(n_1464),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1471),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1476),
.B(n_1455),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1496),
.B(n_1467),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1492),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1492),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1494),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1483),
.B(n_1464),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1471),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1484),
.B(n_1446),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1471),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1484),
.B(n_1418),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1461),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1483),
.B(n_1455),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1488),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1490),
.B(n_1422),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1483),
.B(n_1442),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_L g1536 ( 
.A(n_1480),
.B(n_1460),
.C(n_1438),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1470),
.A2(n_1432),
.B1(n_1389),
.B2(n_1399),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1471),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1526),
.B(n_1533),
.Y(n_1539)
);

NAND2x1_ASAP7_75t_L g1540 ( 
.A(n_1520),
.B(n_1491),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1504),
.B(n_1513),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1502),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1507),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1520),
.B(n_1488),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1520),
.B(n_1488),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1507),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1532),
.B(n_1488),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1509),
.B(n_1473),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1508),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1508),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1532),
.B(n_1483),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1510),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1514),
.B(n_1503),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1532),
.B(n_1483),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1526),
.B(n_1480),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1533),
.Y(n_1558)
);

NAND2x1p5_ASAP7_75t_L g1559 ( 
.A(n_1497),
.B(n_1487),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1506),
.B(n_1470),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1510),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1524),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1524),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1499),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1506),
.B(n_1477),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1515),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1505),
.B(n_1480),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1497),
.B(n_1487),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1516),
.B(n_1477),
.Y(n_1571)
);

OAI21xp33_ASAP7_75t_L g1572 ( 
.A1(n_1500),
.A2(n_1390),
.B(n_1479),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1522),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1566),
.B(n_1502),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1541),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1566),
.B(n_1529),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1539),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_1497),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1560),
.B(n_1516),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1560),
.B(n_1517),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1565),
.B(n_1517),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1518),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1545),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1572),
.B(n_1528),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1548),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1539),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1539),
.B(n_1527),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1558),
.B(n_1529),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1550),
.B(n_1531),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1551),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1558),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1552),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1569),
.B(n_1530),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1554),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1542),
.B(n_1527),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1540),
.B(n_1527),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1559),
.B(n_1519),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1574),
.B(n_1555),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1592),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1601)
);

NOR4xp25_ASAP7_75t_L g1602 ( 
.A(n_1587),
.B(n_1543),
.C(n_1568),
.D(n_1567),
.Y(n_1602)
);

OAI32xp33_ASAP7_75t_L g1603 ( 
.A1(n_1597),
.A2(n_1570),
.A3(n_1585),
.B1(n_1592),
.B2(n_1589),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1597),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1581),
.Y(n_1605)
);

OAI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1587),
.A2(n_1570),
.B1(n_1557),
.B2(n_1543),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1590),
.B(n_1571),
.Y(n_1608)
);

OAI31xp33_ASAP7_75t_L g1609 ( 
.A1(n_1585),
.A2(n_1512),
.A3(n_1547),
.B(n_1546),
.Y(n_1609)
);

XNOR2xp5_ASAP7_75t_L g1610 ( 
.A(n_1580),
.B(n_1546),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1547),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1596),
.A2(n_1536),
.B1(n_1537),
.B2(n_1571),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

INVxp33_ASAP7_75t_L g1614 ( 
.A(n_1596),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1578),
.B(n_1564),
.Y(n_1615)
);

OAI31xp33_ASAP7_75t_L g1616 ( 
.A1(n_1598),
.A2(n_1549),
.A3(n_1553),
.B(n_1556),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1598),
.A2(n_1557),
.B(n_1538),
.C(n_1519),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1613),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1605),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1604),
.B(n_1582),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1615),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1608),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1611),
.B(n_1583),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1601),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1594),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1607),
.Y(n_1628)
);

NOR4xp25_ASAP7_75t_L g1629 ( 
.A(n_1627),
.B(n_1619),
.C(n_1626),
.D(n_1620),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1627),
.A2(n_1603),
.B(n_1609),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1618),
.B(n_1625),
.Y(n_1632)
);

AOI211xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1623),
.A2(n_1606),
.B(n_1601),
.C(n_1588),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1624),
.A2(n_1588),
.B(n_1579),
.Y(n_1634)
);

AOI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1621),
.A2(n_1614),
.B(n_1617),
.C(n_1616),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1621),
.B(n_1612),
.C(n_1588),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1622),
.A2(n_1557),
.B1(n_1599),
.B2(n_1519),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1625),
.A2(n_1612),
.B(n_1583),
.Y(n_1638)
);

OAI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1629),
.A2(n_1579),
.B(n_1628),
.Y(n_1639)
);

AOI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1630),
.A2(n_1584),
.B(n_1576),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1632),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1634),
.Y(n_1642)
);

NOR3xp33_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1591),
.C(n_1586),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1642),
.Y(n_1644)
);

AO221x1_ASAP7_75t_L g1645 ( 
.A1(n_1641),
.A2(n_1637),
.B1(n_1633),
.B2(n_1593),
.C(n_1595),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1639),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1643),
.B(n_1635),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1640),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1643),
.B(n_1636),
.C(n_1638),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1644),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1646),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1645),
.B(n_1573),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1647),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1648),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1654),
.B(n_1649),
.C(n_1647),
.D(n_1549),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1651),
.B(n_1653),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_SL g1657 ( 
.A(n_1650),
.B(n_1538),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1656),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1655),
.B1(n_1652),
.B2(n_1657),
.C(n_1653),
.Y(n_1659)
);

OAI211xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1659),
.A2(n_1658),
.B(n_1538),
.C(n_1562),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1659),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1661),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1660),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1658),
.Y(n_1664)
);

XNOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1663),
.B(n_1553),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1665),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1666),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1667),
.A2(n_1664),
.B1(n_1556),
.B2(n_1561),
.C(n_1563),
.Y(n_1668)
);

AO221x2_ASAP7_75t_L g1669 ( 
.A1(n_1668),
.A2(n_1501),
.B1(n_1523),
.B2(n_1534),
.C(n_1482),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1669),
.A2(n_1535),
.B1(n_1471),
.B2(n_1518),
.Y(n_1670)
);

AOI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1535),
.B(n_1501),
.C(n_1525),
.Y(n_1671)
);


endmodule