module fake_ariane_1647_n_372 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_106, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_372);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_106;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_372;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_347;
wire n_183;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_245;
wire n_319;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_117;
wire n_139;
wire n_130;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_327;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_339;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_173;
wire n_242;
wire n_320;
wire n_309;
wire n_115;
wire n_331;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_303;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_333;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_343;
wire n_287;
wire n_302;
wire n_284;
wire n_249;
wire n_212;
wire n_123;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_150;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_118;
wire n_121;
wire n_353;
wire n_241;
wire n_357;
wire n_191;
wire n_211;
wire n_322;
wire n_251;
wire n_116;
wire n_351;
wire n_359;
wire n_155;
wire n_127;

INVx1_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_14),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_49),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_32),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_39),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_29),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_19),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_36),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_47),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_12),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_15),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_28),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_57),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_1),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_62),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_87),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_11),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_4),
.Y(n_155)
);

BUFx2_ASAP7_75t_SL g156 ( 
.A(n_22),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_20),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_30),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_56),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_24),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_21),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_44),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_17),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_25),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_43),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_0),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx11_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_5),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_112),
.B(n_9),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_10),
.B1(n_16),
.B2(n_18),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_118),
.B(n_26),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_27),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_33),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_184),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_154),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_185),
.B1(n_176),
.B2(n_170),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_119),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_186),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_154),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_164),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_111),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_123),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_117),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_135),
.Y(n_218)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_198),
.Y(n_219)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

OR2x6_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_156),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_129),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_214),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_159),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_R g227 ( 
.A(n_190),
.B(n_115),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_120),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_121),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_141),
.Y(n_230)
);

AND2x4_ASAP7_75t_SL g231 ( 
.A(n_200),
.B(n_122),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_144),
.B1(n_163),
.B2(n_147),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_127),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_124),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_125),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_195),
.B(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_126),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_130),
.B1(n_138),
.B2(n_166),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_165),
.C(n_133),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_131),
.B1(n_143),
.B2(n_134),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_196),
.B(n_132),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_SL g246 ( 
.A(n_206),
.B(n_140),
.C(n_142),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_191),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_192),
.B(n_151),
.Y(n_249)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_152),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

OR2x6_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_150),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_219),
.B(n_168),
.Y(n_253)
);

INVx3_ASAP7_75t_SL g254 ( 
.A(n_218),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_139),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_202),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_161),
.B(n_158),
.C(n_148),
.Y(n_257)
);

NAND2x1p5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_162),
.Y(n_260)
);

INVxp33_ASAP7_75t_SL g261 ( 
.A(n_227),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_146),
.B(n_169),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_220),
.A2(n_169),
.B(n_35),
.C(n_37),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_234),
.B(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_34),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_222),
.A2(n_237),
.B(n_244),
.C(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_109),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_38),
.B(n_41),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_233),
.A2(n_42),
.B(n_46),
.C(n_48),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_230),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_250),
.B(n_245),
.Y(n_280)
);

BUFx4_ASAP7_75t_SL g281 ( 
.A(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_232),
.B1(n_241),
.B2(n_243),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_248),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_246),
.B1(n_51),
.B2(n_52),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_50),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_53),
.Y(n_287)
);

AO21x2_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_54),
.B(n_55),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_58),
.B(n_60),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_61),
.B(n_63),
.Y(n_290)
);

OAI211xp5_ASAP7_75t_L g291 ( 
.A1(n_267),
.A2(n_65),
.B(n_67),
.C(n_68),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_255),
.B1(n_251),
.B2(n_273),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_70),
.B(n_71),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_72),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_272),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

AO31x2_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_74),
.A3(n_76),
.B(n_80),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_82),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_282),
.A2(n_258),
.B1(n_260),
.B2(n_252),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_270),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_254),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_256),
.B1(n_271),
.B2(n_257),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_274),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_107),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

OR2x6_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_84),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_86),
.B(n_90),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_286),
.B(n_290),
.Y(n_316)
);

OAI221xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_291),
.B1(n_289),
.B2(n_293),
.C(n_294),
.Y(n_317)
);

AO21x2_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_294),
.B(n_287),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_297),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

CKINVDCx6p67_ASAP7_75t_R g322 ( 
.A(n_311),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_306),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_305),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_311),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_330),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_332),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_321),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_309),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_331),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_333),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_297),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_309),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_309),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_340),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_335),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_336),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_317),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_342),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_351),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

AOI31xp33_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_348),
.A3(n_344),
.B(n_352),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_354),
.B(n_344),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_SL g360 ( 
.A(n_358),
.B(n_341),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_338),
.B1(n_337),
.B2(n_345),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_359),
.B(n_350),
.Y(n_362)
);

AOI221xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_285),
.B1(n_291),
.B2(n_346),
.C(n_347),
.Y(n_363)
);

NOR4xp25_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_303),
.C(n_289),
.D(n_293),
.Y(n_364)
);

NAND4xp75_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_316),
.C(n_280),
.D(n_288),
.Y(n_365)
);

OR3x1_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_364),
.C(n_316),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_366),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_92),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_95),
.B(n_99),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_100),
.B(n_101),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_372)
);


endmodule