module fake_jpeg_8716_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_27),
.B(n_21),
.Y(n_44)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_20),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_19),
.B1(n_16),
.B2(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_35),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_18),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_55),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_34),
.B1(n_39),
.B2(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_63),
.B1(n_65),
.B2(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_39),
.B1(n_31),
.B2(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_33),
.B(n_24),
.C(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_42),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_51),
.C(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_26),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_77),
.B1(n_31),
.B2(n_36),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_37),
.B1(n_36),
.B2(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_19),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_96),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_42),
.B(n_51),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_72),
.B(n_73),
.C(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_28),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_101),
.C(n_59),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_18),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_115),
.C(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_122),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_54),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_117),
.B(n_119),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_62),
.B1(n_57),
.B2(n_71),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_110),
.B1(n_81),
.B2(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_120),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_69),
.B1(n_58),
.B2(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_31),
.B1(n_61),
.B2(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_67),
.B(n_28),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_78),
.C(n_28),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_15),
.B(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_14),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_0),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_1),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_15),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_131),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_91),
.B(n_107),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_125),
.B1(n_98),
.B2(n_122),
.C(n_126),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_101),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_109),
.CON(n_158),
.SN(n_158)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_143),
.Y(n_149)
);

AOI322xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_103),
.A3(n_98),
.B1(n_95),
.B2(n_93),
.C1(n_96),
.C2(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_105),
.B1(n_109),
.B2(n_124),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_117),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_154),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_108),
.B(n_110),
.C(n_119),
.D(n_115),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_108),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_155),
.C(n_158),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_137),
.B(n_130),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_136),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_105),
.A3(n_109),
.B1(n_96),
.B2(n_123),
.C1(n_99),
.C2(n_81),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_170),
.B(n_11),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_136),
.C(n_127),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_174),
.C(n_150),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_137),
.B1(n_130),
.B2(n_132),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_147),
.B1(n_152),
.B2(n_159),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_128),
.B(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_139),
.C(n_146),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_152),
.B(n_149),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_180),
.B1(n_183),
.B2(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_161),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_166),
.C(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_162),
.B1(n_138),
.B2(n_85),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_85),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_184),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_2),
.B(n_3),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_2),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_191),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_172),
.B1(n_166),
.B2(n_164),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_190),
.B(n_192),
.C(n_10),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_172),
.C(n_5),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

AOI31xp67_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_175),
.A3(n_5),
.B(n_6),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

NAND4xp25_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_4),
.C(n_7),
.D(n_9),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_198),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_187),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_197),
.B(n_186),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_7),
.B(n_9),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_188),
.B(n_191),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_10),
.B(n_11),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_10),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_202),
.C(n_203),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_206),
.Y(n_208)
);


endmodule