module fake_jpeg_31977_n_66 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_66);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_66;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx11_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_27),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_11),
.B1(n_19),
.B2(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_3),
.B1(n_7),
.B2(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_27),
.B1(n_23),
.B2(n_16),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_34),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_16),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_40),
.B(n_43),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_25),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_14),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_19),
.B(n_9),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_32),
.B1(n_35),
.B2(n_10),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_43),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_38),
.B1(n_26),
.B2(n_42),
.Y(n_52)
);

XOR2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_20),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_46),
.C(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_32),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_7),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_50),
.B(n_29),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_53),
.B1(n_62),
.B2(n_29),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_3),
.Y(n_66)
);


endmodule