module fake_ariane_1525_n_2560 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2560);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2560;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_1298;
wire n_737;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_762;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_2557;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_907;
wire n_1454;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_476),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_265),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_66),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_232),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_353),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_415),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_216),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_230),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_141),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_510),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_531),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_489),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_256),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_83),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_423),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_277),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_347),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_193),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_368),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_299),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_293),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_530),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_490),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_52),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_255),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_153),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_98),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_103),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_300),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_317),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_193),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_498),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_484),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_361),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_294),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_526),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_500),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_65),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_527),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_379),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_495),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_516),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_432),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_291),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_157),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_239),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_536),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_157),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_502),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_286),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_504),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_56),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_59),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_307),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_361),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_533),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_46),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_480),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_449),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_262),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_431),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_224),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_337),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_70),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_168),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_354),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_329),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_305),
.Y(n_610)
);

CKINVDCx14_ASAP7_75t_R g611 ( 
.A(n_277),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_12),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_299),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_175),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_381),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_243),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_459),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_218),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_175),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_364),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_12),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_144),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_499),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_385),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_141),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_508),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_512),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_49),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_401),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_225),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_483),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_392),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_109),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_457),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_212),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_473),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_242),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_524),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_325),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_136),
.Y(n_640)
);

BUFx8_ASAP7_75t_SL g641 ( 
.A(n_513),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_195),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_199),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_121),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_501),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_255),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_294),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_62),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_511),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_163),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_503),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_197),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_19),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_13),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_212),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_21),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_62),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_318),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_519),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_523),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_446),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_119),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_353),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_292),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_303),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_225),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_262),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_198),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_33),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_170),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_485),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_487),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_22),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_477),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_73),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_329),
.Y(n_677)
);

BUFx5_ASAP7_75t_L g678 ( 
.A(n_129),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_137),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_14),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_186),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_77),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_327),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_196),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_292),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_460),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_514),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_413),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_518),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_172),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_494),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_406),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_537),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_142),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_468),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_346),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_458),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_234),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_13),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_392),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_505),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_174),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_287),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_522),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_472),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_454),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_275),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_385),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_509),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_104),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_61),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_374),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_14),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_481),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_238),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_401),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_520),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_93),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_148),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_171),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_419),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_269),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_259),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_117),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_365),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_440),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_64),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_521),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_365),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_410),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_388),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_247),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_223),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_309),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_529),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_224),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_406),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_515),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_525),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_260),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_309),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_64),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_152),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_209),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_100),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_497),
.Y(n_746)
);

BUFx2_ASAP7_75t_SL g747 ( 
.A(n_507),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_371),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_427),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_52),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_280),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_322),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_301),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_117),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_24),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_534),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_278),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_50),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_68),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_307),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_51),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_199),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_428),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_328),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_517),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_535),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_493),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_553),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_553),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_678),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_569),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_569),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_611),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_653),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_683),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_683),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_678),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_703),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_661),
.B(n_0),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_703),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_743),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_556),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_743),
.Y(n_783)
);

CKINVDCx16_ASAP7_75t_R g784 ( 
.A(n_611),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_678),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_566),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_678),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_678),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_678),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_678),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_551),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_551),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_551),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_551),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_565),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_596),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_596),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_596),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_566),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_596),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_608),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_736),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_687),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_548),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_540),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_556),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_543),
.Y(n_807)
);

CKINVDCx14_ASAP7_75t_R g808 ( 
.A(n_573),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_545),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_608),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_550),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_554),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_608),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_570),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_623),
.B(n_1),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_588),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_608),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_547),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_696),
.B(n_0),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_592),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_687),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_605),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_562),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_606),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_612),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_640),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_618),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_676),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_628),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_640),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_562),
.Y(n_831)
);

INVxp33_ASAP7_75t_SL g832 ( 
.A(n_711),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_571),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_629),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_539),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_647),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_558),
.Y(n_837)
);

INVx4_ASAP7_75t_R g838 ( 
.A(n_641),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_572),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_648),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_574),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_640),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_650),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_641),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_573),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_581),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_561),
.Y(n_847)
);

CKINVDCx16_ASAP7_75t_R g848 ( 
.A(n_541),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_587),
.B(n_1),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_561),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_640),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_603),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_656),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_603),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_696),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_587),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_574),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_681),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_681),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_626),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_658),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_663),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_668),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_669),
.Y(n_864)
);

INVxp33_ASAP7_75t_SL g865 ( 
.A(n_542),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_671),
.Y(n_866)
);

CKINVDCx14_ASAP7_75t_R g867 ( 
.A(n_626),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_681),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_674),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_770),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_803),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_818),
.B(n_595),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_786),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_803),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_803),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_808),
.B(n_768),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_845),
.B(n_583),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_803),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_785),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_770),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_867),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_771),
.B(n_585),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_803),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_844),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_786),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_821),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_838),
.Y(n_887)
);

INVx5_ASAP7_75t_L g888 ( 
.A(n_821),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_818),
.B(n_595),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_777),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_780),
.B(n_586),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_821),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_777),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_837),
.B(n_635),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_837),
.B(n_635),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_821),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_845),
.B(n_589),
.Y(n_897)
);

CKINVDCx16_ASAP7_75t_R g898 ( 
.A(n_784),
.Y(n_898)
);

BUFx8_ASAP7_75t_SL g899 ( 
.A(n_782),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_855),
.B(n_856),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_844),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_796),
.B(n_593),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_839),
.B(n_654),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_799),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_797),
.Y(n_906)
);

INVx5_ASAP7_75t_L g907 ( 
.A(n_821),
.Y(n_907)
);

NOR2x1_ASAP7_75t_L g908 ( 
.A(n_839),
.B(n_747),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_788),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_787),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_787),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_842),
.Y(n_912)
);

BUFx8_ASAP7_75t_SL g913 ( 
.A(n_782),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_846),
.B(n_654),
.Y(n_914)
);

BUFx12f_ASAP7_75t_L g915 ( 
.A(n_799),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_842),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_846),
.B(n_666),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_810),
.B(n_600),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_855),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_789),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_791),
.Y(n_921)
);

XNOR2x2_ASAP7_75t_L g922 ( 
.A(n_806),
.B(n_607),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_790),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_791),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_792),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_792),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_793),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_820),
.Y(n_928)
);

BUFx8_ASAP7_75t_SL g929 ( 
.A(n_806),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_813),
.B(n_666),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_815),
.B(n_568),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_793),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_794),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_817),
.B(n_700),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_826),
.B(n_601),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_919),
.B(n_879),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_887),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_919),
.B(n_849),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_870),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_870),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_919),
.B(n_804),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_928),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_880),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_910),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_916),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_872),
.B(n_856),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_880),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_890),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_879),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_890),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_893),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_893),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_919),
.B(n_849),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_916),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_919),
.B(n_819),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_908),
.B(n_769),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_881),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_911),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_872),
.B(n_772),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_911),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_909),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_916),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_881),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_931),
.B(n_773),
.Y(n_964)
);

CKINVDCx6p67_ASAP7_75t_R g965 ( 
.A(n_915),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_909),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_872),
.B(n_774),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_920),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_931),
.B(n_773),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_900),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_920),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_923),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_923),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_878),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_931),
.B(n_851),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_925),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_925),
.A2(n_645),
.B(n_568),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_927),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_927),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_915),
.B(n_779),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_924),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_924),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_926),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_898),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_926),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_889),
.B(n_775),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_916),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_921),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_878),
.Y(n_989)
);

AND2x2_ASAP7_75t_SL g990 ( 
.A(n_877),
.B(n_645),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_900),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_921),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_884),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_916),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_921),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_889),
.B(n_776),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_889),
.B(n_778),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_897),
.A2(n_832),
.B1(n_865),
.B2(n_833),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_878),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_902),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_931),
.B(n_868),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_887),
.B(n_691),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_931),
.B(n_830),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_876),
.B(n_804),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_921),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_931),
.B(n_833),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_921),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_894),
.B(n_781),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_932),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_932),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_932),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_932),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_878),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_902),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_932),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_933),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_933),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_933),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_933),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_878),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_886),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_930),
.B(n_865),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_910),
.Y(n_1023)
);

INVxp67_ASAP7_75t_R g1024 ( 
.A(n_984),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_961),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_939),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_961),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_968),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_968),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_972),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_990),
.B(n_910),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_938),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_990),
.B(n_910),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_949),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_945),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_990),
.B(n_910),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_938),
.B(n_882),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_1006),
.B(n_891),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_939),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_973),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_943),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_943),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_947),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_973),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_938),
.B(n_930),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_945),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_947),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_949),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_976),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_958),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_L g1051 ( 
.A(n_966),
.B(n_873),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_938),
.B(n_930),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1004),
.B(n_847),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_953),
.B(n_934),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_944),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_949),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_976),
.Y(n_1057)
);

AND3x2_ASAP7_75t_L g1058 ( 
.A(n_1002),
.B(n_905),
.C(n_885),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1022),
.A2(n_756),
.B1(n_691),
.B2(n_832),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_953),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_949),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_978),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_953),
.A2(n_756),
.B1(n_828),
.B2(n_795),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_953),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_958),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_985),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_985),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_964),
.B(n_651),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_978),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_979),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_985),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_940),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_940),
.Y(n_1073)
);

AND2x6_ASAP7_75t_L g1074 ( 
.A(n_955),
.B(n_894),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_945),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_979),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_1015),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_1015),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_966),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_971),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_942),
.B(n_847),
.Y(n_1081)
);

NAND2xp33_ASAP7_75t_SL g1082 ( 
.A(n_957),
.B(n_758),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_969),
.A2(n_934),
.B1(n_918),
.B2(n_903),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_971),
.B(n_659),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_998),
.B(n_850),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_981),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_942),
.B(n_850),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_993),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_948),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_1015),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_1015),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_948),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_981),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_SL g1094 ( 
.A(n_965),
.B(n_887),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1015),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_950),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1000),
.B(n_852),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_950),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_951),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1014),
.B(n_852),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_951),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_955),
.B(n_1015),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_952),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_952),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_944),
.Y(n_1105)
);

NAND2xp33_ASAP7_75t_SL g1106 ( 
.A(n_957),
.B(n_584),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_960),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_960),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_982),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_955),
.B(n_660),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_982),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_983),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_983),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_988),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_997),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_997),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_945),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_988),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_945),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_955),
.B(n_675),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1007),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_936),
.B(n_686),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1008),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1008),
.Y(n_1125)
);

NOR2x1p5_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_854),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_970),
.B(n_854),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_970),
.B(n_894),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_967),
.B(n_848),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_991),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_L g1131 ( 
.A(n_945),
.B(n_681),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_991),
.B(n_835),
.C(n_860),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_975),
.B(n_689),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1001),
.B(n_705),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_974),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_959),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1007),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1003),
.B(n_735),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1011),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_941),
.B(n_860),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_954),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1011),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_895),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_956),
.B(n_746),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_956),
.B(n_934),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_956),
.B(n_765),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1012),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1012),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_956),
.B(n_904),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_959),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1016),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_SL g1152 ( 
.A(n_980),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1019),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_974),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1019),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_992),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_992),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_946),
.B(n_802),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1049),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1057),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1062),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1066),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1069),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1070),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1032),
.B(n_963),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1076),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1025),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1027),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1028),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1082),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1159),
.B(n_946),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1130),
.B(n_959),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1029),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1030),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1088),
.Y(n_1176)
);

INVxp33_ASAP7_75t_L g1177 ( 
.A(n_1081),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1087),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1129),
.B(n_1053),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1127),
.B(n_959),
.Y(n_1180)
);

XOR2x2_ASAP7_75t_L g1181 ( 
.A(n_1085),
.B(n_922),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1040),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1037),
.B(n_986),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1079),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1116),
.B(n_986),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1149),
.B(n_1136),
.Y(n_1187)
);

INVxp33_ASAP7_75t_L g1188 ( 
.A(n_1097),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1080),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1072),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1038),
.A2(n_1005),
.B(n_995),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1072),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1073),
.Y(n_1193)
);

XOR2x2_ASAP7_75t_L g1194 ( 
.A(n_1059),
.B(n_922),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1073),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1032),
.B(n_986),
.Y(n_1196)
);

XOR2xp5_ASAP7_75t_L g1197 ( 
.A(n_1132),
.B(n_937),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1089),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1066),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1089),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1092),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1128),
.B(n_986),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1092),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1117),
.B(n_996),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1149),
.B(n_996),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1098),
.Y(n_1206)
);

CKINVDCx16_ASAP7_75t_R g1207 ( 
.A(n_1094),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1124),
.B(n_996),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1099),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1099),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1103),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1125),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1103),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1108),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1035),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1031),
.A2(n_1005),
.B(n_995),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1031),
.A2(n_1010),
.B(n_1009),
.Y(n_1217)
);

XNOR2xp5_ASAP7_75t_L g1218 ( 
.A(n_1126),
.B(n_823),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1067),
.Y(n_1219)
);

NOR2x1_ASAP7_75t_L g1220 ( 
.A(n_1051),
.B(n_980),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_L g1221 ( 
.A(n_1100),
.B(n_996),
.Y(n_1221)
);

INVxp33_ASAP7_75t_L g1222 ( 
.A(n_1128),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1108),
.Y(n_1223)
);

XOR2xp5_ASAP7_75t_L g1224 ( 
.A(n_1063),
.B(n_823),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1067),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1149),
.B(n_980),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1086),
.B(n_1009),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1060),
.B(n_584),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1096),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1060),
.B(n_980),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1101),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1093),
.B(n_1010),
.Y(n_1232)
);

CKINVDCx16_ASAP7_75t_R g1233 ( 
.A(n_1082),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1104),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1109),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1150),
.Y(n_1236)
);

INVxp33_ASAP7_75t_L g1237 ( 
.A(n_1143),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1038),
.A2(n_1018),
.B(n_1017),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1157),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1158),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1106),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1058),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1140),
.B(n_980),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1074),
.B(n_1017),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1158),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1110),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1112),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1143),
.B(n_895),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1071),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1113),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1026),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1026),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1064),
.B(n_895),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1024),
.B(n_904),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1039),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1064),
.B(n_1018),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1114),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1039),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1041),
.Y(n_1259)
);

INVxp67_ASAP7_75t_SL g1260 ( 
.A(n_1045),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1052),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1145),
.B(n_935),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1042),
.Y(n_1263)
);

INVxp33_ASAP7_75t_L g1264 ( 
.A(n_1144),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1042),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1043),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1051),
.B(n_904),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1043),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1047),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_1054),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1144),
.B(n_1146),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1146),
.B(n_831),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1050),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1050),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1065),
.Y(n_1275)
);

AND2x6_ASAP7_75t_L g1276 ( 
.A(n_1048),
.B(n_954),
.Y(n_1276)
);

INVxp33_ASAP7_75t_L g1277 ( 
.A(n_1111),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1074),
.B(n_1102),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1065),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1035),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1033),
.B(n_974),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1111),
.B(n_914),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1115),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1106),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1115),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1119),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1033),
.B(n_989),
.Y(n_1287)
);

BUFx8_ASAP7_75t_L g1288 ( 
.A(n_1152),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1074),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1074),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1119),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1036),
.A2(n_977),
.B(n_989),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1121),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1122),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1122),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_1121),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1036),
.B(n_1048),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1152),
.B(n_622),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1137),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1152),
.Y(n_1300)
);

XOR2xp5_ASAP7_75t_L g1301 ( 
.A(n_1083),
.B(n_831),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1137),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_1035),
.B(n_954),
.Y(n_1303)
);

XOR2xp5_ASAP7_75t_L g1304 ( 
.A(n_1133),
.B(n_841),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1139),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1084),
.B(n_914),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1139),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1074),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1074),
.B(n_989),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1142),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1142),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1084),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1048),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1147),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1147),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1148),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1148),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1102),
.Y(n_1318)
);

INVxp33_ASAP7_75t_L g1319 ( 
.A(n_1123),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1133),
.B(n_914),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1151),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1151),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1153),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1035),
.Y(n_1324)
);

XOR2xp5_ASAP7_75t_L g1325 ( 
.A(n_1134),
.B(n_841),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1153),
.Y(n_1326)
);

XOR2xp5_ASAP7_75t_L g1327 ( 
.A(n_1134),
.B(n_857),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1154),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1154),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_SL g1330 ( 
.A(n_1078),
.B(n_622),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1156),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1107),
.Y(n_1332)
);

XOR2xp5_ASAP7_75t_L g1333 ( 
.A(n_1138),
.B(n_857),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1107),
.Y(n_1334)
);

AND2x2_ASAP7_75t_SL g1335 ( 
.A(n_1078),
.B(n_899),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1107),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1056),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1056),
.B(n_989),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1056),
.Y(n_1339)
);

XNOR2x2_ASAP7_75t_L g1340 ( 
.A(n_1138),
.B(n_899),
.Y(n_1340)
);

XOR2x2_ASAP7_75t_L g1341 ( 
.A(n_1068),
.B(n_913),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1135),
.B(n_917),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1061),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1061),
.B(n_999),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1135),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1135),
.B(n_917),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1078),
.B(n_962),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1061),
.B(n_999),
.Y(n_1348)
);

INVxp33_ASAP7_75t_SL g1349 ( 
.A(n_1123),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1034),
.B(n_999),
.Y(n_1350)
);

XNOR2xp5_ASAP7_75t_L g1351 ( 
.A(n_1068),
.B(n_913),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1155),
.B(n_917),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1090),
.B(n_1034),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1251),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1188),
.B(n_1034),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1179),
.B(n_1172),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1330),
.A2(n_619),
.B1(n_620),
.B2(n_590),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1176),
.B(n_929),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1160),
.Y(n_1359)
);

NOR3xp33_ASAP7_75t_L g1360 ( 
.A(n_1243),
.B(n_688),
.C(n_677),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1252),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1330),
.A2(n_619),
.B1(n_620),
.B2(n_590),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1262),
.B(n_1155),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1255),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1288),
.Y(n_1365)
);

NOR2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1178),
.B(n_929),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1243),
.A2(n_1155),
.B(n_1091),
.C(n_1095),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1221),
.B(n_1046),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1215),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1262),
.B(n_1077),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1177),
.B(n_707),
.Y(n_1371)
);

INVxp33_ASAP7_75t_L g1372 ( 
.A(n_1304),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1226),
.B(n_1090),
.Y(n_1373)
);

AOI22x1_ASAP7_75t_L g1374 ( 
.A1(n_1313),
.A2(n_1090),
.B1(n_1091),
.B2(n_1077),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1161),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1181),
.A2(n_719),
.B1(n_748),
.B2(n_707),
.Y(n_1376)
);

AO221x1_ASAP7_75t_L g1377 ( 
.A1(n_1284),
.A2(n_715),
.B1(n_684),
.B2(n_1075),
.C(n_1046),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1237),
.B(n_1349),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1180),
.B(n_1077),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_L g1380 ( 
.A(n_1276),
.B(n_1118),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1183),
.B(n_1091),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1288),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1254),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1272),
.B(n_783),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1162),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1202),
.B(n_1248),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1173),
.B(n_1075),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1186),
.B(n_1095),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1233),
.B(n_719),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1186),
.B(n_1095),
.Y(n_1390)
);

BUFx5_ASAP7_75t_L g1391 ( 
.A(n_1276),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1164),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1205),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1222),
.B(n_1075),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1264),
.B(n_1075),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1204),
.B(n_1118),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1212),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1204),
.B(n_1118),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1194),
.B(n_1205),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1300),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1166),
.B(n_698),
.C(n_690),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1301),
.A2(n_1278),
.B1(n_1228),
.B2(n_1226),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1224),
.A2(n_541),
.B1(n_602),
.B2(n_594),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1260),
.B(n_1120),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1260),
.B(n_1261),
.Y(n_1405)
);

NAND2xp33_ASAP7_75t_L g1406 ( 
.A(n_1276),
.B(n_1120),
.Y(n_1406)
);

INVxp33_ASAP7_75t_L g1407 ( 
.A(n_1325),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1187),
.B(n_1120),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1208),
.B(n_1120),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1241),
.B(n_541),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1187),
.B(n_1278),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1208),
.B(n_1141),
.Y(n_1412)
);

OR2x6_ASAP7_75t_L g1413 ( 
.A(n_1308),
.B(n_805),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1239),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1271),
.B(n_609),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1271),
.B(n_644),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1240),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1261),
.B(n_1055),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1165),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1303),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1270),
.B(n_1190),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1207),
.Y(n_1422)
);

O2A1O1Ixp5_ASAP7_75t_L g1423 ( 
.A1(n_1281),
.A2(n_999),
.B(n_1020),
.C(n_1013),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1215),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1245),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1163),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1345),
.B(n_1055),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1335),
.B(n_1055),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1298),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1270),
.B(n_652),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1267),
.B(n_1167),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1192),
.B(n_1055),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1277),
.B(n_664),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1276),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1168),
.B(n_692),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1174),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1199),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1219),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1318),
.A2(n_721),
.B1(n_731),
.B2(n_694),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1230),
.B(n_1055),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1175),
.Y(n_1442)
);

INVx8_ASAP7_75t_L g1443 ( 
.A(n_1253),
.Y(n_1443)
);

XOR2xp5_ASAP7_75t_L g1444 ( 
.A(n_1218),
.B(n_807),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1340),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1296),
.B(n_1013),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1182),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1298),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1293),
.B(n_594),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1184),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1229),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1225),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1231),
.Y(n_1453)
);

OR2x2_ASAP7_75t_SL g1454 ( 
.A(n_1341),
.B(n_700),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1242),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1327),
.B(n_594),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1230),
.B(n_1105),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1289),
.B(n_1105),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1234),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1289),
.B(n_1105),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1333),
.A2(n_657),
.B1(n_602),
.B2(n_544),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1249),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1235),
.A2(n_713),
.B1(n_729),
.B2(n_720),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1220),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1290),
.B(n_1105),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1193),
.B(n_1105),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1195),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1290),
.B(n_954),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_L g1469 ( 
.A(n_1313),
.B(n_954),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1198),
.B(n_1013),
.Y(n_1470)
);

INVx8_ASAP7_75t_L g1471 ( 
.A(n_1253),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1319),
.B(n_1013),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1351),
.B(n_809),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1200),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1185),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1171),
.B(n_602),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1206),
.B(n_1020),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1189),
.Y(n_1479)
);

AND2x2_ASAP7_75t_SL g1480 ( 
.A(n_1282),
.B(n_1131),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1320),
.A2(n_657),
.B1(n_546),
.B2(n_555),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1209),
.B(n_1020),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1197),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1280),
.B(n_962),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1280),
.B(n_962),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_SL g1486 ( 
.A(n_1253),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1246),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1236),
.B(n_1020),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1297),
.A2(n_1021),
.B(n_749),
.C(n_627),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1306),
.B(n_811),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1196),
.A2(n_557),
.B1(n_559),
.B2(n_552),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1342),
.B(n_812),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1312),
.B(n_1244),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1210),
.B(n_1021),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1247),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1211),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1297),
.A2(n_564),
.B1(n_567),
.B2(n_563),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1337),
.B(n_1021),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1346),
.B(n_657),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1352),
.B(n_814),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1227),
.A2(n_741),
.B1(n_744),
.B2(n_734),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1250),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1213),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1257),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1214),
.B(n_1021),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1223),
.B(n_816),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1339),
.B(n_962),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1343),
.B(n_962),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1324),
.B(n_987),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1332),
.B(n_575),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1258),
.B(n_987),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_SL g1512 ( 
.A(n_1324),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1259),
.A2(n_580),
.B1(n_597),
.B2(n_578),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1334),
.B(n_599),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1227),
.B(n_1232),
.Y(n_1515)
);

NOR2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1244),
.B(n_822),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1309),
.B(n_987),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1263),
.B(n_824),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1353),
.Y(n_1519)
);

NOR2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1309),
.B(n_825),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1265),
.B(n_827),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1256),
.B(n_987),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1232),
.B(n_829),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1266),
.B(n_834),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1256),
.B(n_987),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1268),
.B(n_994),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1269),
.B(n_836),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1273),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1274),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1275),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1279),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1283),
.B(n_840),
.Y(n_1532)
);

AND2x6_ASAP7_75t_SL g1533 ( 
.A(n_1281),
.B(n_843),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1336),
.B(n_994),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1285),
.B(n_994),
.Y(n_1535)
);

NAND2x1_ASAP7_75t_L g1536 ( 
.A(n_1353),
.B(n_994),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1353),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1347),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1286),
.B(n_1316),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1291),
.B(n_994),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_L g1541 ( 
.A(n_1350),
.B(n_994),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1287),
.B(n_604),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1294),
.B(n_944),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1287),
.B(n_610),
.Y(n_1544)
);

NAND2x1_ASAP7_75t_L g1545 ( 
.A(n_1295),
.B(n_944),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1299),
.A2(n_614),
.B1(n_615),
.B2(n_613),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1302),
.B(n_1023),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1305),
.B(n_853),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1356),
.B(n_616),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1384),
.B(n_1307),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1541),
.A2(n_1350),
.B(n_1344),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1430),
.B(n_1310),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1415),
.B(n_1311),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_SL g1554 ( 
.A1(n_1363),
.A2(n_1344),
.B(n_1338),
.C(n_1348),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1542),
.A2(n_1217),
.B(n_1216),
.C(n_1292),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1380),
.A2(n_1348),
.B(n_1338),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1389),
.B(n_861),
.Y(n_1557)
);

NOR3xp33_ASAP7_75t_L g1558 ( 
.A(n_1501),
.B(n_755),
.C(n_753),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1414),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1416),
.B(n_1314),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1370),
.A2(n_1217),
.B(n_1216),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1357),
.B(n_1315),
.Y(n_1562)
);

BUFx4f_ASAP7_75t_L g1563 ( 
.A(n_1537),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1417),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1360),
.A2(n_639),
.B1(n_667),
.B2(n_630),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1405),
.B(n_1317),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1359),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1406),
.A2(n_1131),
.B(n_1321),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1469),
.A2(n_1515),
.B(n_1405),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1370),
.A2(n_1238),
.B(n_1191),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1425),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1378),
.B(n_1322),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1395),
.B(n_1431),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1537),
.B(n_1323),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1393),
.B(n_1326),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1499),
.B(n_1328),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1473),
.B(n_621),
.Y(n_1577)
);

AOI33xp33_ASAP7_75t_L g1578 ( 
.A1(n_1461),
.A2(n_760),
.A3(n_754),
.B1(n_759),
.B2(n_752),
.B3(n_862),
.Y(n_1578)
);

NOR3xp33_ASAP7_75t_L g1579 ( 
.A(n_1501),
.B(n_864),
.C(n_863),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1433),
.B(n_1329),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1397),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1537),
.B(n_1394),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1393),
.B(n_1490),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1519),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1376),
.A2(n_1331),
.B1(n_869),
.B2(n_866),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1420),
.A2(n_977),
.B(n_1023),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1544),
.A2(n_798),
.B(n_800),
.C(n_794),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1467),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1520),
.A2(n_906),
.B(n_901),
.C(n_625),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1363),
.A2(n_977),
.B(n_1023),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_R g1591 ( 
.A(n_1422),
.B(n_901),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1399),
.B(n_1476),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1375),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1418),
.A2(n_977),
.B(n_1023),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_L g1595 ( 
.A(n_1382),
.B(n_901),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1362),
.A2(n_680),
.B1(n_699),
.B2(n_633),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1373),
.B(n_906),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1418),
.A2(n_800),
.B(n_798),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1369),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1434),
.A2(n_1404),
.B(n_1381),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1383),
.B(n_624),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1373),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1434),
.A2(n_1404),
.B(n_1412),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1367),
.A2(n_858),
.B(n_801),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1423),
.A2(n_637),
.B(n_632),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1396),
.B(n_933),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1523),
.B(n_642),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1366),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1373),
.B(n_906),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1436),
.B(n_643),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1372),
.B(n_646),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_SL g1612 ( 
.A1(n_1388),
.A2(n_859),
.B(n_4),
.C(n_2),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1385),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1398),
.A2(n_665),
.B(n_655),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1386),
.A2(n_679),
.B1(n_682),
.B2(n_670),
.Y(n_1615)
);

AO21x1_ASAP7_75t_L g1616 ( 
.A1(n_1421),
.A2(n_859),
.B(n_715),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1409),
.B(n_538),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1371),
.B(n_685),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1392),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1419),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1410),
.B(n_702),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1379),
.B(n_549),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1518),
.B(n_708),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1527),
.B(n_710),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1390),
.A2(n_716),
.B(n_712),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1510),
.A2(n_722),
.B(n_718),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1374),
.A2(n_714),
.B(n_687),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1489),
.A2(n_724),
.B(n_725),
.C(n_723),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1548),
.B(n_727),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1492),
.B(n_730),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1369),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1500),
.B(n_732),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1432),
.A2(n_714),
.B(n_687),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1514),
.A2(n_737),
.B(n_733),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1432),
.A2(n_767),
.B(n_714),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1516),
.A2(n_742),
.B(n_745),
.C(n_740),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1449),
.B(n_750),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1477),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1474),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1407),
.B(n_751),
.Y(n_1640)
);

O2A1O1Ixp33_ASAP7_75t_SL g1641 ( 
.A1(n_1355),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1533),
.B(n_757),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1466),
.A2(n_767),
.B(n_714),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1497),
.A2(n_761),
.B1(n_764),
.B2(n_762),
.Y(n_1644)
);

NOR2x1p5_ASAP7_75t_L g1645 ( 
.A(n_1445),
.B(n_684),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1466),
.A2(n_1525),
.B(n_1522),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1437),
.B(n_684),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1481),
.A2(n_715),
.B1(n_684),
.B2(n_560),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1411),
.B(n_1519),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1442),
.B(n_3),
.Y(n_1650)
);

NOR2x1_ASAP7_75t_L g1651 ( 
.A(n_1428),
.B(n_767),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1447),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1496),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1369),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1536),
.A2(n_912),
.B(n_892),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1480),
.B(n_1402),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1503),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1450),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1451),
.B(n_5),
.Y(n_1659)
);

NOR2xp67_ASAP7_75t_L g1660 ( 
.A(n_1464),
.B(n_429),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1488),
.A2(n_577),
.B1(n_579),
.B2(n_576),
.Y(n_1661)
);

O2A1O1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1463),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1358),
.B(n_582),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1453),
.B(n_6),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1424),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1491),
.A2(n_739),
.B(n_738),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1459),
.B(n_7),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1401),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1484),
.A2(n_1509),
.B(n_1485),
.Y(n_1669)
);

OR2x6_ASAP7_75t_L g1670 ( 
.A(n_1443),
.B(n_886),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1456),
.B(n_10),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1472),
.A2(n_598),
.B(n_617),
.C(n_591),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1429),
.B(n_11),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1424),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1529),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1448),
.B(n_11),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1424),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1455),
.Y(n_1678)
);

BUFx12f_ASAP7_75t_L g1679 ( 
.A(n_1365),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1435),
.B(n_15),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1377),
.A2(n_634),
.B(n_631),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1440),
.A2(n_638),
.B1(n_649),
.B2(n_636),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1538),
.B(n_763),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1446),
.A2(n_672),
.B(n_673),
.C(n_662),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1517),
.A2(n_695),
.B(n_693),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1483),
.B(n_697),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1512),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1475),
.B(n_1479),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1507),
.A2(n_704),
.B(n_701),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1507),
.A2(n_709),
.B(n_706),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1400),
.B(n_717),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1508),
.A2(n_728),
.B(n_726),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1487),
.B(n_15),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1387),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1495),
.B(n_16),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1413),
.B(n_912),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1477),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1444),
.B(n_766),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1538),
.B(n_912),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1508),
.A2(n_892),
.B(n_886),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1513),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1701)
);

CKINVDCx8_ASAP7_75t_R g1702 ( 
.A(n_1443),
.Y(n_1702)
);

AND2x2_ASAP7_75t_SL g1703 ( 
.A(n_1403),
.B(n_20),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1512),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1493),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1502),
.B(n_20),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1511),
.A2(n_892),
.B(n_886),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1470),
.A2(n_874),
.B(n_871),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1511),
.A2(n_892),
.B(n_886),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1526),
.A2(n_892),
.B(n_874),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1526),
.A2(n_874),
.B(n_871),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1408),
.B(n_21),
.C(n_22),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1506),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1443),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1471),
.B(n_23),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1454),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1470),
.A2(n_874),
.B(n_871),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1486),
.B(n_25),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1535),
.A2(n_874),
.B(n_871),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1538),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1530),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1535),
.A2(n_875),
.B(n_871),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1391),
.B(n_912),
.Y(n_1723)
);

AND3x1_ASAP7_75t_L g1724 ( 
.A(n_1546),
.B(n_26),
.C(n_27),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1413),
.B(n_912),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1540),
.A2(n_883),
.B(n_875),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1540),
.A2(n_883),
.B(n_875),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1478),
.A2(n_883),
.B(n_875),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1441),
.A2(n_883),
.B(n_875),
.Y(n_1729)
);

OAI21xp33_ASAP7_75t_L g1730 ( 
.A1(n_1498),
.A2(n_26),
.B(n_27),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1471),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1457),
.A2(n_888),
.B(n_883),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1504),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1413),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1471),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1493),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1703),
.A2(n_1486),
.B1(n_1493),
.B2(n_1368),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1583),
.B(n_1521),
.Y(n_1738)
);

OR2x6_ASAP7_75t_SL g1739 ( 
.A(n_1642),
.B(n_1524),
.Y(n_1739)
);

OAI321xp33_ASAP7_75t_L g1740 ( 
.A1(n_1730),
.A2(n_1532),
.A3(n_1539),
.B1(n_1528),
.B2(n_1482),
.C(n_1494),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1608),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1569),
.A2(n_1427),
.B(n_1478),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1688),
.Y(n_1743)
);

AO21x2_ASAP7_75t_L g1744 ( 
.A1(n_1616),
.A2(n_1539),
.B(n_1468),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1577),
.A2(n_1458),
.B1(n_1460),
.B2(n_1465),
.Y(n_1745)
);

AOI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1627),
.A2(n_1534),
.B(n_1505),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1556),
.A2(n_1494),
.B(n_1482),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1565),
.A2(n_1543),
.B1(n_1547),
.B2(n_1531),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1702),
.B(n_1426),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1626),
.A2(n_1634),
.B(n_1680),
.C(n_1662),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1550),
.B(n_1438),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1551),
.A2(n_1547),
.B(n_1543),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1663),
.B(n_28),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1592),
.A2(n_1361),
.B1(n_1364),
.B2(n_1354),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1559),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1572),
.B(n_1439),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1696),
.B(n_1391),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1563),
.B(n_1452),
.Y(n_1758)
);

O2A1O1Ixp33_ASAP7_75t_SL g1759 ( 
.A1(n_1555),
.A2(n_1545),
.B(n_1391),
.C(n_1462),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1696),
.B(n_1391),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1628),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1714),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1599),
.Y(n_1763)
);

NAND2x1p5_ASAP7_75t_L g1764 ( 
.A(n_1563),
.B(n_888),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1557),
.B(n_1638),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_R g1766 ( 
.A(n_1679),
.B(n_888),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1565),
.A2(n_1724),
.B1(n_1596),
.B2(n_1625),
.Y(n_1767)
);

AO21x2_ASAP7_75t_L g1768 ( 
.A1(n_1570),
.A2(n_896),
.B(n_888),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1558),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.C(n_34),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1725),
.B(n_888),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1697),
.B(n_32),
.Y(n_1771)
);

BUFx4f_ASAP7_75t_SL g1772 ( 
.A(n_1581),
.Y(n_1772)
);

OR2x6_ASAP7_75t_L g1773 ( 
.A(n_1715),
.B(n_430),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1564),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1580),
.B(n_1553),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1698),
.A2(n_907),
.B1(n_896),
.B2(n_36),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_L g1777 ( 
.A(n_1714),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1591),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1567),
.Y(n_1779)
);

NOR2x1p5_ASAP7_75t_SL g1780 ( 
.A(n_1593),
.B(n_1613),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1668),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1714),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1596),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1649),
.B(n_37),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1686),
.B(n_38),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1701),
.A2(n_1734),
.B(n_1644),
.C(n_1713),
.Y(n_1786)
);

OAI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1712),
.A2(n_39),
.B(n_40),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1600),
.A2(n_907),
.B(n_896),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1603),
.A2(n_907),
.B(n_896),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1607),
.A2(n_907),
.B(n_896),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1554),
.A2(n_907),
.B(n_39),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1571),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1578),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1735),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1611),
.B(n_41),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1619),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1671),
.B(n_42),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1687),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1568),
.A2(n_43),
.B(n_44),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1588),
.Y(n_1800)
);

AO22x1_ASAP7_75t_L g1801 ( 
.A1(n_1718),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1708),
.A2(n_1728),
.B(n_1717),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1560),
.B(n_45),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1618),
.B(n_46),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1614),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1552),
.B(n_47),
.Y(n_1806)
);

AOI22x1_ASAP7_75t_L g1807 ( 
.A1(n_1689),
.A2(n_1690),
.B1(n_1692),
.B2(n_1605),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1561),
.A2(n_48),
.B(n_50),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1715),
.A2(n_1549),
.B1(n_1621),
.B2(n_1636),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1599),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1707),
.A2(n_51),
.B(n_53),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1637),
.B(n_53),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1656),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_1813)
);

O2A1O1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1682),
.A2(n_57),
.B(n_54),
.C(n_55),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1639),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1709),
.A2(n_57),
.B(n_58),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1715),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1666),
.A2(n_63),
.B(n_60),
.C(n_61),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1610),
.A2(n_66),
.B1(n_63),
.B2(n_65),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1612),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1820)
);

OAI21xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1650),
.A2(n_1664),
.B(n_1659),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1725),
.B(n_67),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1672),
.A2(n_69),
.B(n_70),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1700),
.A2(n_71),
.B(n_72),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1630),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1825)
);

AOI22x1_ASAP7_75t_L g1826 ( 
.A1(n_1646),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1590),
.A2(n_74),
.B(n_75),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1615),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1673),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1620),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1652),
.B(n_79),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1594),
.A2(n_80),
.B(n_81),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1584),
.B(n_81),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1632),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1584),
.B(n_1599),
.Y(n_1835)
);

AOI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1681),
.A2(n_434),
.B(n_433),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1658),
.B(n_82),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1586),
.A2(n_84),
.B(n_85),
.Y(n_1838)
);

INVx5_ASAP7_75t_L g1839 ( 
.A(n_1670),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1676),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1566),
.A2(n_86),
.B(n_87),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1669),
.A2(n_1723),
.B(n_1635),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1684),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1633),
.A2(n_88),
.B(n_89),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1640),
.B(n_90),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1694),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1643),
.A2(n_91),
.B(n_92),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1733),
.B(n_94),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1710),
.A2(n_94),
.B(n_95),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1653),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1576),
.B(n_95),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1606),
.A2(n_96),
.B(n_97),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1573),
.B(n_96),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1661),
.A2(n_97),
.B(n_98),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1716),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1704),
.Y(n_1856)
);

BUFx8_ASAP7_75t_L g1857 ( 
.A(n_1631),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1631),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1657),
.B(n_99),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1691),
.B(n_101),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1711),
.A2(n_102),
.B(n_103),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1675),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1649),
.B(n_435),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1631),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1719),
.A2(n_102),
.B(n_104),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1623),
.B(n_105),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1721),
.B(n_105),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1585),
.B(n_106),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1678),
.B(n_106),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1602),
.B(n_107),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1562),
.B(n_107),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1595),
.B(n_108),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1654),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1575),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1687),
.B(n_108),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1722),
.A2(n_109),
.B(n_110),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1575),
.B(n_110),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1731),
.B(n_111),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1654),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1726),
.A2(n_111),
.B(n_112),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1667),
.A2(n_1693),
.B1(n_1706),
.B2(n_1695),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1727),
.A2(n_112),
.B(n_113),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1654),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1617),
.A2(n_113),
.B(n_114),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1645),
.B(n_114),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1589),
.A2(n_118),
.B1(n_115),
.B2(n_116),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1624),
.B(n_115),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1674),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1629),
.B(n_116),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1720),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1647),
.Y(n_1891)
);

OAI21xp33_ASAP7_75t_L g1892 ( 
.A1(n_1579),
.A2(n_118),
.B(n_119),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1655),
.A2(n_120),
.B(n_121),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1641),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1731),
.B(n_122),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1705),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1597),
.B(n_123),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1842),
.A2(n_1604),
.B(n_1598),
.Y(n_1898)
);

CKINVDCx20_ASAP7_75t_R g1899 ( 
.A(n_1772),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1747),
.A2(n_1651),
.B(n_1736),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1765),
.B(n_1720),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1857),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1775),
.B(n_1665),
.Y(n_1903)
);

OAI21xp33_ASAP7_75t_L g1904 ( 
.A1(n_1753),
.A2(n_1648),
.B(n_1601),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1802),
.A2(n_1670),
.B(n_1685),
.Y(n_1905)
);

NAND3x1_ASAP7_75t_L g1906 ( 
.A(n_1795),
.B(n_1736),
.C(n_1677),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1779),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1743),
.B(n_1665),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1857),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1759),
.A2(n_1670),
.B(n_1699),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1821),
.B(n_1881),
.Y(n_1911)
);

INVx8_ASAP7_75t_L g1912 ( 
.A(n_1773),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1752),
.A2(n_1732),
.B(n_1729),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1741),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1785),
.B(n_1683),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1742),
.A2(n_1838),
.B(n_1832),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1796),
.B(n_1582),
.Y(n_1917)
);

BUFx8_ASAP7_75t_L g1918 ( 
.A(n_1812),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1804),
.B(n_1677),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1762),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1762),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1738),
.B(n_1674),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1746),
.A2(n_1574),
.B(n_1587),
.Y(n_1923)
);

AO31x2_ASAP7_75t_L g1924 ( 
.A1(n_1748),
.A2(n_1660),
.A3(n_1622),
.B(n_1674),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1827),
.A2(n_1609),
.B(n_1597),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1830),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1756),
.B(n_1751),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1896),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1771),
.B(n_1609),
.Y(n_1929)
);

A2O1A1Ixp33_ASAP7_75t_L g1930 ( 
.A1(n_1750),
.A2(n_1860),
.B(n_1767),
.C(n_1845),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1780),
.B(n_436),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1808),
.A2(n_124),
.B(n_125),
.Y(n_1932)
);

OAI21x1_ASAP7_75t_L g1933 ( 
.A1(n_1791),
.A2(n_438),
.B(n_437),
.Y(n_1933)
);

OAI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1823),
.A2(n_124),
.B(n_125),
.Y(n_1934)
);

NAND2xp33_ASAP7_75t_L g1935 ( 
.A(n_1787),
.B(n_126),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1790),
.A2(n_1740),
.B(n_1799),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1794),
.B(n_126),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1858),
.B(n_442),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1806),
.B(n_127),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1858),
.Y(n_1940)
);

AOI21x1_ASAP7_75t_SL g1941 ( 
.A1(n_1895),
.A2(n_1853),
.B(n_1878),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1762),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1778),
.B(n_127),
.Y(n_1943)
);

AO31x2_ASAP7_75t_L g1944 ( 
.A1(n_1891),
.A2(n_444),
.A3(n_445),
.B(n_443),
.Y(n_1944)
);

BUFx12f_ASAP7_75t_L g1945 ( 
.A(n_1773),
.Y(n_1945)
);

OAI21x1_ASAP7_75t_L g1946 ( 
.A1(n_1836),
.A2(n_448),
.B(n_447),
.Y(n_1946)
);

OAI21x1_ASAP7_75t_L g1947 ( 
.A1(n_1789),
.A2(n_451),
.B(n_450),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1858),
.Y(n_1948)
);

AO21x2_ASAP7_75t_L g1949 ( 
.A1(n_1744),
.A2(n_453),
.B(n_452),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1854),
.A2(n_128),
.B(n_129),
.Y(n_1950)
);

OAI21x1_ASAP7_75t_L g1951 ( 
.A1(n_1788),
.A2(n_456),
.B(n_455),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1803),
.B(n_128),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1856),
.B(n_130),
.Y(n_1953)
);

NOR2x1_ASAP7_75t_L g1954 ( 
.A(n_1798),
.B(n_130),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1768),
.A2(n_131),
.B(n_132),
.Y(n_1955)
);

OAI21x1_ASAP7_75t_L g1956 ( 
.A1(n_1893),
.A2(n_1816),
.B(n_1811),
.Y(n_1956)
);

INVxp67_ASAP7_75t_SL g1957 ( 
.A(n_1874),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1757),
.A2(n_131),
.B(n_132),
.Y(n_1958)
);

AOI211x1_ASAP7_75t_L g1959 ( 
.A1(n_1801),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1887),
.B(n_133),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1818),
.A2(n_134),
.B(n_135),
.Y(n_1961)
);

OAI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1793),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1760),
.A2(n_138),
.B(n_139),
.Y(n_1963)
);

AOI21x1_ASAP7_75t_L g1964 ( 
.A1(n_1849),
.A2(n_139),
.B(n_140),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1888),
.Y(n_1965)
);

NAND3xp33_ASAP7_75t_SL g1966 ( 
.A(n_1855),
.B(n_140),
.C(n_142),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1786),
.A2(n_143),
.B(n_144),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1784),
.B(n_143),
.Y(n_1968)
);

A2O1A1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1781),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1850),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1755),
.Y(n_1971)
);

OR2x6_ASAP7_75t_L g1972 ( 
.A(n_1863),
.B(n_1784),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1871),
.B(n_145),
.Y(n_1973)
);

AND3x4_ASAP7_75t_L g1974 ( 
.A(n_1870),
.B(n_146),
.C(n_147),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1851),
.B(n_148),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1774),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1777),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1792),
.Y(n_1978)
);

CKINVDCx8_ASAP7_75t_R g1979 ( 
.A(n_1777),
.Y(n_1979)
);

A2O1A1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1892),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1839),
.B(n_461),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1800),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1839),
.B(n_1763),
.Y(n_1983)
);

A2O1A1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1809),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_1984)
);

BUFx3_ASAP7_75t_L g1985 ( 
.A(n_1777),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1839),
.B(n_462),
.Y(n_1986)
);

OAI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1824),
.A2(n_464),
.B(n_463),
.Y(n_1987)
);

NAND2x1p5_ASAP7_75t_L g1988 ( 
.A(n_1782),
.B(n_465),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1815),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1863),
.A2(n_152),
.B(n_153),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1739),
.B(n_154),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1820),
.A2(n_154),
.B(n_155),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1846),
.A2(n_155),
.B(n_156),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1870),
.B(n_156),
.Y(n_1994)
);

NOR2xp67_ASAP7_75t_L g1995 ( 
.A(n_1763),
.B(n_158),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1877),
.B(n_158),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1782),
.Y(n_1997)
);

AO31x2_ASAP7_75t_L g1998 ( 
.A1(n_1862),
.A2(n_1890),
.A3(n_1805),
.B(n_1865),
.Y(n_1998)
);

OAI21xp33_ASAP7_75t_L g1999 ( 
.A1(n_1783),
.A2(n_159),
.B(n_160),
.Y(n_1999)
);

AOI21x1_ASAP7_75t_L g2000 ( 
.A1(n_1861),
.A2(n_1880),
.B(n_1876),
.Y(n_2000)
);

OAI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1882),
.A2(n_467),
.B(n_466),
.Y(n_2001)
);

NOR2xp67_ASAP7_75t_L g2002 ( 
.A(n_1810),
.B(n_159),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1814),
.A2(n_160),
.B(n_161),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1919),
.B(n_1797),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1907),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1899),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_SL g2007 ( 
.A(n_1902),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1965),
.B(n_1810),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1926),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1928),
.B(n_1878),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1922),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1972),
.Y(n_2012)
);

A2O1A1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_1930),
.A2(n_1840),
.B(n_1829),
.C(n_1828),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1914),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1970),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1903),
.B(n_1911),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1972),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1971),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1982),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1935),
.A2(n_1868),
.B1(n_1817),
.B2(n_1769),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1916),
.A2(n_1835),
.B(n_1894),
.Y(n_2021)
);

O2A1O1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1984),
.A2(n_1761),
.B(n_1813),
.C(n_1825),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1929),
.B(n_1873),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1901),
.B(n_1873),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1913),
.A2(n_1900),
.B(n_1910),
.Y(n_2025)
);

NAND2x1p5_ASAP7_75t_L g2026 ( 
.A(n_1983),
.B(n_1864),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1936),
.A2(n_1847),
.B(n_1844),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1960),
.A2(n_1843),
.B1(n_1886),
.B2(n_1737),
.Y(n_2028)
);

CKINVDCx20_ASAP7_75t_R g2029 ( 
.A(n_1918),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1927),
.B(n_1831),
.Y(n_2030)
);

A2O1A1Ixp33_ASAP7_75t_L g2031 ( 
.A1(n_1904),
.A2(n_1776),
.B(n_1885),
.C(n_1841),
.Y(n_2031)
);

A2O1A1Ixp33_ASAP7_75t_SL g2032 ( 
.A1(n_1932),
.A2(n_1869),
.B(n_1819),
.C(n_1834),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1934),
.A2(n_1826),
.B1(n_1875),
.B2(n_1822),
.Y(n_2033)
);

AND2x2_ASAP7_75t_SL g2034 ( 
.A(n_1981),
.B(n_1749),
.Y(n_2034)
);

O2A1O1Ixp5_ASAP7_75t_L g2035 ( 
.A1(n_1950),
.A2(n_1833),
.B(n_1770),
.C(n_1852),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1908),
.Y(n_2036)
);

NAND2xp33_ASAP7_75t_L g2037 ( 
.A(n_1999),
.B(n_1864),
.Y(n_2037)
);

OR2x2_ASAP7_75t_SL g2038 ( 
.A(n_1991),
.B(n_1782),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1905),
.A2(n_1758),
.B(n_1884),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1983),
.B(n_1864),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1918),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1925),
.A2(n_1807),
.B(n_1745),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1977),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1976),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1978),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2003),
.A2(n_1848),
.B(n_1837),
.Y(n_2046)
);

INVx1_ASAP7_75t_SL g2047 ( 
.A(n_1985),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_1917),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1955),
.A2(n_1879),
.B(n_1897),
.Y(n_2049)
);

NAND2x1p5_ASAP7_75t_L g2050 ( 
.A(n_1981),
.B(n_1883),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1909),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1993),
.A2(n_1992),
.B(n_1961),
.Y(n_2052)
);

BUFx2_ASAP7_75t_SL g2053 ( 
.A(n_1979),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1912),
.Y(n_2054)
);

INVx2_ASAP7_75t_SL g2055 ( 
.A(n_1912),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1956),
.A2(n_1889),
.B(n_1883),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1968),
.B(n_1883),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1973),
.B(n_1866),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1998),
.Y(n_2059)
);

CKINVDCx12_ASAP7_75t_R g2060 ( 
.A(n_1945),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1943),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1915),
.B(n_1872),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1989),
.Y(n_2063)
);

INVxp67_ASAP7_75t_SL g2064 ( 
.A(n_1957),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1942),
.B(n_1859),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1937),
.B(n_1867),
.Y(n_2066)
);

INVxp67_ASAP7_75t_SL g2067 ( 
.A(n_1898),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1931),
.B(n_1754),
.Y(n_2068)
);

BUFx4f_ASAP7_75t_SL g2069 ( 
.A(n_2029),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2005),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2020),
.A2(n_1980),
.B1(n_1974),
.B2(n_1959),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_2051),
.Y(n_2072)
);

BUFx2_ASAP7_75t_L g2073 ( 
.A(n_2036),
.Y(n_2073)
);

OAI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2028),
.A2(n_1966),
.B1(n_1967),
.B2(n_1990),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_2052),
.A2(n_1962),
.B1(n_1931),
.B2(n_1949),
.Y(n_2075)
);

INVx6_ASAP7_75t_L g2076 ( 
.A(n_2012),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_SL g2077 ( 
.A1(n_2034),
.A2(n_2046),
.B1(n_2033),
.B2(n_2062),
.Y(n_2077)
);

INVx4_ASAP7_75t_L g2078 ( 
.A(n_2043),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_SL g2079 ( 
.A1(n_2034),
.A2(n_1952),
.B1(n_1939),
.B2(n_1996),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_2012),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_SL g2081 ( 
.A1(n_2060),
.A2(n_1994),
.B1(n_1954),
.B2(n_1975),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2009),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2036),
.B(n_1953),
.Y(n_2083)
);

INVx1_ASAP7_75t_SL g2084 ( 
.A(n_2006),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2004),
.B(n_1942),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_SL g2086 ( 
.A1(n_2062),
.A2(n_1986),
.B1(n_1933),
.B2(n_1906),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_2041),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_2014),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_2061),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2016),
.B(n_1924),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2048),
.B(n_1924),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_SL g2092 ( 
.A1(n_2042),
.A2(n_1986),
.B1(n_1958),
.B2(n_1963),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_2054),
.Y(n_2093)
);

INVx4_ASAP7_75t_L g2094 ( 
.A(n_2007),
.Y(n_2094)
);

BUFx2_ASAP7_75t_SL g2095 ( 
.A(n_2007),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_2068),
.A2(n_2002),
.B1(n_1995),
.B2(n_1987),
.Y(n_2096)
);

INVx8_ASAP7_75t_L g2097 ( 
.A(n_2065),
.Y(n_2097)
);

OAI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_2039),
.A2(n_2021),
.B1(n_2068),
.B2(n_2027),
.Y(n_2098)
);

AOI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_2020),
.A2(n_1923),
.B1(n_2001),
.B2(n_1946),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2058),
.A2(n_1938),
.B1(n_1948),
.B2(n_1940),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2063),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_2047),
.Y(n_2102)
);

INVx1_ASAP7_75t_SL g2103 ( 
.A(n_2008),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_2057),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2011),
.A2(n_1920),
.B1(n_1921),
.B2(n_1942),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2013),
.A2(n_1969),
.B1(n_1964),
.B2(n_2000),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2031),
.A2(n_1988),
.B(n_1951),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2103),
.B(n_2048),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2091),
.Y(n_2109)
);

NOR2xp67_ASAP7_75t_L g2110 ( 
.A(n_2094),
.B(n_2055),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2073),
.B(n_2104),
.Y(n_2111)
);

CKINVDCx11_ASAP7_75t_R g2112 ( 
.A(n_2087),
.Y(n_2112)
);

O2A1O1Ixp33_ASAP7_75t_L g2113 ( 
.A1(n_2098),
.A2(n_2032),
.B(n_2031),
.C(n_2022),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2070),
.Y(n_2114)
);

O2A1O1Ixp33_ASAP7_75t_L g2115 ( 
.A1(n_2071),
.A2(n_2032),
.B(n_2022),
.C(n_2037),
.Y(n_2115)
);

OA21x2_ASAP7_75t_L g2116 ( 
.A1(n_2090),
.A2(n_2025),
.B(n_2059),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_2069),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2085),
.B(n_2024),
.Y(n_2118)
);

A2O1A1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_2077),
.A2(n_2049),
.B(n_2066),
.C(n_2030),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_2106),
.A2(n_2056),
.B(n_2067),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_SL g2121 ( 
.A(n_2094),
.B(n_2012),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2082),
.B(n_2023),
.Y(n_2122)
);

OR2x6_ASAP7_75t_L g2123 ( 
.A(n_2097),
.B(n_2012),
.Y(n_2123)
);

AOI21x1_ASAP7_75t_SL g2124 ( 
.A1(n_2083),
.A2(n_2010),
.B(n_2040),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2101),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2076),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2080),
.Y(n_2127)
);

AOI211xp5_ASAP7_75t_L g2128 ( 
.A1(n_2074),
.A2(n_2010),
.B(n_2015),
.C(n_2017),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2077),
.B(n_2064),
.Y(n_2129)
);

O2A1O1Ixp5_ASAP7_75t_L g2130 ( 
.A1(n_2074),
.A2(n_2065),
.B(n_2035),
.C(n_2067),
.Y(n_2130)
);

NOR2xp67_ASAP7_75t_R g2131 ( 
.A(n_2121),
.B(n_2078),
.Y(n_2131)
);

NAND2xp33_ASAP7_75t_R g2132 ( 
.A(n_2129),
.B(n_2102),
.Y(n_2132)
);

AO31x2_ASAP7_75t_L g2133 ( 
.A1(n_2120),
.A2(n_2019),
.A3(n_2044),
.B(n_2018),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_2116),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2114),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2108),
.B(n_2038),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2111),
.B(n_2072),
.Y(n_2137)
);

BUFx3_ASAP7_75t_L g2138 ( 
.A(n_2117),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2135),
.Y(n_2139)
);

OR2x6_ASAP7_75t_L g2140 ( 
.A(n_2138),
.B(n_2095),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2137),
.B(n_2111),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2135),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2137),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2136),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2143),
.B(n_2144),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2141),
.B(n_2119),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2139),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2140),
.A2(n_2113),
.B1(n_2128),
.B2(n_2115),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2140),
.B(n_2110),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2139),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_2142),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2139),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2141),
.B(n_2138),
.Y(n_2153)
);

AND2x4_ASAP7_75t_L g2154 ( 
.A(n_2153),
.B(n_2117),
.Y(n_2154)
);

AOI211xp5_ASAP7_75t_L g2155 ( 
.A1(n_2148),
.A2(n_2081),
.B(n_2134),
.C(n_2107),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2150),
.Y(n_2156)
);

AO21x2_ASAP7_75t_L g2157 ( 
.A1(n_2147),
.A2(n_2150),
.B(n_2152),
.Y(n_2157)
);

OA21x2_ASAP7_75t_L g2158 ( 
.A1(n_2147),
.A2(n_2130),
.B(n_2109),
.Y(n_2158)
);

AOI211xp5_ASAP7_75t_L g2159 ( 
.A1(n_2146),
.A2(n_2134),
.B(n_2132),
.C(n_2136),
.Y(n_2159)
);

NOR2x1p5_ASAP7_75t_L g2160 ( 
.A(n_2145),
.B(n_2078),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2151),
.A2(n_2134),
.B1(n_2075),
.B2(n_2086),
.Y(n_2161)
);

AOI222xp33_ASAP7_75t_L g2162 ( 
.A1(n_2151),
.A2(n_2134),
.B1(n_2109),
.B2(n_2096),
.C1(n_2059),
.C2(n_2133),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2149),
.A2(n_2079),
.B1(n_2086),
.B2(n_2092),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2153),
.B(n_2112),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2154),
.B(n_2084),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2157),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2157),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2156),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2154),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2164),
.B(n_2114),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2160),
.B(n_2161),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2159),
.B(n_2093),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2155),
.B(n_2089),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2166),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2170),
.B(n_2169),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2166),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2167),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2175),
.B(n_2170),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2177),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2174),
.A2(n_2163),
.B1(n_2158),
.B2(n_2173),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2176),
.B(n_2168),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_SL g2182 ( 
.A1(n_2179),
.A2(n_2158),
.B1(n_2173),
.B2(n_2172),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2178),
.B(n_2165),
.Y(n_2183)
);

NAND2x2_ASAP7_75t_L g2184 ( 
.A(n_2181),
.B(n_2171),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2180),
.B(n_2165),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2178),
.B(n_2172),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2178),
.B(n_2088),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2182),
.B(n_2163),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_2187),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2183),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2184),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2185),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2186),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2187),
.B(n_2162),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2184),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2186),
.B(n_2133),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2186),
.B(n_2133),
.Y(n_2197)
);

OAI221xp5_ASAP7_75t_L g2198 ( 
.A1(n_2188),
.A2(n_2192),
.B1(n_2195),
.B2(n_2191),
.C(n_2196),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2189),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2190),
.A2(n_2079),
.B1(n_2092),
.B2(n_2100),
.Y(n_2200)
);

INVx1_ASAP7_75t_SL g2201 ( 
.A(n_2190),
.Y(n_2201)
);

O2A1O1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2188),
.A2(n_2035),
.B(n_2108),
.C(n_2099),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2194),
.A2(n_2053),
.B1(n_2126),
.B2(n_2116),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2193),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2197),
.Y(n_2205)
);

OAI21xp5_ASAP7_75t_SL g2206 ( 
.A1(n_2192),
.A2(n_2131),
.B(n_2127),
.Y(n_2206)
);

NOR3xp33_ASAP7_75t_L g2207 ( 
.A(n_2192),
.B(n_1766),
.C(n_2127),
.Y(n_2207)
);

OAI22xp33_ASAP7_75t_SL g2208 ( 
.A1(n_2188),
.A2(n_2076),
.B1(n_2050),
.B2(n_2123),
.Y(n_2208)
);

OAI32xp33_ASAP7_75t_L g2209 ( 
.A1(n_2188),
.A2(n_2050),
.A3(n_2122),
.B1(n_2118),
.B2(n_2026),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_2189),
.Y(n_2210)
);

NAND3xp33_ASAP7_75t_L g2211 ( 
.A(n_2199),
.B(n_2116),
.C(n_2017),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_2210),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2201),
.Y(n_2213)
);

O2A1O1Ixp33_ASAP7_75t_L g2214 ( 
.A1(n_2198),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2204),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2205),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2200),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_2203),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2202),
.B(n_2133),
.Y(n_2219)
);

OAI211xp5_ASAP7_75t_L g2220 ( 
.A1(n_2206),
.A2(n_165),
.B(n_162),
.C(n_164),
.Y(n_2220)
);

INVxp33_ASAP7_75t_L g2221 ( 
.A(n_2207),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2209),
.A2(n_2116),
.B1(n_2122),
.B2(n_2118),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2208),
.A2(n_2017),
.B1(n_2125),
.B2(n_2076),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2210),
.B(n_2133),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_SL g2225 ( 
.A1(n_2201),
.A2(n_2017),
.B1(n_1920),
.B2(n_1921),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_2212),
.B(n_1997),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2219),
.A2(n_2080),
.B1(n_2125),
.B2(n_1997),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2213),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2215),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2214),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2216),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2221),
.B(n_2133),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2224),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2220),
.B(n_164),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2218),
.B(n_165),
.Y(n_2235)
);

NAND2xp33_ASAP7_75t_L g2236 ( 
.A(n_2217),
.B(n_2222),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2211),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2225),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2223),
.B(n_2123),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2231),
.B(n_166),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2234),
.Y(n_2241)
);

NOR3xp33_ASAP7_75t_L g2242 ( 
.A(n_2228),
.B(n_166),
.C(n_167),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2235),
.B(n_167),
.Y(n_2243)
);

NAND3xp33_ASAP7_75t_SL g2244 ( 
.A(n_2230),
.B(n_1764),
.C(n_2105),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2229),
.B(n_1997),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2226),
.B(n_2123),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2237),
.B(n_168),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2236),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_2238),
.B(n_169),
.Y(n_2249)
);

AOI211x1_ASAP7_75t_L g2250 ( 
.A1(n_2233),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2232),
.A2(n_2080),
.B1(n_2123),
.B2(n_2040),
.Y(n_2251)
);

AOI221xp5_ASAP7_75t_L g2252 ( 
.A1(n_2227),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.C(n_176),
.Y(n_2252)
);

INVxp67_ASAP7_75t_L g2253 ( 
.A(n_2239),
.Y(n_2253)
);

NOR3xp33_ASAP7_75t_L g2254 ( 
.A(n_2239),
.B(n_173),
.C(n_176),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2234),
.B(n_177),
.Y(n_2255)
);

INVxp33_ASAP7_75t_L g2256 ( 
.A(n_2235),
.Y(n_2256)
);

INVxp67_ASAP7_75t_SL g2257 ( 
.A(n_2235),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_SL g2258 ( 
.A(n_2228),
.B(n_177),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_2234),
.B(n_178),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2231),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2234),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2248),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2260),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_2258),
.B(n_178),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2250),
.Y(n_2265)
);

O2A1O1Ixp5_ASAP7_75t_L g2266 ( 
.A1(n_2245),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_2266)
);

NAND4xp25_ASAP7_75t_L g2267 ( 
.A(n_2249),
.B(n_2254),
.C(n_2259),
.D(n_2255),
.Y(n_2267)
);

NAND2xp33_ASAP7_75t_SL g2268 ( 
.A(n_2240),
.B(n_179),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2256),
.B(n_2247),
.Y(n_2269)
);

NOR4xp25_ASAP7_75t_L g2270 ( 
.A(n_2241),
.B(n_182),
.C(n_180),
.D(n_181),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2243),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2257),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2246),
.B(n_182),
.Y(n_2273)
);

XNOR2xp5_ASAP7_75t_L g2274 ( 
.A(n_2261),
.B(n_183),
.Y(n_2274)
);

O2A1O1Ixp5_ASAP7_75t_SL g2275 ( 
.A1(n_2253),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2242),
.Y(n_2276)
);

OAI211xp5_ASAP7_75t_SL g2277 ( 
.A1(n_2252),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2244),
.B(n_187),
.Y(n_2278)
);

OAI211xp5_ASAP7_75t_L g2279 ( 
.A1(n_2251),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_2279)
);

AOI221xp5_ASAP7_75t_L g2280 ( 
.A1(n_2260),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2248),
.Y(n_2281)
);

AOI222xp33_ASAP7_75t_L g2282 ( 
.A1(n_2253),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.C1(n_194),
.C2(n_195),
.Y(n_2282)
);

INVxp67_ASAP7_75t_SL g2283 ( 
.A(n_2248),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2250),
.B(n_192),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_2258),
.Y(n_2285)
);

NAND3xp33_ASAP7_75t_SL g2286 ( 
.A(n_2258),
.B(n_194),
.C(n_196),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2248),
.Y(n_2287)
);

XNOR2xp5_ASAP7_75t_L g2288 ( 
.A(n_2250),
.B(n_197),
.Y(n_2288)
);

OAI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2260),
.A2(n_1947),
.B(n_1941),
.Y(n_2289)
);

NOR3xp33_ASAP7_75t_L g2290 ( 
.A(n_2260),
.B(n_198),
.C(n_200),
.Y(n_2290)
);

NOR2x1_ASAP7_75t_L g2291 ( 
.A(n_2248),
.B(n_200),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2248),
.B(n_201),
.Y(n_2292)
);

NAND5xp2_ASAP7_75t_L g2293 ( 
.A(n_2248),
.B(n_203),
.C(n_201),
.D(n_202),
.E(n_204),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_2258),
.B(n_202),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2248),
.B(n_2080),
.Y(n_2295)
);

AOI221x1_ASAP7_75t_L g2296 ( 
.A1(n_2248),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.C(n_206),
.Y(n_2296)
);

AOI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2248),
.A2(n_205),
.B(n_206),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_2248),
.Y(n_2298)
);

AOI221xp5_ASAP7_75t_L g2299 ( 
.A1(n_2263),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.C(n_210),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2263),
.B(n_207),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2291),
.B(n_208),
.Y(n_2301)
);

OAI221xp5_ASAP7_75t_L g2302 ( 
.A1(n_2283),
.A2(n_213),
.B1(n_210),
.B2(n_211),
.C(n_214),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2263),
.A2(n_2097),
.B1(n_2064),
.B2(n_2026),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2270),
.B(n_211),
.Y(n_2304)
);

AOI222xp33_ASAP7_75t_L g2305 ( 
.A1(n_2272),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.C1(n_216),
.C2(n_217),
.Y(n_2305)
);

NOR3xp33_ASAP7_75t_L g2306 ( 
.A(n_2262),
.B(n_2287),
.C(n_2281),
.Y(n_2306)
);

OAI322xp33_ASAP7_75t_L g2307 ( 
.A1(n_2295),
.A2(n_215),
.A3(n_217),
.B1(n_218),
.B2(n_219),
.C1(n_220),
.C2(n_221),
.Y(n_2307)
);

NAND2x1_ASAP7_75t_SL g2308 ( 
.A(n_2265),
.B(n_219),
.Y(n_2308)
);

A2O1A1Ixp33_ASAP7_75t_L g2309 ( 
.A1(n_2264),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2269),
.A2(n_2097),
.B1(n_2124),
.B2(n_2045),
.Y(n_2310)
);

AOI211xp5_ASAP7_75t_L g2311 ( 
.A1(n_2279),
.A2(n_226),
.B(n_222),
.C(n_223),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2288),
.Y(n_2312)
);

AOI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2271),
.A2(n_2298),
.B1(n_2273),
.B2(n_2294),
.Y(n_2313)
);

OAI21xp5_ASAP7_75t_SL g2314 ( 
.A1(n_2284),
.A2(n_226),
.B(n_227),
.Y(n_2314)
);

OR3x1_ASAP7_75t_L g2315 ( 
.A(n_2286),
.B(n_227),
.C(n_228),
.Y(n_2315)
);

OAI221xp5_ASAP7_75t_L g2316 ( 
.A1(n_2266),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_2316)
);

NAND3xp33_ASAP7_75t_L g2317 ( 
.A(n_2268),
.B(n_229),
.C(n_231),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2297),
.A2(n_2293),
.B(n_2274),
.Y(n_2318)
);

NAND4xp75_ASAP7_75t_L g2319 ( 
.A(n_2276),
.B(n_234),
.C(n_232),
.D(n_233),
.Y(n_2319)
);

AOI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2292),
.A2(n_233),
.B(n_235),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2296),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2282),
.B(n_235),
.Y(n_2322)
);

NOR2x1_ASAP7_75t_L g2323 ( 
.A(n_2267),
.B(n_236),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2290),
.B(n_236),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_SL g2325 ( 
.A(n_2285),
.B(n_237),
.Y(n_2325)
);

AOI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2277),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_2326)
);

NAND5xp2_ASAP7_75t_L g2327 ( 
.A(n_2278),
.B(n_2280),
.C(n_2289),
.D(n_2275),
.E(n_242),
.Y(n_2327)
);

OAI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2283),
.A2(n_243),
.B1(n_240),
.B2(n_241),
.C(n_244),
.Y(n_2328)
);

NAND4xp25_ASAP7_75t_L g2329 ( 
.A(n_2262),
.B(n_244),
.C(n_240),
.D(n_241),
.Y(n_2329)
);

O2A1O1Ixp5_ASAP7_75t_L g2330 ( 
.A1(n_2283),
.A2(n_248),
.B(n_245),
.C(n_246),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2283),
.A2(n_248),
.B1(n_245),
.B2(n_246),
.Y(n_2331)
);

AOI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2306),
.A2(n_249),
.B(n_250),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2321),
.B(n_249),
.Y(n_2333)
);

AOI322xp5_ASAP7_75t_L g2334 ( 
.A1(n_2312),
.A2(n_1944),
.A3(n_251),
.B1(n_252),
.B2(n_253),
.C1(n_254),
.C2(n_256),
.Y(n_2334)
);

NOR3xp33_ASAP7_75t_L g2335 ( 
.A(n_2313),
.B(n_250),
.C(n_251),
.Y(n_2335)
);

AOI22xp33_ASAP7_75t_SL g2336 ( 
.A1(n_2304),
.A2(n_1944),
.B1(n_254),
.B2(n_252),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2301),
.B(n_253),
.C(n_257),
.Y(n_2337)
);

OAI211xp5_ASAP7_75t_SL g2338 ( 
.A1(n_2323),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2308),
.B(n_258),
.Y(n_2339)
);

NOR3xp33_ASAP7_75t_SL g2340 ( 
.A(n_2314),
.B(n_260),
.C(n_261),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2300),
.B(n_261),
.C(n_263),
.Y(n_2341)
);

AOI211xp5_ASAP7_75t_L g2342 ( 
.A1(n_2316),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_2305),
.B(n_264),
.Y(n_2343)
);

NOR4xp25_ASAP7_75t_L g2344 ( 
.A(n_2322),
.B(n_268),
.C(n_266),
.D(n_267),
.Y(n_2344)
);

XNOR2x2_ASAP7_75t_L g2345 ( 
.A(n_2329),
.B(n_266),
.Y(n_2345)
);

AOI211xp5_ASAP7_75t_SL g2346 ( 
.A1(n_2307),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2311),
.B(n_2330),
.Y(n_2347)
);

NOR3xp33_ASAP7_75t_SL g2348 ( 
.A(n_2327),
.B(n_2317),
.C(n_2318),
.Y(n_2348)
);

NAND5xp2_ASAP7_75t_L g2349 ( 
.A(n_2326),
.B(n_270),
.C(n_271),
.D(n_272),
.E(n_273),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_L g2350 ( 
.A(n_2325),
.B(n_270),
.C(n_271),
.Y(n_2350)
);

NOR2x1_ASAP7_75t_L g2351 ( 
.A(n_2319),
.B(n_2331),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2315),
.B(n_272),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2299),
.B(n_273),
.Y(n_2353)
);

AOI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2324),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.C(n_278),
.Y(n_2354)
);

NOR3xp33_ASAP7_75t_L g2355 ( 
.A(n_2320),
.B(n_274),
.C(n_276),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2309),
.B(n_279),
.Y(n_2356)
);

NOR3xp33_ASAP7_75t_L g2357 ( 
.A(n_2302),
.B(n_279),
.C(n_280),
.Y(n_2357)
);

NOR3xp33_ASAP7_75t_L g2358 ( 
.A(n_2328),
.B(n_281),
.C(n_282),
.Y(n_2358)
);

NOR3xp33_ASAP7_75t_SL g2359 ( 
.A(n_2303),
.B(n_281),
.C(n_282),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2310),
.B(n_283),
.Y(n_2360)
);

NAND4xp25_ASAP7_75t_L g2361 ( 
.A(n_2306),
.B(n_285),
.C(n_283),
.D(n_284),
.Y(n_2361)
);

NOR3xp33_ASAP7_75t_L g2362 ( 
.A(n_2306),
.B(n_284),
.C(n_285),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2321),
.B(n_286),
.Y(n_2363)
);

NAND3xp33_ASAP7_75t_SL g2364 ( 
.A(n_2306),
.B(n_287),
.C(n_288),
.Y(n_2364)
);

OAI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2321),
.A2(n_288),
.B(n_289),
.Y(n_2365)
);

NAND4xp25_ASAP7_75t_L g2366 ( 
.A(n_2306),
.B(n_291),
.C(n_289),
.D(n_290),
.Y(n_2366)
);

AOI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2306),
.A2(n_290),
.B(n_293),
.Y(n_2367)
);

AND2x2_ASAP7_75t_SL g2368 ( 
.A(n_2306),
.B(n_295),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2308),
.Y(n_2369)
);

NAND3xp33_ASAP7_75t_L g2370 ( 
.A(n_2306),
.B(n_295),
.C(n_296),
.Y(n_2370)
);

AOI21xp33_ASAP7_75t_SL g2371 ( 
.A1(n_2306),
.A2(n_296),
.B(n_297),
.Y(n_2371)
);

NAND4xp25_ASAP7_75t_SL g2372 ( 
.A(n_2306),
.B(n_300),
.C(n_297),
.D(n_298),
.Y(n_2372)
);

NOR2x1_ASAP7_75t_L g2373 ( 
.A(n_2300),
.B(n_298),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2321),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_2374)
);

OAI221xp5_ASAP7_75t_L g2375 ( 
.A1(n_2306),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.C(n_306),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2306),
.B(n_304),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2321),
.A2(n_310),
.B1(n_306),
.B2(n_308),
.Y(n_2377)
);

OAI211xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2313),
.A2(n_311),
.B(n_308),
.C(n_310),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2308),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2306),
.A2(n_311),
.B(n_312),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2306),
.A2(n_312),
.B(n_313),
.Y(n_2381)
);

AOI221xp5_ASAP7_75t_L g2382 ( 
.A1(n_2306),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.C(n_316),
.Y(n_2382)
);

CKINVDCx16_ASAP7_75t_R g2383 ( 
.A(n_2369),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2348),
.B(n_314),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2379),
.B(n_315),
.Y(n_2385)
);

NAND2xp33_ASAP7_75t_R g2386 ( 
.A(n_2376),
.B(n_2333),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2339),
.Y(n_2387)
);

OAI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2363),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2388)
);

NAND2xp33_ASAP7_75t_SL g2389 ( 
.A(n_2340),
.B(n_319),
.Y(n_2389)
);

NAND2xp33_ASAP7_75t_L g2390 ( 
.A(n_2335),
.B(n_319),
.Y(n_2390)
);

OAI211xp5_ASAP7_75t_L g2391 ( 
.A1(n_2365),
.A2(n_2352),
.B(n_2367),
.C(n_2332),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2344),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.C(n_323),
.Y(n_2392)
);

AOI31xp33_ASAP7_75t_L g2393 ( 
.A1(n_2346),
.A2(n_2370),
.A3(n_2342),
.B(n_2373),
.Y(n_2393)
);

AOI221x1_ASAP7_75t_L g2394 ( 
.A1(n_2357),
.A2(n_320),
.B1(n_321),
.B2(n_323),
.C(n_324),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2359),
.B(n_324),
.Y(n_2395)
);

OAI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_2338),
.A2(n_325),
.B(n_326),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2368),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2345),
.Y(n_2398)
);

AOI221x1_ASAP7_75t_L g2399 ( 
.A1(n_2358),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.C(n_330),
.Y(n_2399)
);

NOR2xp67_ASAP7_75t_L g2400 ( 
.A(n_2372),
.B(n_2361),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_2349),
.B(n_330),
.Y(n_2401)
);

NAND2xp33_ASAP7_75t_L g2402 ( 
.A(n_2362),
.B(n_331),
.Y(n_2402)
);

AOI222xp33_ASAP7_75t_L g2403 ( 
.A1(n_2347),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.C1(n_334),
.C2(n_335),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2355),
.Y(n_2404)
);

INVx5_ASAP7_75t_L g2405 ( 
.A(n_2337),
.Y(n_2405)
);

XOR2xp5_ASAP7_75t_L g2406 ( 
.A(n_2366),
.B(n_332),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_SL g2407 ( 
.A(n_2371),
.B(n_333),
.C(n_334),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2378),
.B(n_2364),
.Y(n_2408)
);

AOI22x1_ASAP7_75t_L g2409 ( 
.A1(n_2380),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_2409)
);

OAI22x1_ASAP7_75t_L g2410 ( 
.A1(n_2350),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2336),
.B(n_338),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2341),
.B(n_339),
.Y(n_2412)
);

NAND4xp75_ASAP7_75t_L g2413 ( 
.A(n_2351),
.B(n_340),
.C(n_341),
.D(n_342),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2343),
.Y(n_2414)
);

AO22x2_ASAP7_75t_L g2415 ( 
.A1(n_2374),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2356),
.B(n_2381),
.Y(n_2416)
);

OAI221xp5_ASAP7_75t_L g2417 ( 
.A1(n_2377),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.C(n_346),
.Y(n_2417)
);

HB1xp67_ASAP7_75t_L g2418 ( 
.A(n_2375),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2353),
.Y(n_2419)
);

AOI211xp5_ASAP7_75t_L g2420 ( 
.A1(n_2354),
.A2(n_2382),
.B(n_2360),
.C(n_2334),
.Y(n_2420)
);

INVx1_ASAP7_75t_SL g2421 ( 
.A(n_2368),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2369),
.B(n_343),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2339),
.Y(n_2423)
);

A2O1A1Ixp33_ASAP7_75t_L g2424 ( 
.A1(n_2346),
.A2(n_344),
.B(n_345),
.C(n_347),
.Y(n_2424)
);

OAI211xp5_ASAP7_75t_L g2425 ( 
.A1(n_2365),
.A2(n_348),
.B(n_349),
.C(n_350),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2339),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_2373),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_L g2428 ( 
.A(n_2369),
.B(n_348),
.Y(n_2428)
);

NAND2xp33_ASAP7_75t_SL g2429 ( 
.A(n_2340),
.B(n_349),
.Y(n_2429)
);

NOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2398),
.B(n_350),
.Y(n_2430)
);

OR2x2_ASAP7_75t_L g2431 ( 
.A(n_2383),
.B(n_351),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2421),
.B(n_351),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2384),
.B(n_352),
.Y(n_2433)
);

HB1xp67_ASAP7_75t_L g2434 ( 
.A(n_2427),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2395),
.Y(n_2435)
);

OAI21xp5_ASAP7_75t_SL g2436 ( 
.A1(n_2401),
.A2(n_352),
.B(n_354),
.Y(n_2436)
);

XOR2x1_ASAP7_75t_L g2437 ( 
.A(n_2384),
.B(n_355),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2395),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2415),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2400),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2415),
.Y(n_2441)
);

XOR2xp5_ASAP7_75t_L g2442 ( 
.A(n_2406),
.B(n_2404),
.Y(n_2442)
);

XNOR2x1_ASAP7_75t_L g2443 ( 
.A(n_2387),
.B(n_356),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_SL g2444 ( 
.A(n_2428),
.B(n_357),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2423),
.B(n_358),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2405),
.B(n_358),
.Y(n_2446)
);

NOR3xp33_ASAP7_75t_SL g2447 ( 
.A(n_2386),
.B(n_359),
.C(n_360),
.Y(n_2447)
);

NOR2x1_ASAP7_75t_L g2448 ( 
.A(n_2413),
.B(n_359),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2397),
.Y(n_2449)
);

AOI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2408),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_2450)
);

NAND4xp75_ASAP7_75t_L g2451 ( 
.A(n_2414),
.B(n_362),
.C(n_363),
.D(n_364),
.Y(n_2451)
);

XNOR2xp5_ASAP7_75t_L g2452 ( 
.A(n_2426),
.B(n_366),
.Y(n_2452)
);

AOI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2389),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2407),
.B(n_367),
.Y(n_2454)
);

NAND4xp75_ASAP7_75t_L g2455 ( 
.A(n_2394),
.B(n_369),
.C(n_370),
.D(n_371),
.Y(n_2455)
);

NOR2x1_ASAP7_75t_L g2456 ( 
.A(n_2385),
.B(n_2422),
.Y(n_2456)
);

NAND4xp75_ASAP7_75t_L g2457 ( 
.A(n_2399),
.B(n_369),
.C(n_370),
.D(n_372),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2405),
.B(n_372),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2405),
.Y(n_2459)
);

XNOR2x1_ASAP7_75t_L g2460 ( 
.A(n_2410),
.B(n_373),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2396),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2429),
.B(n_373),
.Y(n_2462)
);

NAND2x1p5_ASAP7_75t_L g2463 ( 
.A(n_2419),
.B(n_374),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2409),
.Y(n_2464)
);

NAND2x1p5_ASAP7_75t_L g2465 ( 
.A(n_2416),
.B(n_375),
.Y(n_2465)
);

NOR2x1_ASAP7_75t_L g2466 ( 
.A(n_2425),
.B(n_375),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2393),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2434),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2459),
.B(n_2418),
.Y(n_2469)
);

NAND4xp75_ASAP7_75t_L g2470 ( 
.A(n_2456),
.B(n_2412),
.C(n_2392),
.D(n_2411),
.Y(n_2470)
);

NOR5xp2_ASAP7_75t_L g2471 ( 
.A(n_2467),
.B(n_2391),
.C(n_2417),
.D(n_2424),
.E(n_2420),
.Y(n_2471)
);

INVxp67_ASAP7_75t_L g2472 ( 
.A(n_2430),
.Y(n_2472)
);

NOR3xp33_ASAP7_75t_L g2473 ( 
.A(n_2449),
.B(n_2388),
.C(n_2402),
.Y(n_2473)
);

AO22x2_ASAP7_75t_L g2474 ( 
.A1(n_2439),
.A2(n_2390),
.B1(n_2403),
.B2(n_378),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_2438),
.B(n_376),
.C(n_377),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2437),
.Y(n_2476)
);

NOR3xp33_ASAP7_75t_L g2477 ( 
.A(n_2435),
.B(n_376),
.C(n_377),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2441),
.B(n_378),
.Y(n_2478)
);

AO211x2_ASAP7_75t_L g2479 ( 
.A1(n_2446),
.A2(n_379),
.B(n_380),
.C(n_381),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_L g2480 ( 
.A(n_2458),
.B(n_380),
.C(n_382),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2462),
.B(n_382),
.Y(n_2481)
);

NOR4xp25_ASAP7_75t_L g2482 ( 
.A(n_2436),
.B(n_383),
.C(n_384),
.D(n_386),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2465),
.Y(n_2483)
);

NAND3xp33_ASAP7_75t_L g2484 ( 
.A(n_2431),
.B(n_383),
.C(n_384),
.Y(n_2484)
);

NOR4xp25_ASAP7_75t_L g2485 ( 
.A(n_2433),
.B(n_386),
.C(n_387),
.D(n_388),
.Y(n_2485)
);

A2O1A1Ixp33_ASAP7_75t_L g2486 ( 
.A1(n_2432),
.A2(n_387),
.B(n_389),
.C(n_390),
.Y(n_2486)
);

NOR3xp33_ASAP7_75t_SL g2487 ( 
.A(n_2455),
.B(n_389),
.C(n_390),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2463),
.Y(n_2488)
);

AND2x2_ASAP7_75t_SL g2489 ( 
.A(n_2454),
.B(n_391),
.Y(n_2489)
);

NAND3xp33_ASAP7_75t_SL g2490 ( 
.A(n_2442),
.B(n_391),
.C(n_393),
.Y(n_2490)
);

CKINVDCx16_ASAP7_75t_R g2491 ( 
.A(n_2444),
.Y(n_2491)
);

XOR2xp5_ASAP7_75t_L g2492 ( 
.A(n_2443),
.B(n_393),
.Y(n_2492)
);

NAND3xp33_ASAP7_75t_SL g2493 ( 
.A(n_2453),
.B(n_394),
.C(n_395),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2447),
.B(n_394),
.Y(n_2494)
);

INVx3_ASAP7_75t_L g2495 ( 
.A(n_2445),
.Y(n_2495)
);

AOI22xp33_ASAP7_75t_L g2496 ( 
.A1(n_2468),
.A2(n_2448),
.B1(n_2466),
.B2(n_2464),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2489),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2476),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2491),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2492),
.Y(n_2500)
);

CKINVDCx20_ASAP7_75t_R g2501 ( 
.A(n_2469),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_2472),
.Y(n_2502)
);

HB1xp67_ASAP7_75t_L g2503 ( 
.A(n_2495),
.Y(n_2503)
);

NOR2x1p5_ASAP7_75t_L g2504 ( 
.A(n_2490),
.B(n_2457),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2488),
.B(n_2461),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2483),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2487),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2485),
.B(n_2445),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2494),
.B(n_2452),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2474),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2478),
.B(n_2460),
.Y(n_2511)
);

INVx1_ASAP7_75t_SL g2512 ( 
.A(n_2481),
.Y(n_2512)
);

INVx2_ASAP7_75t_SL g2513 ( 
.A(n_2479),
.Y(n_2513)
);

BUFx2_ASAP7_75t_L g2514 ( 
.A(n_2474),
.Y(n_2514)
);

HB1xp67_ASAP7_75t_L g2515 ( 
.A(n_2470),
.Y(n_2515)
);

AOI22xp5_ASAP7_75t_SL g2516 ( 
.A1(n_2499),
.A2(n_2471),
.B1(n_2482),
.B2(n_2480),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_SL g2517 ( 
.A1(n_2501),
.A2(n_2484),
.B1(n_2473),
.B2(n_2493),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2503),
.B(n_2477),
.Y(n_2518)
);

OAI322xp33_ASAP7_75t_L g2519 ( 
.A1(n_2502),
.A2(n_2440),
.A3(n_2450),
.B1(n_2475),
.B2(n_2486),
.C1(n_2451),
.C2(n_400),
.Y(n_2519)
);

OAI322xp33_ASAP7_75t_L g2520 ( 
.A1(n_2497),
.A2(n_395),
.A3(n_396),
.B1(n_397),
.B2(n_398),
.C1(n_399),
.C2(n_400),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2505),
.B(n_396),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2510),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2514),
.Y(n_2523)
);

HB1xp67_ASAP7_75t_L g2524 ( 
.A(n_2515),
.Y(n_2524)
);

NAND3xp33_ASAP7_75t_L g2525 ( 
.A(n_2506),
.B(n_397),
.C(n_398),
.Y(n_2525)
);

AOI322xp5_ASAP7_75t_L g2526 ( 
.A1(n_2505),
.A2(n_399),
.A3(n_402),
.B1(n_403),
.B2(n_404),
.C1(n_405),
.C2(n_407),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2506),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2506),
.B(n_402),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_2498),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_L g2530 ( 
.A1(n_2513),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_2530)
);

AOI322xp5_ASAP7_75t_L g2531 ( 
.A1(n_2496),
.A2(n_407),
.A3(n_408),
.B1(n_409),
.B2(n_410),
.C1(n_411),
.C2(n_412),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2524),
.A2(n_2500),
.B1(n_2507),
.B2(n_2504),
.Y(n_2532)
);

AO22x2_ASAP7_75t_L g2533 ( 
.A1(n_2527),
.A2(n_2512),
.B1(n_2508),
.B2(n_2511),
.Y(n_2533)
);

AO22x2_ASAP7_75t_L g2534 ( 
.A1(n_2523),
.A2(n_2509),
.B1(n_409),
.B2(n_411),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2529),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2522),
.Y(n_2536)
);

AOI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2518),
.A2(n_408),
.B1(n_412),
.B2(n_413),
.Y(n_2537)
);

OAI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2517),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2538)
);

NAND5xp2_ASAP7_75t_L g2539 ( 
.A(n_2532),
.B(n_2516),
.C(n_2530),
.D(n_2519),
.E(n_2528),
.Y(n_2539)
);

OAI221xp5_ASAP7_75t_L g2540 ( 
.A1(n_2536),
.A2(n_2535),
.B1(n_2525),
.B2(n_2538),
.C(n_2537),
.Y(n_2540)
);

NAND3xp33_ASAP7_75t_L g2541 ( 
.A(n_2533),
.B(n_2521),
.C(n_2531),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2534),
.A2(n_2520),
.B1(n_2526),
.B2(n_417),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2536),
.A2(n_414),
.B1(n_416),
.B2(n_417),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2541),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2542),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2540),
.B(n_418),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_L g2547 ( 
.A(n_2544),
.B(n_2539),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_SL g2548 ( 
.A1(n_2545),
.A2(n_2543),
.B1(n_420),
.B2(n_421),
.Y(n_2548)
);

OAI21xp5_ASAP7_75t_L g2549 ( 
.A1(n_2546),
.A2(n_418),
.B(n_420),
.Y(n_2549)
);

AOI22xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2547),
.A2(n_2549),
.B1(n_2548),
.B2(n_423),
.Y(n_2550)
);

OAI22xp33_ASAP7_75t_L g2551 ( 
.A1(n_2547),
.A2(n_421),
.B1(n_422),
.B2(n_424),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2550),
.B(n_422),
.Y(n_2552)
);

NOR2x1_ASAP7_75t_L g2553 ( 
.A(n_2551),
.B(n_424),
.Y(n_2553)
);

AOI22xp5_ASAP7_75t_SL g2554 ( 
.A1(n_2552),
.A2(n_425),
.B1(n_426),
.B2(n_469),
.Y(n_2554)
);

AOI22xp33_ASAP7_75t_L g2555 ( 
.A1(n_2553),
.A2(n_425),
.B1(n_426),
.B2(n_470),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2554),
.B(n_471),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2556),
.B(n_2555),
.Y(n_2557)
);

AOI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2557),
.A2(n_474),
.B1(n_475),
.B2(n_478),
.C(n_479),
.Y(n_2558)
);

AOI21xp33_ASAP7_75t_L g2559 ( 
.A1(n_2558),
.A2(n_482),
.B(n_486),
.Y(n_2559)
);

AOI211xp5_ASAP7_75t_L g2560 ( 
.A1(n_2559),
.A2(n_488),
.B(n_491),
.C(n_492),
.Y(n_2560)
);


endmodule