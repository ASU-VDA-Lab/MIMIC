module fake_netlist_6_2144_n_1755 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1755);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1755;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_61),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_84),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_69),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_5),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_35),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_105),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_125),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_64),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_98),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_18),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_75),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_24),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_94),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_26),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_43),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_17),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_143),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_81),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_66),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_117),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_104),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_41),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_133),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_169),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_124),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_58),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_53),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_130),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_107),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_118),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_142),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_90),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_68),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_74),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_172),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_147),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_33),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_37),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_29),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_165),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_162),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_57),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_95),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_157),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_145),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_34),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_176),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_85),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_45),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_144),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_178),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_137),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_139),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_4),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_67),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_88),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_76),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_72),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_79),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_114),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_99),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_62),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_103),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_115),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_89),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_92),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_80),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_56),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_33),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_159),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_21),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_5),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_49),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_152),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_58),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_170),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_38),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_59),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_17),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_44),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_113),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_146),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_60),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_96),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_111),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_100),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_86),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_93),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_50),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_148),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_65),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_20),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_28),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_56),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_97),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_25),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_29),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_18),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_59),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_163),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_87),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_168),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_110),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_155),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_52),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_21),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_36),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_134),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_3),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_173),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_15),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_38),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_164),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_106),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_32),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_19),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_13),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_36),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_120),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_46),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_32),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_10),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_112),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_70),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_158),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_16),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_0),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_131),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_177),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_48),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_27),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_6),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_47),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_31),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_27),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_41),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_192),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_217),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_276),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_188),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_183),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_238),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_0),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_213),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_184),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_213),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_238),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_213),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_186),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_238),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_213),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_213),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_236),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_213),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_236),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_261),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_213),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_214),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_216),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_195),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_195),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_298),
.B(n_1),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_185),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_222),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_207),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_229),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_231),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_261),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_251),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_285),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_2),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_201),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_191),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_207),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_228),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_192),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_228),
.B(n_2),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_234),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_235),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_247),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_239),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_247),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_240),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_285),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_286),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_326),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_201),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_194),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_283),
.B(n_3),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_243),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_201),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_189),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_326),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_209),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_280),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_280),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_328),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_206),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_328),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_283),
.B(n_4),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_244),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_226),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_197),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_189),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_245),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_232),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_233),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_227),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_248),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_246),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_262),
.B(n_6),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_197),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_279),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_250),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_254),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_256),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_255),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_227),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_263),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_262),
.B(n_11),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_319),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_201),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_287),
.B(n_13),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_442),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_R g456 ( 
.A(n_443),
.B(n_264),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_366),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_370),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_374),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_377),
.B(n_319),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_384),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_237),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_418),
.B(n_287),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_379),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_418),
.B(n_314),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_385),
.B(n_182),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_376),
.A2(n_314),
.B(n_202),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_363),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_390),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_392),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_378),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g476 ( 
.A(n_415),
.B(n_252),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_378),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_393),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_404),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_418),
.B(n_190),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_381),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_380),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_383),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_437),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_405),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_208),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_407),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_431),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_382),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_409),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_451),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_R g497 ( 
.A(n_416),
.B(n_193),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_428),
.B(n_265),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_436),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_211),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_434),
.B(n_266),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_439),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_444),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_446),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_451),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_436),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_395),
.B(n_218),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_372),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_363),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_364),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_362),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_394),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_398),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_365),
.B(n_411),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_427),
.B(n_230),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_445),
.B(n_237),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_364),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_449),
.B(n_219),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_389),
.B(n_225),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_396),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_386),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_273),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_464),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_464),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_515),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_490),
.A2(n_440),
.B1(n_452),
.B2(n_397),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_386),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_490),
.B(n_241),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_490),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_517),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_267),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_454),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_512),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_501),
.A2(n_449),
.B1(n_368),
.B2(n_388),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_461),
.B(n_402),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_512),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_501),
.B(n_271),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_478),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_481),
.B(n_465),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_495),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_501),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_512),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_521),
.B(n_253),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_484),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_486),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_496),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_469),
.B(n_272),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_508),
.B(n_201),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_458),
.B(n_432),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

INVx4_ASAP7_75t_SL g562 ( 
.A(n_512),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_458),
.B(n_459),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_459),
.B(n_441),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_512),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_457),
.B(n_277),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_462),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_496),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_L g571 ( 
.A(n_462),
.B(n_201),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_481),
.B(n_368),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_465),
.B(n_282),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_471),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_466),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_476),
.A2(n_388),
.B1(n_403),
.B2(n_288),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_471),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_475),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_521),
.B(n_465),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_513),
.B(n_425),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_475),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_506),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_525),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_467),
.B(n_399),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_506),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_467),
.B(n_284),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_460),
.B(n_375),
.Y(n_590)
);

AO22x2_ASAP7_75t_L g591 ( 
.A1(n_521),
.A2(n_320),
.B1(n_331),
.B2(n_358),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_467),
.B(n_297),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_460),
.B(n_463),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_456),
.B(n_463),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_477),
.B(n_258),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_462),
.B(n_299),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_506),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_523),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_509),
.B(n_414),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_522),
.B(n_420),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_483),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_487),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_473),
.B(n_259),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_472),
.B(n_268),
.Y(n_606)
);

INVx4_ASAP7_75t_SL g607 ( 
.A(n_488),
.Y(n_607)
);

AND2x2_ASAP7_75t_SL g608 ( 
.A(n_470),
.B(n_278),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_499),
.B(n_502),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_473),
.B(n_289),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_474),
.B(n_252),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_474),
.B(n_410),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_479),
.B(n_293),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_470),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_470),
.Y(n_616)
);

OAI221xp5_ASAP7_75t_L g617 ( 
.A1(n_500),
.A2(n_403),
.B1(n_294),
.B2(n_357),
.C(n_352),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_470),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_498),
.A2(n_292),
.B1(n_347),
.B2(n_343),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_479),
.B(n_305),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_525),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_507),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_509),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_500),
.B(n_448),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_468),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_516),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_480),
.B(n_308),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_526),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_480),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_489),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_489),
.B(n_306),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_455),
.B(n_429),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_491),
.B(n_429),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_491),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_494),
.B(n_307),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_494),
.Y(n_639)
);

BUFx10_ASAP7_75t_L g640 ( 
.A(n_503),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_503),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_497),
.A2(n_210),
.B1(n_205),
.B2(n_203),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_504),
.A2(n_274),
.B1(n_304),
.B2(n_303),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_504),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_505),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_505),
.B(n_387),
.Y(n_646)
);

NOR2x1p5_ASAP7_75t_L g647 ( 
.A(n_510),
.B(n_204),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_510),
.B(n_312),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_511),
.B(n_387),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_511),
.A2(n_302),
.B1(n_317),
.B2(n_334),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_520),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_520),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_514),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_493),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_495),
.B(n_391),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_456),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_519),
.B(n_391),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_453),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_515),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_453),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_470),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_518),
.A2(n_296),
.B1(n_327),
.B2(n_315),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_515),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_453),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_515),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_518),
.B(n_309),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_518),
.B(n_310),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_604),
.Y(n_669)
);

BUFx6f_ASAP7_75t_SL g670 ( 
.A(n_640),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_616),
.B(n_220),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_536),
.B(n_325),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_552),
.B(n_530),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_657),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_530),
.B(n_344),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_L g676 ( 
.A(n_609),
.B(n_311),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_552),
.B(n_220),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_536),
.B(n_350),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_616),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_615),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_627),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_549),
.B(n_528),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_608),
.A2(n_223),
.B1(n_220),
.B2(n_353),
.Y(n_683)
);

AO22x1_ASAP7_75t_L g684 ( 
.A1(n_543),
.A2(n_345),
.B1(n_346),
.B2(n_355),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_531),
.B(n_412),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_533),
.B(n_275),
.C(n_270),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_549),
.B(n_324),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_531),
.B(n_332),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_532),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_608),
.A2(n_220),
.B1(n_223),
.B2(n_353),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_542),
.B(n_335),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_554),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_561),
.Y(n_693)
);

BUFx8_ASAP7_75t_L g694 ( 
.A(n_633),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_667),
.A2(n_426),
.B1(n_424),
.B2(n_419),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_660),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_631),
.B(n_338),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_660),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_611),
.B(n_413),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_547),
.B(n_400),
.Y(n_700)
);

BUFx8_ASAP7_75t_L g701 ( 
.A(n_633),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_668),
.B(n_614),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_547),
.B(n_400),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_664),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_547),
.A2(n_339),
.B1(n_203),
.B2(n_200),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_629),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_664),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_529),
.B(n_220),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_662),
.B(n_618),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_538),
.B(n_220),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_629),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_623),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_560),
.B(n_301),
.C(n_215),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_659),
.B(n_220),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_580),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_662),
.B(n_223),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_623),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_618),
.B(n_223),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_625),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_661),
.B(n_223),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_561),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_665),
.B(n_223),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_666),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_662),
.B(n_223),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_666),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_537),
.B(n_193),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_625),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_651),
.B(n_196),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_537),
.B(n_196),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_540),
.B(n_353),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_580),
.A2(n_353),
.B1(n_417),
.B2(n_237),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_636),
.B(n_353),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_636),
.B(n_353),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_580),
.Y(n_734)
);

AND2x2_ASAP7_75t_SL g735 ( 
.A(n_606),
.B(n_401),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_603),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_603),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_646),
.B(n_353),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_602),
.A2(n_342),
.B1(n_341),
.B2(n_290),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_556),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_646),
.B(n_198),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_625),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_553),
.B(n_198),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_624),
.B(n_401),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_557),
.B(n_199),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_596),
.A2(n_348),
.B(n_200),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_642),
.B(n_199),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_624),
.B(n_423),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_555),
.B(n_205),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_566),
.B(n_210),
.Y(n_750)
);

NOR2x1p5_ASAP7_75t_L g751 ( 
.A(n_599),
.B(n_204),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_575),
.Y(n_752)
);

BUFx12f_ASAP7_75t_SL g753 ( 
.A(n_651),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_572),
.B(n_406),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_572),
.A2(n_348),
.B1(n_349),
.B2(n_341),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_567),
.A2(n_349),
.B(n_422),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_572),
.A2(n_342),
.B1(n_187),
.B2(n_323),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_546),
.Y(n_758)
);

BUFx6f_ASAP7_75t_SL g759 ( 
.A(n_640),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_527),
.B(n_423),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_556),
.Y(n_761)
);

O2A1O1Ixp5_ASAP7_75t_L g762 ( 
.A1(n_545),
.A2(n_422),
.B(n_421),
.C(n_408),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_527),
.B(n_221),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_575),
.Y(n_764)
);

AOI22x1_ASAP7_75t_L g765 ( 
.A1(n_534),
.A2(n_290),
.B1(n_291),
.B2(n_345),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_546),
.B(n_224),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_569),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_534),
.B(n_421),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_606),
.B(n_242),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_658),
.B(n_249),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_658),
.B(n_406),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_539),
.B(n_257),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_574),
.B(n_260),
.Y(n_774)
);

AND2x6_ASAP7_75t_SL g775 ( 
.A(n_612),
.B(n_408),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_599),
.B(n_291),
.Y(n_776)
);

BUFx5_ASAP7_75t_L g777 ( 
.A(n_535),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_578),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_569),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_535),
.B(n_269),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_635),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_535),
.B(n_281),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_535),
.B(n_295),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_579),
.B(n_300),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_577),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_577),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_548),
.B(n_313),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_582),
.B(n_316),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_653),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_544),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_635),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_649),
.B(n_336),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_653),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_535),
.B(n_337),
.Y(n_794)
);

AND2x6_ASAP7_75t_SL g795 ( 
.A(n_590),
.B(n_564),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_535),
.B(n_333),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_589),
.B(n_340),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_572),
.A2(n_330),
.B1(n_359),
.B2(n_321),
.Y(n_798)
);

AO221x1_ASAP7_75t_L g799 ( 
.A1(n_591),
.A2(n_360),
.B1(n_356),
.B2(n_355),
.C(n_346),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_583),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_544),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_550),
.B(n_329),
.Y(n_802)
);

O2A1O1Ixp5_ASAP7_75t_L g803 ( 
.A1(n_573),
.A2(n_322),
.B(n_318),
.C(n_360),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_653),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_663),
.A2(n_356),
.B1(n_180),
.B2(n_179),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_587),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_656),
.B(n_22),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_570),
.B(n_174),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_654),
.Y(n_810)
);

INVxp33_ASAP7_75t_SL g811 ( 
.A(n_563),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_656),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_570),
.B(n_167),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_586),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_SL g815 ( 
.A1(n_655),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_601),
.B(n_166),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_588),
.A2(n_154),
.B(n_153),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_632),
.B(n_23),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_673),
.A2(n_559),
.B(n_605),
.C(n_610),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_682),
.B(n_634),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_768),
.B(n_651),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_789),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_685),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_747),
.A2(n_576),
.B(n_592),
.C(n_632),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_702),
.A2(n_551),
.B(n_568),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_673),
.A2(n_628),
.B(n_621),
.C(n_613),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_732),
.A2(n_628),
.B(n_621),
.C(n_613),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_679),
.A2(n_610),
.B(n_605),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_805),
.A2(n_639),
.B1(n_593),
.B2(n_644),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_699),
.B(n_639),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_671),
.A2(n_598),
.B(n_600),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_679),
.B(n_638),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_726),
.A2(n_643),
.B(n_650),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_732),
.A2(n_648),
.B(n_617),
.C(n_602),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_718),
.A2(n_598),
.B(n_600),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_733),
.A2(n_738),
.B(n_677),
.C(n_763),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_719),
.A2(n_645),
.B(n_637),
.C(n_641),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_718),
.A2(n_600),
.B(n_541),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_734),
.A2(n_652),
.B1(n_594),
.B2(n_602),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_744),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_758),
.B(n_586),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_716),
.A2(n_541),
.B(n_584),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_716),
.A2(n_541),
.B(n_584),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_724),
.A2(n_541),
.B(n_584),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_699),
.B(n_640),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_733),
.A2(n_738),
.B(n_677),
.C(n_771),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_715),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_693),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_811),
.B(n_585),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_781),
.Y(n_850)
);

OAI321xp33_ASAP7_75t_L g851 ( 
.A1(n_815),
.A2(n_648),
.A3(n_602),
.B1(n_620),
.B2(n_594),
.C(n_586),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_734),
.A2(n_652),
.B1(n_586),
.B2(n_558),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_693),
.Y(n_853)
);

OAI21xp33_ASAP7_75t_L g854 ( 
.A1(n_729),
.A2(n_591),
.B(n_622),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_679),
.A2(n_541),
.B(n_565),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_789),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_715),
.A2(n_565),
.B(n_584),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_735),
.B(n_654),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_721),
.A2(n_715),
.B1(n_727),
.B2(n_742),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_735),
.A2(n_647),
.B1(n_601),
.B2(n_595),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_811),
.B(n_630),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_736),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_793),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_810),
.Y(n_864)
);

OR2x6_ASAP7_75t_SL g865 ( 
.A(n_752),
.B(n_674),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_736),
.B(n_597),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_737),
.B(n_597),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_L g868 ( 
.A1(n_787),
.A2(n_792),
.B(n_812),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_700),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_791),
.B(n_764),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_793),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_791),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_812),
.A2(n_591),
.B1(n_619),
.B2(n_626),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_752),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_695),
.B(n_571),
.C(n_607),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_803),
.A2(n_595),
.B(n_562),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_802),
.A2(n_562),
.B(n_595),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_777),
.B(n_595),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_760),
.B(n_562),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_686),
.A2(n_595),
.B(n_28),
.C(n_30),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_687),
.A2(n_595),
.B(n_151),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_773),
.A2(n_136),
.B1(n_135),
.B2(n_132),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_795),
.B(n_770),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_804),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_672),
.A2(n_129),
.B(n_127),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_770),
.B(n_26),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_706),
.A2(n_31),
.B(n_34),
.C(n_35),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_678),
.A2(n_126),
.B(n_123),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_741),
.B(n_37),
.C(n_39),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_748),
.B(n_40),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_L g891 ( 
.A(n_674),
.B(n_122),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_703),
.A2(n_102),
.B(n_101),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_804),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_769),
.B(n_772),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_790),
.A2(n_83),
.B(n_82),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_712),
.B(n_71),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_711),
.B(n_42),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_790),
.A2(n_46),
.B(n_47),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_745),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_762),
.A2(n_54),
.B(n_55),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_669),
.B(n_54),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_755),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_683),
.A2(n_690),
.B(n_707),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_801),
.A2(n_697),
.B(n_796),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_780),
.A2(n_783),
.B(n_782),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_745),
.A2(n_750),
.B(n_806),
.C(n_784),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_670),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_794),
.A2(n_688),
.B(n_730),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_754),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_818),
.A2(n_691),
.B(n_680),
.C(n_681),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_740),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_717),
.B(n_728),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_740),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_754),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_708),
.A2(n_720),
.B(n_722),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_L g916 ( 
.A(n_684),
.B(n_739),
.C(n_713),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_675),
.A2(n_731),
.B1(n_754),
.B2(n_705),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_676),
.B(n_757),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_798),
.B(n_776),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_808),
.B(n_773),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_670),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_778),
.B(n_707),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_710),
.A2(n_714),
.B(n_816),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_753),
.B(n_766),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_761),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_809),
.A2(n_813),
.B(n_807),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_750),
.A2(n_797),
.B(n_784),
.C(n_774),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_761),
.A2(n_767),
.B(n_807),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_774),
.A2(n_788),
.B(n_797),
.C(n_675),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_814),
.B(n_754),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_767),
.A2(n_779),
.B(n_785),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_689),
.A2(n_704),
.B(n_725),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_SL g933 ( 
.A(n_753),
.B(n_670),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_675),
.A2(n_751),
.B1(n_788),
.B2(n_766),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_779),
.A2(n_785),
.B(n_786),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_786),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_675),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_800),
.A2(n_692),
.B(n_723),
.Y(n_938)
);

AOI33xp33_ASAP7_75t_L g939 ( 
.A1(n_799),
.A2(n_765),
.A3(n_775),
.B1(n_698),
.B2(n_696),
.B3(n_704),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_800),
.A2(n_723),
.B(n_749),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_743),
.Y(n_941)
);

OR2x6_ASAP7_75t_SL g942 ( 
.A(n_694),
.B(n_701),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_756),
.A2(n_746),
.B1(n_817),
.B2(n_759),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_694),
.B(n_701),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_777),
.A2(n_759),
.B(n_810),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_810),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_777),
.A2(n_673),
.B(n_733),
.C(n_732),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_777),
.B(n_715),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_682),
.B(n_528),
.Y(n_951)
);

AO32x2_ASAP7_75t_L g952 ( 
.A1(n_815),
.A2(n_812),
.A3(n_806),
.B1(n_536),
.B2(n_549),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_699),
.B(n_530),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_726),
.A2(n_518),
.B(n_528),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_721),
.Y(n_955)
);

NAND2x1_ASAP7_75t_L g956 ( 
.A(n_715),
.B(n_679),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_700),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_682),
.B(n_528),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_709),
.A2(n_662),
.B(n_614),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_673),
.A2(n_732),
.B(n_738),
.C(n_733),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_747),
.A2(n_528),
.B(n_518),
.C(n_682),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_702),
.A2(n_734),
.B1(n_682),
.B2(n_549),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_951),
.B(n_961),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_840),
.B(n_823),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_894),
.B(n_820),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_955),
.Y(n_970)
);

INVx5_ASAP7_75t_L g971 ( 
.A(n_847),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_965),
.B(n_954),
.Y(n_972)
);

AOI211x1_ASAP7_75t_L g973 ( 
.A1(n_854),
.A2(n_833),
.B(n_828),
.C(n_900),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_903),
.A2(n_958),
.B(n_950),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_823),
.B(n_849),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_903),
.A2(n_962),
.B(n_959),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_922),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_827),
.A2(n_826),
.B(n_902),
.C(n_906),
.Y(n_978)
);

AO31x2_ASAP7_75t_L g979 ( 
.A1(n_910),
.A2(n_966),
.A3(n_873),
.B(n_852),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_868),
.B(n_941),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_886),
.A2(n_824),
.B1(n_917),
.B2(n_934),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_918),
.A2(n_905),
.B(n_943),
.C(n_908),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_850),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_872),
.B(n_858),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_832),
.B(n_828),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_864),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_830),
.B(n_953),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_851),
.B(n_829),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_955),
.B(n_960),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_960),
.B(n_963),
.Y(n_990)
);

AOI21x1_ASAP7_75t_L g991 ( 
.A1(n_825),
.A2(n_904),
.B(n_926),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_847),
.B(n_869),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_963),
.B(n_890),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_923),
.A2(n_835),
.B(n_831),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_878),
.A2(n_846),
.B(n_836),
.Y(n_995)
);

AND3x4_ASAP7_75t_L g996 ( 
.A(n_919),
.B(n_916),
.C(n_821),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_841),
.B(n_870),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_869),
.B(n_862),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_920),
.A2(n_859),
.B(n_838),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_863),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_947),
.A2(n_964),
.B(n_915),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_956),
.A2(n_948),
.B(n_879),
.Y(n_1002)
);

AOI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_819),
.A2(n_834),
.B(n_851),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_863),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_870),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_938),
.A2(n_940),
.B(n_932),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_866),
.A2(n_867),
.B(n_935),
.Y(n_1007)
);

CKINVDCx8_ASAP7_75t_R g1008 ( 
.A(n_874),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_870),
.B(n_839),
.Y(n_1009)
);

OAI22x1_ASAP7_75t_L g1010 ( 
.A1(n_883),
.A2(n_946),
.B1(n_930),
.B2(n_845),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_928),
.A2(n_931),
.B(n_877),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_841),
.B(n_822),
.Y(n_1012)
);

BUFx12f_ASAP7_75t_L g1013 ( 
.A(n_907),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_909),
.Y(n_1014)
);

CKINVDCx8_ASAP7_75t_R g1015 ( 
.A(n_921),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_909),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_857),
.A2(n_855),
.B(n_844),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_929),
.A2(n_927),
.B(n_837),
.C(n_939),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_842),
.A2(n_843),
.B(n_912),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_937),
.B(n_848),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_876),
.A2(n_860),
.B(n_936),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_909),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_SL g1023 ( 
.A1(n_889),
.A2(n_882),
.B(n_899),
.Y(n_1023)
);

NAND2xp33_ASAP7_75t_L g1024 ( 
.A(n_937),
.B(n_893),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_863),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_930),
.B(n_856),
.Y(n_1026)
);

AO31x2_ASAP7_75t_L g1027 ( 
.A1(n_880),
.A2(n_897),
.A3(n_887),
.B(n_881),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_848),
.B(n_853),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_924),
.B(n_848),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_911),
.A2(n_925),
.B(n_900),
.Y(n_1031)
);

AO21x1_ASAP7_75t_L g1032 ( 
.A1(n_898),
.A2(n_892),
.B(n_901),
.Y(n_1032)
);

INVx6_ASAP7_75t_L g1033 ( 
.A(n_893),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_853),
.B(n_957),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_853),
.B(n_914),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_895),
.A2(n_888),
.B(n_885),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_871),
.B(n_884),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_871),
.B(n_884),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_937),
.B(n_896),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_944),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_914),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_875),
.A2(n_861),
.B(n_945),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_891),
.A2(n_933),
.B(n_952),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_933),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_942),
.B(n_865),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_952),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_952),
.A2(n_963),
.B(n_960),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_870),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_903),
.A2(n_950),
.B(n_949),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_849),
.B(n_811),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_847),
.A2(n_662),
.B(n_709),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_847),
.B(n_734),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_894),
.A2(n_965),
.B1(n_902),
.B2(n_833),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_870),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_903),
.A2(n_950),
.B(n_949),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_951),
.B(n_961),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_930),
.B(n_841),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_910),
.A2(n_966),
.A3(n_873),
.B(n_852),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_951),
.B(n_961),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_847),
.A2(n_662),
.B(n_709),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_849),
.B(n_811),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_951),
.B(n_961),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_870),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_902),
.A2(n_954),
.B1(n_919),
.B2(n_868),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_870),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_L g1066 ( 
.A(n_864),
.Y(n_1066)
);

NAND2x1_ASAP7_75t_L g1067 ( 
.A(n_955),
.B(n_715),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_840),
.B(n_805),
.Y(n_1068)
);

NAND2x1p5_ASAP7_75t_L g1069 ( 
.A(n_847),
.B(n_734),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_910),
.A2(n_966),
.A3(n_873),
.B(n_852),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_922),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_SL g1072 ( 
.A1(n_902),
.A2(n_381),
.B1(n_382),
.B2(n_379),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_910),
.A2(n_966),
.A3(n_873),
.B(n_852),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_847),
.A2(n_662),
.B(n_709),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_913),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_902),
.A2(n_954),
.B1(n_886),
.B2(n_916),
.Y(n_1076)
);

NAND3xp33_ASAP7_75t_SL g1077 ( 
.A(n_954),
.B(n_611),
.C(n_833),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_864),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_870),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_951),
.B(n_961),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_840),
.B(n_805),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_847),
.B(n_734),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_916),
.A2(n_886),
.B1(n_854),
.B2(n_954),
.C(n_873),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_847),
.A2(n_662),
.B(n_709),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_SL g1085 ( 
.A1(n_945),
.A2(n_964),
.B(n_947),
.Y(n_1085)
);

OA22x2_ASAP7_75t_L g1086 ( 
.A1(n_854),
.A2(n_799),
.B1(n_815),
.B2(n_833),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_903),
.A2(n_950),
.B(n_949),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_955),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_863),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_847),
.A2(n_662),
.B(n_709),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_913),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_870),
.Y(n_1092)
);

O2A1O1Ixp5_ASAP7_75t_L g1093 ( 
.A1(n_965),
.A2(n_918),
.B(n_905),
.C(n_943),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_894),
.B(n_699),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_903),
.A2(n_950),
.B(n_949),
.Y(n_1095)
);

INVx3_ASAP7_75t_SL g1096 ( 
.A(n_1078),
.Y(n_1096)
);

INVx3_ASAP7_75t_SL g1097 ( 
.A(n_1026),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_975),
.B(n_968),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1013),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1033),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1076),
.A2(n_1056),
.B(n_967),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_967),
.B(n_1056),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1008),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1059),
.B(n_1062),
.Y(n_1104)
);

NOR2x1p5_ASAP7_75t_L g1105 ( 
.A(n_1044),
.B(n_1045),
.Y(n_1105)
);

INVx6_ASAP7_75t_L g1106 ( 
.A(n_1040),
.Y(n_1106)
);

INVx8_ASAP7_75t_L g1107 ( 
.A(n_1016),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1059),
.B(n_1062),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1080),
.B(n_969),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1080),
.B(n_1030),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_981),
.A2(n_1077),
.B1(n_1053),
.B2(n_1086),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1068),
.B(n_1081),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1016),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_986),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1057),
.B(n_1029),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1026),
.Y(n_1117)
);

INVx3_ASAP7_75t_SL g1118 ( 
.A(n_1029),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_969),
.B(n_977),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_1012),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1001),
.A2(n_1093),
.B(n_978),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_SL g1122 ( 
.A(n_1079),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_997),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1071),
.B(n_1053),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1033),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1035),
.B(n_1034),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1050),
.B(n_1061),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1064),
.A2(n_1003),
.B(n_1023),
.C(n_972),
.Y(n_1128)
);

BUFx4_ASAP7_75t_SL g1129 ( 
.A(n_1054),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_980),
.B1(n_984),
.B2(n_1044),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1075),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_972),
.B(n_985),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1035),
.B(n_1005),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1014),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_974),
.A2(n_1095),
.B(n_1055),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_985),
.B(n_973),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1094),
.B(n_987),
.Y(n_1137)
);

OAI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_1086),
.A2(n_1023),
.B(n_1003),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1065),
.B(n_1092),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_987),
.B(n_993),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1091),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_983),
.B(n_1072),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1048),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_970),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_L g1145 ( 
.A(n_1016),
.B(n_1022),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_974),
.A2(n_1087),
.B(n_976),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1018),
.A2(n_1009),
.B(n_1063),
.C(n_1043),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1028),
.B(n_1037),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1016),
.B(n_1022),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1028),
.B(n_1020),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1038),
.B(n_1014),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1010),
.B(n_1004),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1004),
.B(n_1025),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1004),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_993),
.A2(n_990),
.B1(n_1046),
.B2(n_1047),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_976),
.A2(n_1087),
.B(n_1049),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1083),
.B(n_990),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1025),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_989),
.B(n_970),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1015),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1085),
.A2(n_1032),
.B1(n_1041),
.B2(n_1088),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_989),
.B(n_1088),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1049),
.A2(n_1042),
.B1(n_1021),
.B2(n_1000),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1000),
.B(n_1089),
.Y(n_1165)
);

AO21x1_ASAP7_75t_L g1166 ( 
.A1(n_1042),
.A2(n_1021),
.B(n_1031),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_R g1167 ( 
.A(n_1022),
.B(n_1089),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1025),
.B(n_1022),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1031),
.B(n_979),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_979),
.B(n_1070),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_1024),
.Y(n_1171)
);

OAI321xp33_ASAP7_75t_L g1172 ( 
.A1(n_1045),
.A2(n_1006),
.A3(n_999),
.B1(n_991),
.B2(n_1007),
.C(n_994),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1066),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_992),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1066),
.B(n_1027),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1027),
.B(n_979),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_992),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1027),
.B(n_1058),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1052),
.B(n_1082),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_1052),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1069),
.A2(n_1060),
.B1(n_1084),
.B2(n_1074),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1067),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1058),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1019),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1073),
.B(n_1011),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1051),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1090),
.A2(n_1002),
.B(n_1073),
.C(n_1036),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1017),
.B(n_975),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_SL g1189 ( 
.A1(n_1050),
.A2(n_811),
.B1(n_1061),
.B2(n_381),
.Y(n_1189)
);

AOI21xp33_ASAP7_75t_L g1190 ( 
.A1(n_981),
.A2(n_988),
.B(n_1076),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1013),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_988),
.A2(n_902),
.B1(n_916),
.B2(n_886),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_967),
.A2(n_1056),
.B1(n_1062),
.B2(n_1059),
.Y(n_1193)
);

NAND2x1p5_ASAP7_75t_L g1194 ( 
.A(n_971),
.B(n_1016),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_992),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_974),
.A2(n_1049),
.B(n_976),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_967),
.B(n_1056),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1014),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_967),
.B(n_1056),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_L g1202 ( 
.A1(n_981),
.A2(n_1093),
.B(n_1003),
.C(n_988),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_967),
.B(n_1056),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1013),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_968),
.Y(n_1205)
);

INVx3_ASAP7_75t_SL g1206 ( 
.A(n_1078),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1014),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_975),
.B(n_805),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_967),
.B(n_633),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_967),
.B(n_1056),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_967),
.B(n_1056),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_988),
.A2(n_902),
.B1(n_916),
.B2(n_886),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_988),
.A2(n_902),
.B1(n_916),
.B2(n_886),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_986),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_982),
.A2(n_995),
.B(n_1001),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_1008),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_988),
.A2(n_560),
.B(n_564),
.C(n_883),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_975),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1014),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1014),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_967),
.B(n_1056),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_975),
.B(n_805),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_968),
.Y(n_1225)
);

OR2x6_ASAP7_75t_L g1226 ( 
.A(n_1054),
.B(n_870),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1215),
.A2(n_1121),
.B(n_1202),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1112),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1110),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1183),
.Y(n_1231)
);

BUFx2_ASAP7_75t_R g1232 ( 
.A(n_1096),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1131),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1150),
.B(n_1113),
.Y(n_1234)
);

INVx11_ASAP7_75t_L g1235 ( 
.A(n_1115),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1098),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1150),
.B(n_1113),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1107),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1108),
.A2(n_1201),
.B1(n_1222),
.B2(n_1198),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1097),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1190),
.A2(n_1213),
.B1(n_1192),
.B2(n_1212),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1102),
.B(n_1109),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1108),
.B(n_1198),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1216),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1123),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1146),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1201),
.A2(n_1203),
.B1(n_1211),
.B2(n_1210),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1190),
.A2(n_1138),
.B1(n_1111),
.B2(n_1101),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_SL g1249 ( 
.A(n_1214),
.B(n_1106),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1134),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1189),
.A2(n_1127),
.B1(n_1130),
.B2(n_1142),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1215),
.A2(n_1121),
.B(n_1172),
.Y(n_1252)
);

AO21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1124),
.A2(n_1170),
.B(n_1169),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1203),
.B(n_1210),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1188),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1119),
.Y(n_1256)
);

INVx4_ASAP7_75t_SL g1257 ( 
.A(n_1134),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1211),
.A2(n_1222),
.B1(n_1104),
.B2(n_1193),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1119),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1218),
.B(n_1208),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1160),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1184),
.A2(n_1175),
.B1(n_1171),
.B2(n_1106),
.Y(n_1262)
);

CKINVDCx14_ASAP7_75t_R g1263 ( 
.A(n_1099),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1154),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1160),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1151),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1163),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1163),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1205),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1166),
.A2(n_1147),
.B1(n_1157),
.B2(n_1135),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1223),
.B(n_1225),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1140),
.B(n_1137),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1206),
.Y(n_1273)
);

AO21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1170),
.A2(n_1169),
.B(n_1158),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1144),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1209),
.B(n_1120),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1137),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1107),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1107),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1148),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1226),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1136),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1136),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1149),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1135),
.A2(n_1157),
.B1(n_1197),
.B2(n_1164),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1178),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1134),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1129),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1153),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1105),
.A2(n_1126),
.B1(n_1200),
.B2(n_1195),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1140),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1180),
.B(n_1174),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1103),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1152),
.A2(n_1122),
.B1(n_1217),
.B2(n_1227),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1176),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1126),
.B(n_1227),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1194),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1132),
.Y(n_1298)
);

BUFx5_ASAP7_75t_L g1299 ( 
.A(n_1185),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1132),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_SL g1301 ( 
.A(n_1161),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1158),
.A2(n_1143),
.B1(n_1226),
.B2(n_1139),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1139),
.Y(n_1303)
);

CKINVDCx14_ASAP7_75t_R g1304 ( 
.A(n_1191),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1226),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1177),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1133),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1133),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1172),
.A2(n_1187),
.B(n_1181),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1128),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1162),
.A2(n_1118),
.B1(n_1117),
.B2(n_1174),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1114),
.B(n_1224),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1122),
.A2(n_1156),
.B1(n_1221),
.B2(n_1114),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1168),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1195),
.A2(n_1224),
.B1(n_1221),
.B2(n_1200),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1204),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1199),
.A2(n_1220),
.B1(n_1219),
.B2(n_1207),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1194),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1159),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1155),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1173),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1116),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1199),
.B(n_1220),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1207),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1219),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1219),
.A2(n_1220),
.B1(n_1145),
.B2(n_1180),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1156),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1100),
.B(n_1125),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1186),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1196),
.A2(n_1179),
.B1(n_1165),
.B2(n_1180),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1196),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1167),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1182),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1182),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1150),
.B(n_971),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1141),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1112),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1189),
.A2(n_611),
.B1(n_379),
.B2(n_382),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1216),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1183),
.Y(n_1340)
);

BUFx8_ASAP7_75t_L g1341 ( 
.A(n_1115),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1141),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1115),
.Y(n_1343)
);

OAI22x1_ASAP7_75t_L g1344 ( 
.A1(n_1130),
.A2(n_988),
.B1(n_996),
.B2(n_1064),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1107),
.Y(n_1345)
);

INVx2_ASAP7_75t_R g1346 ( 
.A(n_1327),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1251),
.B(n_1293),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1329),
.B(n_1255),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1255),
.B(n_1295),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1253),
.B(n_1274),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1286),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1231),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1270),
.B(n_1261),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1281),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1231),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1286),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1229),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1340),
.Y(n_1358)
);

NAND2x1_ASAP7_75t_L g1359 ( 
.A(n_1329),
.B(n_1280),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1340),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1269),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1299),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_SL g1363 ( 
.A(n_1232),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1228),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1265),
.B(n_1268),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1228),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1228),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1241),
.A2(n_1344),
.B1(n_1310),
.B2(n_1248),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1285),
.B(n_1267),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1337),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1241),
.A2(n_1248),
.B1(n_1338),
.B2(n_1262),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1305),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1285),
.B(n_1277),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1313),
.A2(n_1283),
.B(n_1282),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1299),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1294),
.A2(n_1302),
.B1(n_1313),
.B2(n_1236),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1252),
.A2(n_1332),
.B(n_1246),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1299),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1299),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1299),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1302),
.A2(n_1300),
.B(n_1298),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1292),
.B(n_1311),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1292),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1266),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1296),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1242),
.B(n_1243),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1244),
.B(n_1312),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1230),
.B(n_1289),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1258),
.B(n_1272),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1309),
.A2(n_1239),
.B(n_1247),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1334),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1345),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1276),
.A2(n_1239),
.B(n_1330),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1245),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1276),
.A2(n_1301),
.B1(n_1322),
.B2(n_1307),
.Y(n_1396)
);

CKINVDCx16_ASAP7_75t_R g1397 ( 
.A(n_1301),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1271),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1291),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1319),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1336),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1342),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1256),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1259),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1254),
.A2(n_1331),
.B(n_1306),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1284),
.B(n_1296),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1264),
.B(n_1275),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1314),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1233),
.B(n_1260),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1308),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1333),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1303),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1297),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1318),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1320),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1240),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1296),
.B(n_1290),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1379),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1346),
.B(n_1323),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1379),
.B(n_1380),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1379),
.B(n_1326),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1372),
.A2(n_1315),
.B1(n_1321),
.B2(n_1320),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1359),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1351),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1380),
.B(n_1325),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1356),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1368),
.A2(n_1249),
.B1(n_1273),
.B2(n_1240),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1362),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1356),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1430)
);

NAND4xp25_ASAP7_75t_L g1431 ( 
.A(n_1347),
.B(n_1328),
.C(n_1317),
.D(n_1250),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1394),
.B(n_1273),
.C(n_1244),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1378),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1390),
.A2(n_1321),
.B1(n_1343),
.B2(n_1324),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1391),
.A2(n_1341),
.B1(n_1304),
.B2(n_1263),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1384),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1352),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1390),
.B(n_1353),
.Y(n_1438)
);

NOR2x1_ASAP7_75t_L g1439 ( 
.A(n_1405),
.B(n_1278),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1377),
.A2(n_1335),
.B(n_1237),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1364),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1366),
.B(n_1287),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1383),
.B(n_1345),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1353),
.B(n_1234),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1376),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1366),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1374),
.B(n_1257),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_L g1449 ( 
.A(n_1392),
.B(n_1238),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1348),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1374),
.B(n_1257),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1398),
.A2(n_1343),
.B1(n_1324),
.B2(n_1304),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1370),
.B(n_1279),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1435),
.B(n_1384),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1450),
.B(n_1370),
.Y(n_1455)
);

NOR3xp33_ASAP7_75t_L g1456 ( 
.A(n_1432),
.B(n_1397),
.C(n_1388),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1450),
.B(n_1350),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1438),
.B(n_1385),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1444),
.A2(n_1383),
.B(n_1392),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1438),
.B(n_1361),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1422),
.A2(n_1383),
.B1(n_1397),
.B2(n_1415),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1435),
.B(n_1396),
.C(n_1387),
.Y(n_1462)
);

OAI21xp33_ASAP7_75t_L g1463 ( 
.A1(n_1422),
.A2(n_1427),
.B(n_1432),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1427),
.A2(n_1383),
.B1(n_1371),
.B2(n_1357),
.C(n_1415),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1430),
.B(n_1349),
.Y(n_1465)
);

OAI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1434),
.A2(n_1416),
.B1(n_1373),
.B2(n_1354),
.C(n_1383),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1434),
.A2(n_1417),
.B1(n_1409),
.B2(n_1354),
.C(n_1373),
.Y(n_1467)
);

NAND4xp25_ASAP7_75t_L g1468 ( 
.A(n_1452),
.B(n_1409),
.C(n_1389),
.D(n_1407),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1440),
.B(n_1375),
.C(n_1412),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1440),
.B(n_1431),
.C(n_1439),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1424),
.B(n_1395),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1452),
.A2(n_1417),
.B1(n_1389),
.B2(n_1412),
.C(n_1403),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1431),
.B(n_1375),
.C(n_1400),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1426),
.A2(n_1407),
.B1(n_1408),
.B2(n_1406),
.C(n_1403),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1426),
.B(n_1365),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1448),
.B(n_1363),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1442),
.A2(n_1367),
.B(n_1369),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1423),
.B(n_1384),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1448),
.B(n_1386),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1444),
.A2(n_1406),
.B1(n_1386),
.B2(n_1391),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1420),
.B(n_1348),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1451),
.B(n_1408),
.C(n_1411),
.D(n_1402),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1447),
.Y(n_1483)
);

NAND2x1_ASAP7_75t_L g1484 ( 
.A(n_1423),
.B(n_1355),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1420),
.B(n_1348),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1429),
.B(n_1365),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1429),
.B(n_1365),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1439),
.B(n_1375),
.C(n_1382),
.Y(n_1488)
);

NAND4xp25_ASAP7_75t_L g1489 ( 
.A(n_1419),
.B(n_1411),
.C(n_1401),
.D(n_1402),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1442),
.B(n_1382),
.C(n_1410),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1453),
.B(n_1365),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1420),
.B(n_1348),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1425),
.B(n_1404),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1418),
.B(n_1358),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1421),
.A2(n_1399),
.B(n_1406),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1421),
.B(n_1414),
.C(n_1413),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1444),
.A2(n_1406),
.B1(n_1386),
.B2(n_1399),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1421),
.B(n_1414),
.C(n_1413),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1425),
.B(n_1404),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1418),
.B(n_1360),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1477),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1483),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1483),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1494),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1477),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1494),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1500),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1500),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1455),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1493),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1460),
.B(n_1437),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1499),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1458),
.B(n_1428),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1485),
.B(n_1446),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1484),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1455),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1471),
.B(n_1443),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1465),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1492),
.B(n_1433),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1480),
.B(n_1457),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1488),
.B(n_1446),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1457),
.B(n_1433),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1491),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1475),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1487),
.B(n_1437),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1489),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1459),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1502),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

NOR2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1530),
.B(n_1468),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1530),
.B(n_1470),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1518),
.B(n_1459),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1527),
.B(n_1474),
.Y(n_1537)
);

NAND4xp25_ASAP7_75t_L g1538 ( 
.A(n_1523),
.B(n_1463),
.C(n_1456),
.D(n_1473),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1508),
.B(n_1454),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1508),
.B(n_1454),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1508),
.B(n_1479),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1517),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1524),
.B(n_1478),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1527),
.B(n_1495),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1517),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1504),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1524),
.B(n_1496),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1504),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1506),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1528),
.B(n_1482),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1506),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1507),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1529),
.B(n_1469),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1507),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1514),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1509),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1514),
.B(n_1436),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1516),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1512),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1509),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1511),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1511),
.B(n_1445),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1501),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1520),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1520),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1535),
.B(n_1341),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1534),
.A2(n_1464),
.B1(n_1467),
.B2(n_1472),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1546),
.B(n_1524),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1567),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1553),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1568),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1568),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1531),
.B(n_1521),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1526),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1569),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1567),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1556),
.Y(n_1582)
);

CKINVDCx16_ASAP7_75t_R g1583 ( 
.A(n_1531),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1569),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1563),
.B(n_1526),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1549),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1551),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1547),
.B(n_1526),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1536),
.B(n_1521),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1536),
.B(n_1525),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1539),
.B(n_1525),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1538),
.B(n_1513),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1539),
.B(n_1525),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1546),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1546),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1551),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1552),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1556),
.B(n_1515),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1561),
.B(n_1552),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1540),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1561),
.B(n_1515),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1542),
.B(n_1522),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1550),
.A2(n_1461),
.B(n_1462),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1554),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1540),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1542),
.B(n_1522),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1558),
.B(n_1522),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1555),
.Y(n_1611)
);

NAND2x1p5_ASAP7_75t_L g1612 ( 
.A(n_1550),
.B(n_1524),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1612),
.B(n_1558),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1582),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1584),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1596),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1612),
.B(n_1550),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1605),
.A2(n_1572),
.B1(n_1575),
.B2(n_1593),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1572),
.A2(n_1466),
.B1(n_1523),
.B2(n_1476),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1612),
.B(n_1562),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1583),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1582),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1574),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1576),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1574),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1573),
.B(n_1562),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1596),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1600),
.B(n_1541),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1576),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1571),
.B(n_1235),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1577),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1583),
.A2(n_1444),
.B1(n_1523),
.B2(n_1524),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1573),
.B(n_1505),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1574),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1581),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1596),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1577),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1600),
.B(n_1541),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1581),
.Y(n_1640)
);

INVx3_ASAP7_75t_SL g1641 ( 
.A(n_1597),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1580),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1596),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1581),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1591),
.B(n_1544),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1580),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1618),
.A2(n_1603),
.B(n_1597),
.C(n_1589),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1621),
.A2(n_1603),
.B1(n_1578),
.B2(n_1590),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1621),
.B(n_1570),
.C(n_1602),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1624),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.B(n_1595),
.Y(n_1653)
);

NOR2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1646),
.B(n_1578),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1619),
.A2(n_1601),
.B(n_1590),
.C(n_1608),
.Y(n_1655)
);

AND2x4_ASAP7_75t_SL g1656 ( 
.A(n_1617),
.B(n_1316),
.Y(n_1656)
);

OA22x2_ASAP7_75t_L g1657 ( 
.A1(n_1619),
.A2(n_1548),
.B1(n_1587),
.B2(n_1606),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1624),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1591),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1622),
.B(n_1586),
.Y(n_1660)
);

AOI222xp33_ASAP7_75t_L g1661 ( 
.A1(n_1622),
.A2(n_1615),
.B1(n_1646),
.B2(n_1617),
.C1(n_1632),
.C2(n_1641),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1628),
.B(n_1601),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1604),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1641),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_L g1666 ( 
.A(n_1617),
.B(n_1288),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1613),
.A2(n_1609),
.B1(n_1592),
.B2(n_1594),
.Y(n_1668)
);

NAND2x1_ASAP7_75t_L g1669 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1629),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1594),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1638),
.A2(n_1610),
.B1(n_1497),
.B2(n_1608),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1641),
.A2(n_1607),
.B1(n_1444),
.B2(n_1498),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1638),
.A2(n_1444),
.B1(n_1608),
.B2(n_1602),
.Y(n_1674)
);

OAI211xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1615),
.A2(n_1602),
.B(n_1587),
.C(n_1606),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1662),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1664),
.B(n_1645),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1664),
.B(n_1645),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1663),
.B(n_1645),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1652),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1627),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1659),
.B(n_1628),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1654),
.B(n_1661),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1649),
.B(n_1630),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1657),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1661),
.B(n_1636),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1660),
.B(n_1263),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1656),
.B(n_1636),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1658),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_SL g1691 ( 
.A(n_1655),
.B(n_1675),
.C(n_1673),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1653),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1636),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1657),
.A2(n_1666),
.B1(n_1667),
.B2(n_1665),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1613),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1616),
.Y(n_1696)
);

NAND3x2_ASAP7_75t_L g1697 ( 
.A(n_1683),
.B(n_1620),
.C(n_1628),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1689),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1677),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1691),
.B(n_1674),
.C(n_1669),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1684),
.A2(n_1620),
.B1(n_1648),
.B2(n_1642),
.C(n_1631),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_SL g1702 ( 
.A(n_1687),
.B(n_1672),
.C(n_1620),
.D(n_1639),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1691),
.A2(n_1626),
.B1(n_1633),
.B2(n_1643),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1686),
.A2(n_1643),
.B(n_1616),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_SL g1705 ( 
.A(n_1692),
.B(n_1339),
.C(n_1639),
.Y(n_1705)
);

AOI222xp33_ASAP7_75t_L g1706 ( 
.A1(n_1686),
.A2(n_1633),
.B1(n_1629),
.B2(n_1631),
.C1(n_1648),
.C2(n_1637),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1678),
.B(n_1616),
.Y(n_1707)
);

NAND2x2_ASAP7_75t_L g1708 ( 
.A(n_1682),
.B(n_1643),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1694),
.A2(n_1633),
.B1(n_1642),
.B2(n_1637),
.C(n_1626),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1676),
.B(n_1694),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1705),
.B(n_1685),
.C(n_1693),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1698),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1699),
.B(n_1679),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1707),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1710),
.A2(n_1688),
.B(n_1680),
.Y(n_1716)
);

OAI322xp33_ASAP7_75t_L g1717 ( 
.A1(n_1703),
.A2(n_1690),
.A3(n_1696),
.B1(n_1695),
.B2(n_1639),
.C1(n_1625),
.C2(n_1635),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_L g1718 ( 
.A(n_1704),
.B(n_1689),
.Y(n_1718)
);

NAND2x1_ASAP7_75t_SL g1719 ( 
.A(n_1708),
.B(n_1626),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1709),
.B(n_1633),
.C(n_1625),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1700),
.A2(n_1625),
.B(n_1623),
.Y(n_1721)
);

OAI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1712),
.A2(n_1702),
.B(n_1706),
.Y(n_1722)
);

NAND4xp25_ASAP7_75t_SL g1723 ( 
.A(n_1711),
.B(n_1701),
.C(n_1697),
.D(n_1623),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1713),
.Y(n_1724)
);

NAND4xp75_ASAP7_75t_L g1725 ( 
.A(n_1718),
.B(n_1644),
.C(n_1623),
.D(n_1634),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1716),
.B(n_1633),
.C(n_1634),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1715),
.B(n_1626),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1725),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1726),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1722),
.A2(n_1714),
.B1(n_1720),
.B2(n_1716),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1727),
.B(n_1721),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1724),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1723),
.B(n_1626),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1725),
.Y(n_1734)
);

XNOR2xp5_ASAP7_75t_L g1735 ( 
.A(n_1730),
.B(n_1339),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1733),
.B(n_1719),
.Y(n_1736)
);

NAND4xp75_ASAP7_75t_L g1737 ( 
.A(n_1728),
.B(n_1717),
.C(n_1634),
.D(n_1644),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1316),
.C(n_1635),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1729),
.B(n_1607),
.Y(n_1739)
);

NAND5xp2_ASAP7_75t_L g1740 ( 
.A(n_1734),
.B(n_1610),
.C(n_1585),
.D(n_1598),
.E(n_1611),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1736),
.A2(n_1731),
.B1(n_1644),
.B2(n_1640),
.C(n_1635),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1739),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1735),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1731),
.B(n_1738),
.Y(n_1744)
);

OR5x1_ASAP7_75t_L g1745 ( 
.A(n_1744),
.B(n_1737),
.C(n_1741),
.D(n_1740),
.E(n_1743),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1745),
.B(n_1640),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1640),
.B(n_1588),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_SL g1748 ( 
.A1(n_1747),
.A2(n_1588),
.B(n_1585),
.Y(n_1748)
);

AO22x2_ASAP7_75t_L g1749 ( 
.A1(n_1746),
.A2(n_1611),
.B1(n_1598),
.B2(n_1599),
.Y(n_1749)
);

AOI221x1_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1599),
.B1(n_1532),
.B2(n_1533),
.C(n_1557),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1748),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1751),
.B(n_1449),
.C(n_1393),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1750),
.B1(n_1257),
.B2(n_1564),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_R g1754 ( 
.A1(n_1753),
.A2(n_1564),
.B1(n_1559),
.B2(n_1557),
.C(n_1555),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1238),
.B(n_1392),
.C(n_1393),
.Y(n_1755)
);


endmodule