module real_aes_17299_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1872;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_1380;
wire n_488;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_1499;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_1856;
wire n_658;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_1840;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_1772;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1761;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1842;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_0), .A2(n_62), .B1(n_708), .B2(n_1155), .Y(n_1154) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_0), .Y(n_1173) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1), .Y(n_1211) );
OAI22xp33_ASAP7_75t_L g1426 ( .A1(n_2), .A2(n_337), .B1(n_496), .B2(n_766), .Y(n_1426) );
OAI22xp33_ASAP7_75t_SL g1436 ( .A1(n_2), .A2(n_337), .B1(n_458), .B2(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g983 ( .A(n_3), .Y(n_983) );
INVx1_ASAP7_75t_L g391 ( .A(n_4), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_4), .B(n_401), .Y(n_539) );
AND2x2_ASAP7_75t_L g1789 ( .A(n_4), .B(n_268), .Y(n_1789) );
AND2x2_ASAP7_75t_L g1805 ( .A(n_4), .B(n_501), .Y(n_1805) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_5), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_6), .A2(n_272), .B1(n_546), .B2(n_942), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_6), .A2(n_219), .B1(n_448), .B2(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g1038 ( .A(n_7), .Y(n_1038) );
OAI22xp33_ASAP7_75t_L g1489 ( .A1(n_8), .A2(n_61), .B1(n_393), .B2(n_766), .Y(n_1489) );
OAI22xp33_ASAP7_75t_L g1518 ( .A1(n_8), .A2(n_61), .B1(n_721), .B2(n_745), .Y(n_1518) );
OAI22xp5_ASAP7_75t_SL g1054 ( .A1(n_9), .A2(n_242), .B1(n_715), .B2(n_761), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_9), .A2(n_242), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
INVx1_ASAP7_75t_L g1393 ( .A(n_10), .Y(n_1393) );
OAI22xp33_ASAP7_75t_SL g851 ( .A1(n_11), .A2(n_362), .B1(n_496), .B2(n_852), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_11), .A2(n_198), .B1(n_458), .B2(n_479), .Y(n_867) );
INVx1_ASAP7_75t_L g1025 ( .A(n_12), .Y(n_1025) );
INVx1_ASAP7_75t_L g933 ( .A(n_13), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_13), .A2(n_272), .B1(n_418), .B2(n_962), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_14), .A2(n_165), .B1(n_393), .B2(n_766), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_14), .A2(n_165), .B1(n_479), .B2(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1218 ( .A(n_15), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_16), .A2(n_162), .B1(n_393), .B2(n_766), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_16), .A2(n_162), .B1(n_745), .B2(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1134 ( .A(n_17), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_18), .A2(n_46), .B1(n_721), .B2(n_745), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g765 ( .A1(n_18), .A2(n_46), .B1(n_393), .B2(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g1286 ( .A(n_19), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g1295 ( .A1(n_19), .A2(n_316), .B1(n_626), .B2(n_1296), .C(n_1297), .Y(n_1295) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_20), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g1433 ( .A1(n_21), .A2(n_318), .B1(n_506), .B2(n_1434), .Y(n_1433) );
OAI22xp33_ASAP7_75t_L g1441 ( .A1(n_21), .A2(n_318), .B1(n_460), .B2(n_481), .Y(n_1441) );
INVx2_ASAP7_75t_L g439 ( .A(n_22), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g1569 ( .A1(n_23), .A2(n_26), .B1(n_1533), .B2(n_1541), .Y(n_1569) );
INVx1_ASAP7_75t_L g470 ( .A(n_24), .Y(n_470) );
INVx1_ASAP7_75t_L g464 ( .A(n_25), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g1124 ( .A(n_26), .B(n_1125), .Y(n_1124) );
OAI22xp33_ASAP7_75t_SL g1344 ( .A1(n_27), .A2(n_284), .B1(n_458), .B2(n_479), .Y(n_1344) );
OAI22xp33_ASAP7_75t_L g1351 ( .A1(n_27), .A2(n_284), .B1(n_496), .B2(n_582), .Y(n_1351) );
INVx1_ASAP7_75t_L g659 ( .A(n_28), .Y(n_659) );
INVx1_ASAP7_75t_L g603 ( .A(n_29), .Y(n_603) );
INVx1_ASAP7_75t_L g1882 ( .A(n_30), .Y(n_1882) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_31), .A2(n_301), .B1(n_1305), .B2(n_1307), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_31), .A2(n_169), .B1(n_1314), .B2(n_1315), .Y(n_1313) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_32), .A2(n_98), .B1(n_426), .B2(n_430), .C(n_435), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_32), .A2(n_43), .B1(n_557), .B2(n_560), .Y(n_556) );
INVx1_ASAP7_75t_L g1251 ( .A(n_33), .Y(n_1251) );
AOI22xp33_ASAP7_75t_SL g1370 ( .A1(n_34), .A2(n_177), .B1(n_546), .B2(n_1170), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_34), .A2(n_225), .B1(n_630), .B2(n_1315), .Y(n_1382) );
INVx1_ASAP7_75t_L g651 ( .A(n_35), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_36), .A2(n_701), .B(n_704), .C(n_710), .Y(n_700) );
INVx1_ASAP7_75t_L g733 ( .A(n_36), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g995 ( .A1(n_37), .A2(n_97), .B1(n_460), .B2(n_479), .C(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1011 ( .A(n_37), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_38), .Y(n_386) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_38), .B(n_384), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1614 ( .A1(n_39), .A2(n_215), .B1(n_1541), .B2(n_1565), .Y(n_1614) );
INVx1_ASAP7_75t_L g1052 ( .A(n_40), .Y(n_1052) );
INVx1_ASAP7_75t_L g1089 ( .A(n_41), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_42), .A2(n_205), .B1(n_723), .B2(n_1260), .Y(n_1259) );
OAI22xp33_ASAP7_75t_L g1268 ( .A1(n_42), .A2(n_205), .B1(n_393), .B2(n_913), .Y(n_1268) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_43), .A2(n_80), .B1(n_426), .B2(n_430), .C(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_SL g1153 ( .A(n_44), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_44), .A2(n_62), .B1(n_859), .B2(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1873 ( .A(n_45), .Y(n_1873) );
INVx1_ASAP7_75t_L g1453 ( .A(n_47), .Y(n_1453) );
INVx1_ASAP7_75t_L g1506 ( .A(n_48), .Y(n_1506) );
INVx1_ASAP7_75t_L g771 ( .A(n_49), .Y(n_771) );
INVx1_ASAP7_75t_L g1265 ( .A(n_50), .Y(n_1265) );
OAI211xp5_ASAP7_75t_L g1269 ( .A1(n_50), .A2(n_701), .B(n_756), .C(n_1270), .Y(n_1269) );
XNOR2x1_ASAP7_75t_L g1321 ( .A(n_51), .B(n_1322), .Y(n_1321) );
AOI22xp5_ASAP7_75t_L g1563 ( .A1(n_51), .A2(n_232), .B1(n_1533), .B2(n_1538), .Y(n_1563) );
AOI22xp5_ASAP7_75t_L g1549 ( .A1(n_52), .A2(n_354), .B1(n_1541), .B2(n_1550), .Y(n_1549) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_53), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_54), .Y(n_929) );
INVx1_ASAP7_75t_L g1414 ( .A(n_55), .Y(n_1414) );
AOI22xp33_ASAP7_75t_SL g1363 ( .A1(n_56), .A2(n_225), .B1(n_916), .B2(n_1364), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_56), .A2(n_177), .B1(n_1374), .B2(n_1375), .Y(n_1373) );
INVx1_ASAP7_75t_L g449 ( .A(n_57), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_57), .A2(n_275), .B1(n_541), .B2(n_546), .Y(n_540) );
INVx1_ASAP7_75t_L g986 ( .A(n_58), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g1564 ( .A1(n_59), .A2(n_327), .B1(n_1541), .B2(n_1565), .Y(n_1564) );
XNOR2xp5_ASAP7_75t_L g1189 ( .A(n_60), .B(n_1190), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_60), .A2(n_136), .B1(n_1533), .B2(n_1538), .Y(n_1573) );
INVx1_ASAP7_75t_L g618 ( .A(n_63), .Y(n_618) );
INVx1_ASAP7_75t_L g1035 ( .A(n_64), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_65), .B(n_438), .Y(n_998) );
INVxp67_ASAP7_75t_SL g1007 ( .A(n_65), .Y(n_1007) );
OAI211xp5_ASAP7_75t_SL g746 ( .A1(n_66), .A2(n_726), .B(n_727), .C(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g759 ( .A(n_66), .Y(n_759) );
OAI211xp5_ASAP7_75t_L g1853 ( .A1(n_67), .A2(n_467), .B(n_1854), .C(n_1856), .Y(n_1853) );
INVx1_ASAP7_75t_L g1864 ( .A(n_67), .Y(n_1864) );
OAI211xp5_ASAP7_75t_L g844 ( .A1(n_68), .A2(n_574), .B(n_845), .C(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g866 ( .A(n_68), .Y(n_866) );
INVx1_ASAP7_75t_L g1250 ( .A(n_69), .Y(n_1250) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_70), .A2(n_192), .B1(n_735), .B2(n_736), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_70), .A2(n_192), .B1(n_761), .B2(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g1033 ( .A(n_71), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_72), .Y(n_813) );
INVx1_ASAP7_75t_L g1157 ( .A(n_73), .Y(n_1157) );
OAI222xp33_ASAP7_75t_L g917 ( .A1(n_74), .A2(n_202), .B1(n_497), .B2(n_850), .C1(n_918), .C2(n_919), .Y(n_917) );
OAI222xp33_ASAP7_75t_L g948 ( .A1(n_74), .A2(n_202), .B1(n_243), .B2(n_949), .C1(n_950), .C2(n_951), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g1291 ( .A1(n_75), .A2(n_133), .B1(n_506), .B2(n_507), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g1298 ( .A1(n_75), .A2(n_133), .B1(n_460), .B2(n_481), .Y(n_1298) );
OAI211xp5_ASAP7_75t_L g1465 ( .A1(n_76), .A2(n_753), .B(n_756), .C(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1474 ( .A(n_76), .Y(n_1474) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_77), .A2(n_320), .B1(n_393), .B2(n_766), .Y(n_1111) );
OAI22xp33_ASAP7_75t_L g1113 ( .A1(n_77), .A2(n_320), .B1(n_745), .B2(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g709 ( .A(n_78), .Y(n_709) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_78), .A2(n_726), .B(n_727), .C(n_728), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g1001 ( .A1(n_79), .A2(n_207), .B1(n_458), .B2(n_1002), .Y(n_1001) );
INVxp67_ASAP7_75t_SL g1009 ( .A(n_79), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_80), .A2(n_98), .B1(n_549), .B2(n_551), .Y(n_548) );
INVx1_ASAP7_75t_L g1388 ( .A(n_81), .Y(n_1388) );
INVx1_ASAP7_75t_L g1413 ( .A(n_82), .Y(n_1413) );
INVx1_ASAP7_75t_L g1881 ( .A(n_83), .Y(n_1881) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_84), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g1266 ( .A1(n_85), .A2(n_190), .B1(n_735), .B2(n_1121), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_85), .A2(n_190), .B1(n_713), .B2(n_1110), .Y(n_1272) );
INVx1_ASAP7_75t_L g1158 ( .A(n_86), .Y(n_1158) );
INVx1_ASAP7_75t_L g1879 ( .A(n_87), .Y(n_1879) );
INVx1_ASAP7_75t_L g784 ( .A(n_88), .Y(n_784) );
INVx1_ASAP7_75t_L g1336 ( .A(n_89), .Y(n_1336) );
INVx1_ASAP7_75t_L g1148 ( .A(n_90), .Y(n_1148) );
XNOR2xp5_ASAP7_75t_L g1276 ( .A(n_91), .B(n_1277), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1779 ( .A1(n_92), .A2(n_340), .B1(n_413), .B2(n_418), .Y(n_1779) );
AOI221xp5_ASAP7_75t_L g1811 ( .A1(n_92), .A2(n_356), .B1(n_549), .B2(n_1812), .C(n_1814), .Y(n_1811) );
INVx1_ASAP7_75t_L g1196 ( .A(n_93), .Y(n_1196) );
OAI211xp5_ASAP7_75t_L g1203 ( .A1(n_93), .A2(n_726), .B(n_727), .C(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g985 ( .A(n_94), .Y(n_985) );
OAI22xp33_ASAP7_75t_L g1349 ( .A1(n_95), .A2(n_126), .B1(n_460), .B2(n_481), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1355 ( .A1(n_95), .A2(n_126), .B1(n_506), .B2(n_507), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_96), .A2(n_365), .B1(n_1533), .B2(n_1538), .Y(n_1554) );
OAI22xp33_ASAP7_75t_L g1013 ( .A1(n_97), .A2(n_207), .B1(n_496), .B2(n_582), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_99), .A2(n_217), .B1(n_458), .B2(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g494 ( .A(n_99), .Y(n_494) );
INVx1_ASAP7_75t_L g664 ( .A(n_100), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_101), .A2(n_292), .B1(n_496), .B2(n_507), .Y(n_895) );
OAI22xp5_ASAP7_75t_SL g903 ( .A1(n_101), .A2(n_143), .B1(n_458), .B2(n_481), .Y(n_903) );
INVx1_ASAP7_75t_L g783 ( .A(n_102), .Y(n_783) );
INVx1_ASAP7_75t_L g1000 ( .A(n_103), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_104), .Y(n_898) );
INVx1_ASAP7_75t_L g1858 ( .A(n_105), .Y(n_1858) );
OAI211xp5_ASAP7_75t_L g1862 ( .A1(n_105), .A2(n_932), .B(n_1193), .C(n_1863), .Y(n_1862) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_106), .Y(n_874) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_107), .A2(n_174), .B1(n_393), .B2(n_582), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_107), .A2(n_174), .B1(n_721), .B2(n_723), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_108), .Y(n_812) );
INVx1_ASAP7_75t_L g474 ( .A(n_109), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g1371 ( .A1(n_110), .A2(n_373), .B1(n_916), .B2(n_1364), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_110), .A2(n_112), .B1(n_1377), .B2(n_1380), .Y(n_1384) );
OAI22xp33_ASAP7_75t_SL g1495 ( .A1(n_111), .A2(n_291), .B1(n_713), .B2(n_1198), .Y(n_1495) );
OAI22xp33_ASAP7_75t_L g1522 ( .A1(n_111), .A2(n_291), .B1(n_736), .B2(n_1476), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_112), .A2(n_341), .B1(n_546), .B2(n_1368), .Y(n_1367) );
AOI22xp5_ASAP7_75t_SL g1555 ( .A1(n_113), .A2(n_240), .B1(n_1541), .B2(n_1550), .Y(n_1555) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_114), .A2(n_261), .B1(n_1305), .B2(n_1309), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_114), .A2(n_183), .B1(n_465), .B2(n_1317), .Y(n_1316) );
XOR2xp5_ASAP7_75t_L g807 ( .A(n_115), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g1407 ( .A(n_116), .Y(n_1407) );
INVx1_ASAP7_75t_L g1136 ( .A(n_117), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_117), .A2(n_312), .B1(n_1164), .B2(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1878 ( .A(n_118), .Y(n_1878) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_119), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g1754 ( .A1(n_120), .A2(n_249), .B1(n_1755), .B2(n_1761), .C(n_1765), .Y(n_1754) );
OAI211xp5_ASAP7_75t_L g1800 ( .A1(n_120), .A2(n_1801), .B(n_1806), .C(n_1815), .Y(n_1800) );
INVx1_ASAP7_75t_L g1095 ( .A(n_121), .Y(n_1095) );
INVx1_ASAP7_75t_L g384 ( .A(n_122), .Y(n_384) );
INVx1_ASAP7_75t_L g1028 ( .A(n_123), .Y(n_1028) );
INVx1_ASAP7_75t_L g1511 ( .A(n_124), .Y(n_1511) );
INVx1_ASAP7_75t_L g1144 ( .A(n_125), .Y(n_1144) );
XOR2xp5_ASAP7_75t_L g909 ( .A(n_127), .B(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g1214 ( .A(n_128), .Y(n_1214) );
INVx1_ASAP7_75t_L g1329 ( .A(n_129), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g1791 ( .A1(n_130), .A2(n_286), .B1(n_1792), .B2(n_1796), .Y(n_1791) );
INVx1_ASAP7_75t_L g1326 ( .A(n_131), .Y(n_1326) );
AOI22xp5_ASAP7_75t_L g1557 ( .A1(n_132), .A2(n_345), .B1(n_1538), .B2(n_1550), .Y(n_1557) );
INVx1_ASAP7_75t_L g1081 ( .A(n_134), .Y(n_1081) );
INVx1_ASAP7_75t_L g1493 ( .A(n_135), .Y(n_1493) );
INVx1_ASAP7_75t_L g1132 ( .A(n_137), .Y(n_1132) );
INVx1_ASAP7_75t_L g1417 ( .A(n_138), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g1460 ( .A1(n_139), .A2(n_211), .B1(n_587), .B2(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1480 ( .A(n_139), .Y(n_1480) );
INVx1_ASAP7_75t_L g1857 ( .A(n_140), .Y(n_1857) );
INVx1_ASAP7_75t_L g611 ( .A(n_141), .Y(n_611) );
OAI22xp33_ASAP7_75t_SL g900 ( .A1(n_142), .A2(n_143), .B1(n_506), .B2(n_582), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_142), .A2(n_147), .B1(n_864), .B2(n_865), .Y(n_907) );
INVx1_ASAP7_75t_L g788 ( .A(n_144), .Y(n_788) );
INVx1_ASAP7_75t_L g616 ( .A(n_145), .Y(n_616) );
INVx1_ASAP7_75t_L g1429 ( .A(n_146), .Y(n_1429) );
INVx1_ASAP7_75t_L g899 ( .A(n_147), .Y(n_899) );
INVx1_ASAP7_75t_L g1248 ( .A(n_148), .Y(n_1248) );
INVx1_ASAP7_75t_L g1876 ( .A(n_149), .Y(n_1876) );
XOR2xp5_ASAP7_75t_L g1846 ( .A(n_150), .B(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g613 ( .A(n_151), .Y(n_613) );
AOI31xp33_ASAP7_75t_L g410 ( .A1(n_152), .A2(n_411), .A3(n_456), .B(n_492), .Y(n_410) );
NAND2xp33_ASAP7_75t_SL g534 ( .A(n_152), .B(n_535), .Y(n_534) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_152), .Y(n_563) );
INVx1_ASAP7_75t_L g1280 ( .A(n_153), .Y(n_1280) );
INVx1_ASAP7_75t_L g1348 ( .A(n_154), .Y(n_1348) );
OAI211xp5_ASAP7_75t_L g1352 ( .A1(n_154), .A2(n_574), .B(n_607), .C(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1774 ( .A(n_155), .Y(n_1774) );
CKINVDCx5p33_ASAP7_75t_R g1347 ( .A(n_156), .Y(n_1347) );
INVx1_ASAP7_75t_L g653 ( .A(n_157), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_158), .Y(n_879) );
OAI22xp33_ASAP7_75t_L g1859 ( .A1(n_159), .A2(n_173), .B1(n_1066), .B2(n_1860), .Y(n_1859) );
OAI22xp33_ASAP7_75t_L g1867 ( .A1(n_159), .A2(n_173), .B1(n_496), .B2(n_766), .Y(n_1867) );
INVx1_ASAP7_75t_L g777 ( .A(n_160), .Y(n_777) );
INVx1_ASAP7_75t_L g1409 ( .A(n_161), .Y(n_1409) );
INVx1_ASAP7_75t_L g748 ( .A(n_163), .Y(n_748) );
INVx1_ASAP7_75t_L g666 ( .A(n_164), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_166), .Y(n_816) );
OAI211xp5_ASAP7_75t_L g1105 ( .A1(n_167), .A2(n_755), .B(n_756), .C(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1119 ( .A(n_167), .Y(n_1119) );
CKINVDCx20_ASAP7_75t_R g1222 ( .A(n_168), .Y(n_1222) );
AOI22xp33_ASAP7_75t_SL g1310 ( .A1(n_169), .A2(n_227), .B1(n_1165), .B2(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1107 ( .A(n_170), .Y(n_1107) );
INVxp67_ASAP7_75t_SL g1769 ( .A(n_171), .Y(n_1769) );
AOI221xp5_ASAP7_75t_L g1827 ( .A1(n_171), .A2(n_274), .B1(n_1366), .B2(n_1812), .C(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1392 ( .A(n_172), .Y(n_1392) );
INVx1_ASAP7_75t_L g981 ( .A(n_175), .Y(n_981) );
OAI211xp5_ASAP7_75t_SL g1050 ( .A1(n_176), .A2(n_701), .B(n_756), .C(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1064 ( .A(n_176), .Y(n_1064) );
INVx1_ASAP7_75t_L g609 ( .A(n_178), .Y(n_609) );
INVx1_ASAP7_75t_L g1195 ( .A(n_179), .Y(n_1195) );
INVx1_ASAP7_75t_L g1494 ( .A(n_180), .Y(n_1494) );
OAI211xp5_ASAP7_75t_L g1519 ( .A1(n_180), .A2(n_726), .B(n_727), .C(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1281 ( .A(n_181), .Y(n_1281) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_182), .A2(n_310), .B1(n_761), .B2(n_1110), .Y(n_1109) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_182), .A2(n_310), .B1(n_735), .B2(n_1121), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_183), .A2(n_279), .B1(n_560), .B2(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1875 ( .A(n_184), .Y(n_1875) );
INVx1_ASAP7_75t_L g1790 ( .A(n_185), .Y(n_1790) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_186), .Y(n_823) );
INVx1_ASAP7_75t_L g1611 ( .A(n_187), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_188), .Y(n_1285) );
AOI22xp5_ASAP7_75t_SL g1572 ( .A1(n_189), .A2(n_200), .B1(n_1541), .B2(n_1550), .Y(n_1572) );
INVx1_ASAP7_75t_L g1094 ( .A(n_191), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_193), .A2(n_270), .B1(n_713), .B2(n_1198), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_193), .A2(n_270), .B1(n_1058), .B2(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g749 ( .A(n_194), .Y(n_749) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_194), .A2(n_753), .B(n_756), .C(n_757), .Y(n_752) );
INVx1_ASAP7_75t_L g1221 ( .A(n_195), .Y(n_1221) );
OAI211xp5_ASAP7_75t_L g1345 ( .A1(n_196), .A2(n_467), .B(n_1143), .C(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1354 ( .A(n_196), .Y(n_1354) );
INVx1_ASAP7_75t_L g1504 ( .A(n_197), .Y(n_1504) );
OAI22xp33_ASAP7_75t_SL g854 ( .A1(n_198), .A2(n_322), .B1(n_714), .B2(n_766), .Y(n_854) );
INVx1_ASAP7_75t_L g1500 ( .A(n_199), .Y(n_1500) );
INVx1_ASAP7_75t_L g1076 ( .A(n_201), .Y(n_1076) );
INVx1_ASAP7_75t_L g595 ( .A(n_203), .Y(n_595) );
INVx2_ASAP7_75t_L g1536 ( .A(n_204), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_204), .B(n_1537), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_204), .B(n_317), .Y(n_1544) );
AO22x2_ASAP7_75t_L g1401 ( .A1(n_206), .A2(n_1402), .B1(n_1442), .B2(n_1443), .Y(n_1401) );
INVx1_ASAP7_75t_L g1442 ( .A(n_206), .Y(n_1442) );
INVx1_ASAP7_75t_L g1510 ( .A(n_208), .Y(n_1510) );
AOI22xp5_ASAP7_75t_SL g1568 ( .A1(n_209), .A2(n_277), .B1(n_1538), .B2(n_1543), .Y(n_1568) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_210), .Y(n_881) );
INVx1_ASAP7_75t_L g1484 ( .A(n_211), .Y(n_1484) );
INVx1_ASAP7_75t_L g1217 ( .A(n_212), .Y(n_1217) );
INVx1_ASAP7_75t_L g773 ( .A(n_213), .Y(n_773) );
INVx1_ASAP7_75t_L g1243 ( .A(n_214), .Y(n_1243) );
XNOR2xp5_ASAP7_75t_L g1018 ( .A(n_216), .B(n_1019), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_217), .A2(n_298), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g1540 ( .A1(n_218), .A2(n_338), .B1(n_1541), .B2(n_1543), .Y(n_1540) );
INVx1_ASAP7_75t_L g934 ( .A(n_219), .Y(n_934) );
XOR2xp5_ASAP7_75t_L g969 ( .A(n_220), .B(n_970), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g1548 ( .A1(n_220), .A2(n_282), .B1(n_1533), .B2(n_1538), .Y(n_1548) );
XNOR2x2_ASAP7_75t_L g645 ( .A(n_221), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g975 ( .A(n_222), .Y(n_975) );
INVx1_ASAP7_75t_L g579 ( .A(n_223), .Y(n_579) );
INVx1_ASAP7_75t_L g1467 ( .A(n_224), .Y(n_1467) );
AOI22xp5_ASAP7_75t_L g1558 ( .A1(n_226), .A2(n_300), .B1(n_1533), .B2(n_1541), .Y(n_1558) );
AOI22xp33_ASAP7_75t_SL g1318 ( .A1(n_227), .A2(n_301), .B1(n_1315), .B2(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1032 ( .A(n_228), .Y(n_1032) );
INVx1_ASAP7_75t_L g1240 ( .A(n_229), .Y(n_1240) );
OAI211xp5_ASAP7_75t_L g912 ( .A1(n_230), .A2(n_913), .B(n_914), .C(n_923), .Y(n_912) );
INVx1_ASAP7_75t_L g955 ( .A(n_230), .Y(n_955) );
INVx1_ASAP7_75t_L g1082 ( .A(n_231), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1852 ( .A1(n_233), .A2(n_250), .B1(n_735), .B2(n_1059), .Y(n_1852) );
OAI22xp5_ASAP7_75t_L g1866 ( .A1(n_233), .A2(n_250), .B1(n_713), .B2(n_715), .Y(n_1866) );
INVx1_ASAP7_75t_L g978 ( .A(n_234), .Y(n_978) );
INVx2_ASAP7_75t_L g437 ( .A(n_235), .Y(n_437) );
INVx1_ASAP7_75t_L g454 ( .A(n_235), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_235), .B(n_439), .Y(n_1753) );
XOR2xp5_ASAP7_75t_L g1234 ( .A(n_236), .B(n_1235), .Y(n_1234) );
XNOR2xp5_ASAP7_75t_L g1486 ( .A(n_237), .B(n_1487), .Y(n_1486) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_238), .A2(n_296), .B1(n_506), .B2(n_507), .Y(n_568) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_238), .A2(n_260), .B1(n_458), .B2(n_460), .Y(n_584) );
INVx1_ASAP7_75t_L g1333 ( .A(n_239), .Y(n_1333) );
INVx1_ASAP7_75t_L g922 ( .A(n_241), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_241), .A2(n_267), .B1(n_460), .B2(n_481), .Y(n_952) );
INVx1_ASAP7_75t_L g915 ( .A(n_243), .Y(n_915) );
BUFx3_ASAP7_75t_L g417 ( .A(n_244), .Y(n_417) );
INVx1_ASAP7_75t_L g1327 ( .A(n_245), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1464 ( .A1(n_246), .A2(n_366), .B1(n_393), .B2(n_766), .Y(n_1464) );
OAI22xp33_ASAP7_75t_L g1471 ( .A1(n_246), .A2(n_366), .B1(n_745), .B2(n_1397), .Y(n_1471) );
XOR2xp5_ASAP7_75t_L g1071 ( .A(n_247), .B(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1468 ( .A(n_248), .Y(n_1468) );
OAI211xp5_ASAP7_75t_L g1472 ( .A1(n_248), .A2(n_727), .B(n_1117), .C(n_1473), .Y(n_1472) );
OAI221xp5_ASAP7_75t_SL g1817 ( .A1(n_249), .A2(n_351), .B1(n_1818), .B2(n_1821), .C(n_1825), .Y(n_1817) );
AOI22xp5_ASAP7_75t_L g1532 ( .A1(n_251), .A2(n_295), .B1(n_1533), .B2(n_1538), .Y(n_1532) );
INVx1_ASAP7_75t_L g1139 ( .A(n_252), .Y(n_1139) );
INVx1_ASAP7_75t_L g1391 ( .A(n_253), .Y(n_1391) );
INVx1_ASAP7_75t_L g927 ( .A(n_254), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_254), .B(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g1430 ( .A(n_255), .Y(n_1430) );
INVx1_ASAP7_75t_L g1079 ( .A(n_256), .Y(n_1079) );
INVx1_ASAP7_75t_L g1246 ( .A(n_257), .Y(n_1246) );
OAI22xp33_ASAP7_75t_L g1199 ( .A1(n_258), .A2(n_336), .B1(n_393), .B2(n_766), .Y(n_1199) );
OAI22xp33_ASAP7_75t_L g1207 ( .A1(n_258), .A2(n_336), .B1(n_721), .B2(n_745), .Y(n_1207) );
INVx1_ASAP7_75t_L g576 ( .A(n_259), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_260), .A2(n_303), .B1(n_496), .B2(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g1320 ( .A1(n_261), .A2(n_279), .B1(n_435), .B2(n_445), .C(n_1317), .Y(n_1320) );
INVx1_ASAP7_75t_L g1142 ( .A(n_262), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_262), .A2(n_319), .B1(n_1163), .B2(n_1164), .Y(n_1162) );
INVx1_ASAP7_75t_L g1406 ( .A(n_263), .Y(n_1406) );
INVx1_ASAP7_75t_L g1332 ( .A(n_264), .Y(n_1332) );
XOR2xp5_ASAP7_75t_L g869 ( .A(n_265), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g1215 ( .A(n_266), .Y(n_1215) );
INVx1_ASAP7_75t_L g924 ( .A(n_267), .Y(n_924) );
BUFx3_ASAP7_75t_L g401 ( .A(n_268), .Y(n_401) );
INVx1_ASAP7_75t_L g501 ( .A(n_268), .Y(n_501) );
INVx1_ASAP7_75t_L g706 ( .A(n_269), .Y(n_706) );
XOR2x2_ASAP7_75t_L g741 ( .A(n_271), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g974 ( .A(n_273), .Y(n_974) );
INVx1_ASAP7_75t_L g1777 ( .A(n_274), .Y(n_1777) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_275), .A2(n_307), .B1(n_413), .B2(n_418), .Y(n_412) );
XNOR2x1_ASAP7_75t_L g1447 ( .A(n_276), .B(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g674 ( .A(n_278), .Y(n_674) );
INVx1_ASAP7_75t_L g1454 ( .A(n_280), .Y(n_1454) );
OAI322xp33_ASAP7_75t_SL g1767 ( .A1(n_281), .A2(n_1090), .A3(n_1127), .B1(n_1768), .B2(n_1773), .C1(n_1776), .C2(n_1780), .Y(n_1767) );
OAI22xp33_ASAP7_75t_SL g1829 ( .A1(n_281), .A2(n_286), .B1(n_1830), .B2(n_1833), .Y(n_1829) );
OAI211xp5_ASAP7_75t_L g1490 ( .A1(n_283), .A2(n_710), .B(n_1491), .C(n_1492), .Y(n_1490) );
INVx1_ASAP7_75t_L g1521 ( .A(n_283), .Y(n_1521) );
INVx1_ASAP7_75t_L g1239 ( .A(n_285), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1455 ( .A1(n_287), .A2(n_369), .B1(n_997), .B2(n_1456), .Y(n_1455) );
INVxp33_ASAP7_75t_SL g1479 ( .A(n_287), .Y(n_1479) );
OAI211xp5_ASAP7_75t_L g569 ( .A1(n_288), .A2(n_570), .B(n_574), .C(n_575), .Y(n_569) );
INVx1_ASAP7_75t_L g589 ( .A(n_288), .Y(n_589) );
INVx1_ASAP7_75t_L g1778 ( .A(n_289), .Y(n_1778) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_290), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_292), .B(n_460), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_293), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_294), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g1743 ( .A1(n_295), .A2(n_1744), .B1(n_1745), .B2(n_1836), .Y(n_1743) );
INVx1_ASAP7_75t_L g1836 ( .A(n_295), .Y(n_1836) );
AOI22xp33_ASAP7_75t_L g1841 ( .A1(n_295), .A2(n_1842), .B1(n_1845), .B2(n_1891), .Y(n_1841) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_296), .A2(n_303), .B1(n_479), .B2(n_481), .Y(n_590) );
XOR2x2_ASAP7_75t_L g1359 ( .A(n_297), .B(n_1360), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_298), .A2(n_339), .B1(n_479), .B2(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g1389 ( .A(n_299), .Y(n_1389) );
INVx1_ASAP7_75t_L g416 ( .A(n_302), .Y(n_416) );
INVx1_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
INVx1_ASAP7_75t_L g673 ( .A(n_304), .Y(n_673) );
INVx1_ASAP7_75t_L g657 ( .A(n_305), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g1469 ( .A1(n_306), .A2(n_357), .B1(n_761), .B2(n_1110), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_306), .A2(n_357), .B1(n_1121), .B2(n_1476), .Y(n_1475) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_307), .A2(n_343), .B1(n_549), .B2(n_551), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_308), .A2(n_358), .B1(n_713), .B2(n_715), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_308), .A2(n_358), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g1458 ( .A(n_309), .Y(n_1458) );
OAI211xp5_ASAP7_75t_L g1261 ( .A1(n_311), .A2(n_727), .B(n_1262), .C(n_1263), .Y(n_1261) );
INVx1_ASAP7_75t_L g1271 ( .A(n_311), .Y(n_1271) );
INVx1_ASAP7_75t_L g1140 ( .A(n_312), .Y(n_1140) );
INVx1_ASAP7_75t_L g847 ( .A(n_313), .Y(n_847) );
OAI211xp5_ASAP7_75t_SL g858 ( .A1(n_313), .A2(n_727), .B(n_859), .C(n_861), .Y(n_858) );
INVx1_ASAP7_75t_L g779 ( .A(n_314), .Y(n_779) );
INVx1_ASAP7_75t_L g977 ( .A(n_315), .Y(n_977) );
INVx1_ASAP7_75t_L g1290 ( .A(n_316), .Y(n_1290) );
INVx1_ASAP7_75t_L g1537 ( .A(n_317), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_317), .B(n_1536), .Y(n_1542) );
INVx1_ASAP7_75t_L g1129 ( .A(n_319), .Y(n_1129) );
INVx1_ASAP7_75t_L g1335 ( .A(n_321), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_322), .A2(n_362), .B1(n_460), .B2(n_481), .Y(n_857) );
INVx1_ASAP7_75t_L g1147 ( .A(n_323), .Y(n_1147) );
INVx1_ASAP7_75t_L g1613 ( .A(n_324), .Y(n_1613) );
INVx1_ASAP7_75t_L g1416 ( .A(n_325), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_326), .Y(n_936) );
OAI211xp5_ASAP7_75t_SL g896 ( .A1(n_328), .A2(n_574), .B(n_845), .C(n_897), .Y(n_896) );
OAI211xp5_ASAP7_75t_SL g904 ( .A1(n_328), .A2(n_727), .B(n_905), .C(n_906), .Y(n_904) );
INVx1_ASAP7_75t_L g1330 ( .A(n_329), .Y(n_1330) );
INVx1_ASAP7_75t_L g601 ( .A(n_330), .Y(n_601) );
INVx1_ASAP7_75t_L g1053 ( .A(n_331), .Y(n_1053) );
OAI211xp5_ASAP7_75t_SL g1060 ( .A1(n_331), .A2(n_727), .B(n_1061), .C(n_1063), .Y(n_1060) );
INVx1_ASAP7_75t_L g999 ( .A(n_332), .Y(n_999) );
INVx1_ASAP7_75t_L g1459 ( .A(n_333), .Y(n_1459) );
INVx1_ASAP7_75t_L g1508 ( .A(n_334), .Y(n_1508) );
XOR2x2_ASAP7_75t_L g565 ( .A(n_335), .B(n_566), .Y(n_565) );
INVxp67_ASAP7_75t_SL g498 ( .A(n_339), .Y(n_498) );
INVxp67_ASAP7_75t_SL g1826 ( .A(n_340), .Y(n_1826) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_341), .A2(n_373), .B1(n_1377), .B2(n_1380), .Y(n_1376) );
INVx1_ASAP7_75t_L g1108 ( .A(n_342), .Y(n_1108) );
OAI211xp5_ASAP7_75t_L g1116 ( .A1(n_342), .A2(n_467), .B(n_1117), .C(n_1118), .Y(n_1116) );
INVx1_ASAP7_75t_L g446 ( .A(n_343), .Y(n_446) );
INVx1_ASAP7_75t_L g1499 ( .A(n_344), .Y(n_1499) );
OAI211xp5_ASAP7_75t_SL g1192 ( .A1(n_346), .A2(n_701), .B(n_1193), .C(n_1194), .Y(n_1192) );
INVx1_ASAP7_75t_L g1206 ( .A(n_346), .Y(n_1206) );
INVx1_ASAP7_75t_L g1212 ( .A(n_347), .Y(n_1212) );
INVx1_ASAP7_75t_L g1871 ( .A(n_348), .Y(n_1871) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_349), .Y(n_829) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_350), .Y(n_397) );
INVxp67_ASAP7_75t_SL g1747 ( .A(n_351), .Y(n_1747) );
INVx1_ASAP7_75t_L g1410 ( .A(n_352), .Y(n_1410) );
INVx1_ASAP7_75t_L g1088 ( .A(n_353), .Y(n_1088) );
INVx1_ASAP7_75t_L g1244 ( .A(n_355), .Y(n_1244) );
INVx1_ASAP7_75t_L g1775 ( .A(n_356), .Y(n_1775) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_359), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_360), .Y(n_878) );
INVx1_ASAP7_75t_L g1432 ( .A(n_361), .Y(n_1432) );
INVx2_ASAP7_75t_L g441 ( .A(n_363), .Y(n_441) );
INVx1_ASAP7_75t_L g491 ( .A(n_363), .Y(n_491) );
INVx1_ASAP7_75t_L g693 ( .A(n_363), .Y(n_693) );
INVx1_ASAP7_75t_L g1264 ( .A(n_364), .Y(n_1264) );
INVx1_ASAP7_75t_L g1503 ( .A(n_367), .Y(n_1503) );
INVx1_ASAP7_75t_L g1024 ( .A(n_368), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1483 ( .A(n_369), .Y(n_1483) );
INVx1_ASAP7_75t_L g1027 ( .A(n_370), .Y(n_1027) );
AOI21xp33_ASAP7_75t_L g938 ( .A1(n_371), .A2(n_549), .B(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g958 ( .A(n_371), .Y(n_958) );
INVx1_ASAP7_75t_L g787 ( .A(n_372), .Y(n_787) );
INVx1_ASAP7_75t_L g1772 ( .A(n_374), .Y(n_1772) );
CKINVDCx5p33_ASAP7_75t_R g920 ( .A(n_375), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_402), .B(n_1524), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_387), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1840 ( .A(n_381), .B(n_390), .Y(n_1840) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g1844 ( .A(n_383), .B(n_386), .Y(n_1844) );
INVx1_ASAP7_75t_L g1895 ( .A(n_383), .Y(n_1895) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g1897 ( .A(n_386), .B(n_1895), .Y(n_1897) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g528 ( .A(n_390), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_SL g911 ( .A1(n_390), .A2(n_912), .B(n_925), .Y(n_911) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g555 ( .A(n_391), .B(n_401), .Y(n_555) );
AND2x4_ASAP7_75t_L g940 ( .A(n_391), .B(n_400), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_392), .A2(n_499), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
AND2x4_ASAP7_75t_SL g1839 ( .A(n_392), .B(n_1840), .Y(n_1839) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .Y(n_393) );
OR2x2_ASAP7_75t_L g506 ( .A(n_394), .B(n_500), .Y(n_506) );
OR2x6_ASAP7_75t_L g714 ( .A(n_394), .B(n_500), .Y(n_714) );
INVx1_ASAP7_75t_L g841 ( .A(n_394), .Y(n_841) );
BUFx4f_ASAP7_75t_L g928 ( .A(n_394), .Y(n_928) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g497 ( .A(n_395), .Y(n_497) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_395), .Y(n_597) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g502 ( .A(n_397), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g511 ( .A(n_397), .Y(n_511) );
INVx1_ASAP7_75t_L g518 ( .A(n_397), .Y(n_518) );
AND2x2_ASAP7_75t_L g524 ( .A(n_397), .B(n_398), .Y(n_524) );
INVx2_ASAP7_75t_L g544 ( .A(n_397), .Y(n_544) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_397), .B(n_398), .Y(n_573) );
INVx2_ASAP7_75t_L g503 ( .A(n_398), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_398), .B(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g515 ( .A(n_398), .Y(n_515) );
INVx1_ASAP7_75t_L g545 ( .A(n_398), .Y(n_545) );
AND2x2_ASAP7_75t_L g547 ( .A(n_398), .B(n_511), .Y(n_547) );
OR2x2_ASAP7_75t_L g606 ( .A(n_398), .B(n_544), .Y(n_606) );
OR2x6_ASAP7_75t_L g496 ( .A(n_399), .B(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_399), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g508 ( .A(n_400), .Y(n_508) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g516 ( .A(n_401), .B(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g578 ( .A(n_401), .Y(n_578) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_1014), .Y(n_402) );
XOR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_804), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_643), .B2(n_803), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
XNOR2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_565), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_531), .Y(n_409) );
INVx1_ASAP7_75t_L g533 ( .A(n_411), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_425), .B(n_442), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g1399 ( .A1(n_413), .A2(n_732), .B1(n_1205), .B2(n_1391), .C1(n_1392), .C2(n_1393), .Y(n_1399) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
INVx2_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
AND2x4_ASAP7_75t_L g468 ( .A(n_414), .B(n_455), .Y(n_468) );
BUFx2_ASAP7_75t_L g587 ( .A(n_414), .Y(n_587) );
BUFx2_ASAP7_75t_L g962 ( .A(n_414), .Y(n_962) );
BUFx2_ASAP7_75t_L g997 ( .A(n_414), .Y(n_997) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
INVx1_ASAP7_75t_L g434 ( .A(n_415), .Y(n_434) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g477 ( .A(n_416), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_416), .B(n_417), .Y(n_483) );
INVx2_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_417), .Y(n_433) );
OR2x2_ASAP7_75t_L g459 ( .A(n_417), .B(n_423), .Y(n_459) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx8_ASAP7_75t_L g1317 ( .A(n_419), .Y(n_1317) );
INVx8_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g448 ( .A(n_420), .Y(n_448) );
BUFx3_ASAP7_75t_L g1379 ( .A(n_420), .Y(n_1379) );
NAND2x1p5_ASAP7_75t_L g1797 ( .A(n_420), .B(n_1759), .Y(n_1797) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AND2x4_ASAP7_75t_L g428 ( .A(n_421), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g429 ( .A(n_424), .Y(n_429) );
INVx1_ASAP7_75t_L g1043 ( .A(n_426), .Y(n_1043) );
INVx1_ASAP7_75t_L g1228 ( .A(n_426), .Y(n_1228) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g480 ( .A(n_427), .B(n_461), .Y(n_480) );
INVx2_ASAP7_75t_L g635 ( .A(n_427), .Y(n_635) );
AND2x4_ASAP7_75t_L g724 ( .A(n_427), .B(n_461), .Y(n_724) );
BUFx6f_ASAP7_75t_L g960 ( .A(n_427), .Y(n_960) );
INVx2_ASAP7_75t_L g1045 ( .A(n_427), .Y(n_1045) );
INVx1_ASAP7_75t_L g1247 ( .A(n_427), .Y(n_1247) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_428), .Y(n_630) );
BUFx8_ASAP7_75t_L g818 ( .A(n_428), .Y(n_818) );
INVx2_ASAP7_75t_L g967 ( .A(n_428), .Y(n_967) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g964 ( .A(n_432), .Y(n_964) );
BUFx12f_ASAP7_75t_L g1315 ( .A(n_432), .Y(n_1315) );
BUFx3_ASAP7_75t_L g1375 ( .A(n_432), .Y(n_1375) );
AND2x4_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
BUFx2_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_433), .B(n_477), .Y(n_627) );
INVx2_ASAP7_75t_L g865 ( .A(n_433), .Y(n_865) );
INVx1_ASAP7_75t_L g863 ( .A(n_434), .Y(n_863) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g1372 ( .A(n_436), .B(n_1373), .C(n_1376), .Y(n_1372) );
AND3x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .C(n_440), .Y(n_436) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_437), .Y(n_486) );
NAND2xp33_ASAP7_75t_SL g622 ( .A(n_437), .B(n_439), .Y(n_622) );
INVx1_ASAP7_75t_L g1760 ( .A(n_437), .Y(n_1760) );
INVx3_ASAP7_75t_L g472 ( .A(n_438), .Y(n_472) );
AND2x2_ASAP7_75t_L g862 ( .A(n_438), .B(n_863), .Y(n_862) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g455 ( .A(n_439), .Y(n_455) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g452 ( .A(n_441), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B1(n_447), .B2(n_449), .C(n_450), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI211xp5_ASAP7_75t_L g1172 ( .A1(n_445), .A2(n_468), .B(n_1173), .C(n_1174), .Y(n_1172) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
AOI32xp33_ASAP7_75t_L g1312 ( .A1(n_450), .A2(n_1313), .A3(n_1316), .B1(n_1318), .B2(n_1320), .Y(n_1312) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI33xp33_ASAP7_75t_L g972 ( .A1(n_451), .A2(n_769), .A3(n_973), .B1(n_976), .B2(n_979), .B3(n_984), .Y(n_972) );
OAI33xp33_ASAP7_75t_L g1418 ( .A1(n_451), .A2(n_769), .A3(n_1419), .B1(n_1420), .B2(n_1421), .B3(n_1424), .Y(n_1418) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AND2x4_ASAP7_75t_L g538 ( .A(n_452), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g637 ( .A(n_452), .B(n_453), .Y(n_637) );
INVx1_ASAP7_75t_L g944 ( .A(n_452), .Y(n_944) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NAND3x1_ASAP7_75t_L g691 ( .A(n_454), .B(n_455), .C(n_692), .Y(n_691) );
OR2x4_ASAP7_75t_L g458 ( .A(n_455), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_455), .Y(n_461) );
OR2x6_ASAP7_75t_L g481 ( .A(n_455), .B(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g1759 ( .A(n_455), .B(n_1760), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_456), .B(n_492), .Y(n_532) );
OAI31xp33_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_462), .A3(n_478), .B(n_484), .Y(n_456) );
INVx2_ASAP7_75t_SL g722 ( .A(n_458), .Y(n_722) );
INVx1_ASAP7_75t_L g954 ( .A(n_458), .Y(n_954) );
INVx1_ASAP7_75t_L g1115 ( .A(n_458), .Y(n_1115) );
INVx2_ASAP7_75t_SL g1177 ( .A(n_458), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_458), .Y(n_1260) );
OR2x4_ASAP7_75t_L g460 ( .A(n_459), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g625 ( .A(n_459), .Y(n_625) );
BUFx4f_ASAP7_75t_L g639 ( .A(n_459), .Y(n_639) );
BUFx3_ASAP7_75t_L g680 ( .A(n_459), .Y(n_680) );
BUFx3_ASAP7_75t_L g772 ( .A(n_459), .Y(n_772) );
BUFx3_ASAP7_75t_L g735 ( .A(n_460), .Y(n_735) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_460), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1179 ( .A(n_460), .Y(n_1179) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_467), .C(n_469), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_464), .A2(n_470), .B1(n_514), .B2(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g1380 ( .A(n_466), .Y(n_1380) );
NAND3xp33_ASAP7_75t_SL g585 ( .A(n_467), .B(n_586), .C(n_588), .Y(n_585) );
CKINVDCx8_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
CKINVDCx8_ASAP7_75t_R g727 ( .A(n_468), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g947 ( .A(n_468), .B(n_948), .C(n_952), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g1294 ( .A(n_468), .B(n_1295), .C(n_1298), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_474), .B2(n_475), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_471), .A2(n_475), .B1(n_576), .B2(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_471), .A2(n_862), .B1(n_898), .B2(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g950 ( .A(n_471), .Y(n_950) );
AOI222xp33_ASAP7_75t_L g996 ( .A1(n_471), .A2(n_475), .B1(n_997), .B2(n_998), .C1(n_999), .C2(n_1000), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_471), .B(n_1285), .Y(n_1297) );
AOI22xp33_ASAP7_75t_SL g1346 ( .A1(n_471), .A2(n_475), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AND2x2_ASAP7_75t_L g475 ( .A(n_472), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g730 ( .A(n_472), .B(n_473), .Y(n_730) );
AND2x4_ASAP7_75t_L g732 ( .A(n_472), .B(n_476), .Y(n_732) );
AND2x4_ASAP7_75t_L g860 ( .A(n_472), .B(n_473), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_474), .B(n_520), .Y(n_519) );
AOI32xp33_ASAP7_75t_L g861 ( .A1(n_475), .A2(n_848), .A3(n_862), .B1(n_864), .B2(n_866), .Y(n_861) );
INVxp67_ASAP7_75t_L g905 ( .A(n_475), .Y(n_905) );
INVxp67_ASAP7_75t_L g951 ( .A(n_475), .Y(n_951) );
INVx1_ASAP7_75t_L g1296 ( .A(n_475), .Y(n_1296) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g953 ( .A1(n_480), .A2(n_920), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g1293 ( .A1(n_480), .A2(n_1177), .B1(n_1280), .B2(n_1281), .Y(n_1293) );
INVx1_ASAP7_75t_L g737 ( .A(n_481), .Y(n_737) );
INVx2_ASAP7_75t_L g1003 ( .A(n_481), .Y(n_1003) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_481), .Y(n_1059) );
INVx1_ASAP7_75t_L g1122 ( .A(n_481), .Y(n_1122) );
BUFx3_ASAP7_75t_L g688 ( .A(n_482), .Y(n_688) );
INVx1_ASAP7_75t_L g820 ( .A(n_482), .Y(n_820) );
BUFx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g633 ( .A(n_483), .Y(n_633) );
OAI31xp33_ASAP7_75t_SL g583 ( .A1(n_484), .A2(n_584), .A3(n_585), .B(n_590), .Y(n_583) );
INVx1_ASAP7_75t_L g1299 ( .A(n_484), .Y(n_1299) );
OAI31xp33_ASAP7_75t_L g1435 ( .A1(n_484), .A2(n_1436), .A3(n_1438), .B(n_1441), .Y(n_1435) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
AND2x2_ASAP7_75t_SL g739 ( .A(n_485), .B(n_487), .Y(n_739) );
AND2x2_ASAP7_75t_L g868 ( .A(n_485), .B(n_487), .Y(n_868) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_485), .B(n_487), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1181 ( .A(n_485), .B(n_487), .Y(n_1181) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_489), .B(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g621 ( .A(n_489), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g670 ( .A(n_489), .Y(n_670) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_489), .B(n_1753), .Y(n_1752) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g530 ( .A(n_490), .Y(n_530) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AO21x1_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_504), .B(n_527), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_498), .B2(n_499), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g1279 ( .A1(n_495), .A2(n_499), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g672 ( .A(n_497), .Y(n_672) );
BUFx3_ASAP7_75t_L g888 ( .A(n_497), .Y(n_888) );
BUFx6f_ASAP7_75t_L g993 ( .A(n_497), .Y(n_993) );
INVx2_ASAP7_75t_SL g1808 ( .A(n_497), .Y(n_1808) );
INVx4_ASAP7_75t_L g582 ( .A(n_499), .Y(n_582) );
CKINVDCx16_ASAP7_75t_R g766 ( .A(n_499), .Y(n_766) );
INVx3_ASAP7_75t_SL g913 ( .A(n_499), .Y(n_913) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
BUFx3_ASAP7_75t_L g1366 ( .A(n_502), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g1012 ( .A(n_507), .Y(n_1012) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_L g514 ( .A(n_508), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g526 ( .A(n_508), .B(n_522), .Y(n_526) );
AND2x2_ASAP7_75t_L g711 ( .A(n_508), .B(n_552), .Y(n_711) );
INVx8_ASAP7_75t_L g600 ( .A(n_509), .Y(n_600) );
OR2x2_ASAP7_75t_L g717 ( .A(n_509), .B(n_578), .Y(n_717) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .C(n_525), .Y(n_512) );
INVx1_ASAP7_75t_L g918 ( .A(n_514), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_514), .A2(n_516), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
AND2x4_ASAP7_75t_L g577 ( .A(n_515), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g758 ( .A(n_515), .B(n_578), .Y(n_758) );
INVx1_ASAP7_75t_L g1823 ( .A(n_515), .Y(n_1823) );
BUFx3_ASAP7_75t_L g580 ( .A(n_516), .Y(n_580) );
INVx2_ASAP7_75t_L g708 ( .A(n_516), .Y(n_708) );
INVx2_ASAP7_75t_L g850 ( .A(n_516), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g1270 ( .A1(n_516), .A2(n_577), .B1(n_1264), .B2(n_1271), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_516), .A2(n_758), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_517), .B(n_1789), .Y(n_1794) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_523), .Y(n_1289) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_524), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g1283 ( .A(n_525), .B(n_1284), .C(n_1287), .Y(n_1283) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
AOI31xp33_ASAP7_75t_SL g1145 ( .A1(n_527), .A2(n_1146), .A3(n_1149), .B(n_1156), .Y(n_1145) );
AO21x1_ASAP7_75t_L g1278 ( .A1(n_527), .A2(n_1279), .B(n_1282), .Y(n_1278) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI31xp33_ASAP7_75t_L g567 ( .A1(n_528), .A2(n_568), .A3(n_569), .B(n_581), .Y(n_567) );
BUFx3_ASAP7_75t_L g718 ( .A(n_528), .Y(n_718) );
BUFx2_ASAP7_75t_L g855 ( .A(n_528), .Y(n_855) );
OAI31xp33_ASAP7_75t_L g894 ( .A1(n_528), .A2(n_895), .A3(n_896), .B(n_900), .Y(n_894) );
OAI21xp5_ASAP7_75t_L g1004 ( .A1(n_528), .A2(n_1005), .B(n_1013), .Y(n_1004) );
BUFx2_ASAP7_75t_SL g1273 ( .A(n_528), .Y(n_1273) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g1793 ( .A(n_530), .B(n_1794), .Y(n_1793) );
INVxp67_ASAP7_75t_L g1798 ( .A(n_530), .Y(n_1798) );
OAI31xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .A3(n_534), .B(n_562), .Y(n_531) );
INVx1_ASAP7_75t_L g564 ( .A(n_535), .Y(n_564) );
AOI33xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_540), .A3(n_548), .B1(n_553), .B2(n_554), .B3(n_556), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
OAI33xp33_ASAP7_75t_L g1209 ( .A1(n_537), .A2(n_667), .A3(n_1210), .B1(n_1213), .B2(n_1216), .B3(n_1219), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1301 ( .A(n_537), .Y(n_1301) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
INVx2_ASAP7_75t_L g649 ( .A(n_538), .Y(n_649) );
INVx2_ASAP7_75t_L g831 ( .A(n_538), .Y(n_831) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g942 ( .A(n_542), .Y(n_942) );
INVx2_ASAP7_75t_L g1163 ( .A(n_542), .Y(n_1163) );
INVx2_ASAP7_75t_SL g1303 ( .A(n_542), .Y(n_1303) );
INVx1_ASAP7_75t_L g1311 ( .A(n_542), .Y(n_1311) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_543), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g1788 ( .A(n_543), .B(n_1789), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1832 ( .A(n_543), .B(n_1805), .Y(n_1832) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g561 ( .A(n_547), .Y(n_561) );
BUFx6f_ASAP7_75t_L g1165 ( .A(n_547), .Y(n_1165) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g1306 ( .A(n_550), .Y(n_1306) );
AND2x4_ASAP7_75t_L g1820 ( .A(n_550), .B(n_1805), .Y(n_1820) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx3_ASAP7_75t_L g916 ( .A(n_552), .Y(n_916) );
BUFx6f_ASAP7_75t_L g1152 ( .A(n_552), .Y(n_1152) );
AND2x4_ASAP7_75t_SL g1804 ( .A(n_552), .B(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1813 ( .A(n_552), .Y(n_1813) );
AND2x6_ASAP7_75t_L g1816 ( .A(n_552), .B(n_1789), .Y(n_1816) );
INVx2_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
INVx2_ASAP7_75t_L g842 ( .A(n_554), .Y(n_842) );
AOI33xp33_ASAP7_75t_L g1300 ( .A1(n_554), .A2(n_1301), .A3(n_1302), .B1(n_1304), .B2(n_1308), .B3(n_1310), .Y(n_1300) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_554), .B(n_1370), .C(n_1371), .Y(n_1369) );
AND2x4_ASAP7_75t_L g668 ( .A(n_555), .B(n_669), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g931 ( .A1(n_555), .A2(n_794), .B1(n_932), .B2(n_933), .C(n_934), .Y(n_931) );
INVx4_ASAP7_75t_L g1814 ( .A(n_555), .Y(n_1814) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g1368 ( .A(n_558), .Y(n_1368) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_559), .B(n_578), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g1170 ( .A(n_559), .Y(n_1170) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g566 ( .A(n_567), .B(n_583), .C(n_591), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_570), .A2(n_661), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_570), .A2(n_658), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_570), .A2(n_661), .B1(n_1503), .B2(n_1506), .Y(n_1514) );
OAI22xp5_ASAP7_75t_L g1515 ( .A1(n_570), .A2(n_1030), .B1(n_1500), .B2(n_1511), .Y(n_1515) );
OAI22xp5_ASAP7_75t_L g1874 ( .A1(n_570), .A2(n_991), .B1(n_1875), .B2(n_1876), .Y(n_1874) );
INVx5_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_572), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
BUFx2_ASAP7_75t_SL g665 ( .A(n_572), .Y(n_665) );
BUFx3_ASAP7_75t_L g755 ( .A(n_572), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_572), .A2(n_661), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_572), .A2(n_661), .B1(n_1240), .B2(n_1251), .Y(n_1256) );
BUFx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
NAND3xp33_ASAP7_75t_SL g1005 ( .A(n_574), .B(n_1006), .C(n_1008), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1386 ( .A(n_574), .B(n_1387), .C(n_1390), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_579), .B2(n_580), .Y(n_575) );
BUFx3_ASAP7_75t_L g705 ( .A(n_577), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_577), .A2(n_580), .B1(n_898), .B2(n_899), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_577), .A2(n_849), .B1(n_1107), .B2(n_1108), .Y(n_1106) );
INVx1_ASAP7_75t_L g1155 ( .A(n_577), .Y(n_1155) );
AOI222xp33_ASAP7_75t_L g1390 ( .A1(n_577), .A2(n_580), .B1(n_916), .B2(n_1391), .C1(n_1392), .C2(n_1393), .Y(n_1390) );
O2A1O1Ixp33_ASAP7_75t_L g914 ( .A1(n_578), .A2(n_915), .B(n_916), .C(n_917), .Y(n_914) );
INVx1_ASAP7_75t_L g921 ( .A(n_578), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_579), .B(n_587), .Y(n_586) );
AOI222xp33_ASAP7_75t_L g1006 ( .A1(n_580), .A2(n_758), .B1(n_916), .B2(n_999), .C1(n_1000), .C2(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_580), .A2(n_705), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_580), .A2(n_705), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_580), .A2(n_758), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_587), .B(n_1430), .Y(n_1440) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_619), .Y(n_591) );
OAI33xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .A3(n_602), .B1(n_610), .B2(n_614), .B3(n_615), .Y(n_592) );
OAI33xp33_ASAP7_75t_L g886 ( .A1(n_593), .A2(n_842), .A3(n_887), .B1(n_889), .B2(n_890), .B3(n_893), .Y(n_886) );
BUFx6f_ASAP7_75t_L g1022 ( .A(n_593), .Y(n_1022) );
OAI33xp33_ASAP7_75t_L g1512 ( .A1(n_593), .A2(n_667), .A3(n_1513), .B1(n_1514), .B2(n_1515), .B3(n_1516), .Y(n_1512) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_601), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_595), .A2(n_611), .B1(n_624), .B2(n_626), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_596), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_596), .A2(n_812), .B1(n_828), .B2(n_833), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_596), .A2(n_1037), .B1(n_1329), .B2(n_1332), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_596), .A2(n_833), .B1(n_1327), .B2(n_1336), .Y(n_1342) );
OAI22xp33_ASAP7_75t_L g1408 ( .A1(n_596), .A2(n_1037), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
INVx4_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx3_ASAP7_75t_L g652 ( .A(n_597), .Y(n_652) );
BUFx6f_ASAP7_75t_L g1103 ( .A(n_597), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_598), .A2(n_874), .B1(n_884), .B2(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_598), .A2(n_978), .B1(n_983), .B2(n_993), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_598), .A2(n_888), .B1(n_1413), .B2(n_1414), .Y(n_1412) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_SL g617 ( .A(n_600), .Y(n_617) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_600), .Y(n_655) );
INVx4_ASAP7_75t_L g833 ( .A(n_600), .Y(n_833) );
INVx1_ASAP7_75t_L g1037 ( .A(n_600), .Y(n_1037) );
INVx1_ASAP7_75t_L g1254 ( .A(n_600), .Y(n_1254) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_601), .A2(n_613), .B1(n_639), .B2(n_640), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_607), .B2(n_609), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_603), .A2(n_616), .B1(n_629), .B2(n_631), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_604), .A2(n_611), .B1(n_612), .B2(n_613), .Y(n_610) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g658 ( .A(n_605), .Y(n_658) );
BUFx2_ASAP7_75t_L g795 ( .A(n_605), .Y(n_795) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g663 ( .A(n_606), .Y(n_663) );
INVx1_ASAP7_75t_L g836 ( .A(n_606), .Y(n_836) );
BUFx3_ASAP7_75t_L g891 ( .A(n_606), .Y(n_891) );
BUFx2_ASAP7_75t_L g1340 ( .A(n_606), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_607), .A2(n_975), .B1(n_986), .B2(n_991), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_607), .A2(n_835), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_608), .Y(n_612) );
BUFx4f_ASAP7_75t_L g703 ( .A(n_608), .Y(n_703) );
INVx4_ASAP7_75t_L g797 ( .A(n_608), .Y(n_797) );
BUFx4f_ASAP7_75t_L g845 ( .A(n_608), .Y(n_845) );
BUFx4f_ASAP7_75t_L g937 ( .A(n_608), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_609), .A2(n_618), .B1(n_635), .B2(n_636), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_612), .A2(n_835), .B1(n_878), .B2(n_881), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_612), .A2(n_1099), .B1(n_1243), .B2(n_1246), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_612), .A2(n_1326), .B1(n_1335), .B2(n_1340), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_612), .A2(n_891), .B1(n_1416), .B2(n_1417), .Y(n_1415) );
OAI33xp33_ASAP7_75t_L g1404 ( .A1(n_614), .A2(n_1405), .A3(n_1408), .B1(n_1411), .B2(n_1412), .B3(n_1415), .Y(n_1404) );
OAI33xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .A3(n_628), .B1(n_634), .B2(n_637), .B3(n_638), .Y(n_619) );
OAI33xp33_ASAP7_75t_L g810 ( .A1(n_620), .A2(n_637), .A3(n_811), .B1(n_815), .B2(n_822), .B3(n_827), .Y(n_810) );
OAI33xp33_ASAP7_75t_L g872 ( .A1(n_620), .A2(n_637), .A3(n_873), .B1(n_877), .B2(n_880), .B3(n_883), .Y(n_872) );
BUFx3_ASAP7_75t_L g1127 ( .A(n_620), .Y(n_1127) );
OAI33xp33_ASAP7_75t_L g1324 ( .A1(n_620), .A2(n_637), .A3(n_1325), .B1(n_1328), .B2(n_1331), .B3(n_1334), .Y(n_1324) );
OAI33xp33_ASAP7_75t_L g1497 ( .A1(n_620), .A2(n_689), .A3(n_1498), .B1(n_1502), .B2(n_1505), .B3(n_1509), .Y(n_1497) );
BUFx4f_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx4f_ASAP7_75t_L g676 ( .A(n_621), .Y(n_676) );
BUFx2_ASAP7_75t_L g769 ( .A(n_621), .Y(n_769) );
BUFx8_ASAP7_75t_L g1224 ( .A(n_621), .Y(n_1224) );
INVx2_ASAP7_75t_SL g1131 ( .A(n_624), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1141 ( .A1(n_624), .A2(n_1142), .B1(n_1143), .B2(n_1144), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1780 ( .A(n_624), .B(n_1781), .Y(n_1780) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g1078 ( .A(n_625), .Y(n_1078) );
INVx2_ASAP7_75t_L g682 ( .A(n_626), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_626), .A2(n_639), .B1(n_828), .B2(n_829), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_626), .A2(n_639), .B1(n_884), .B2(n_885), .Y(n_883) );
BUFx6f_ASAP7_75t_L g1143 ( .A(n_626), .Y(n_1143) );
HB1xp67_ASAP7_75t_L g1226 ( .A(n_626), .Y(n_1226) );
HB1xp67_ASAP7_75t_L g1241 ( .A(n_626), .Y(n_1241) );
OAI22xp33_ASAP7_75t_L g1331 ( .A1(n_626), .A2(n_639), .B1(n_1332), .B2(n_1333), .Y(n_1331) );
OAI22xp33_ASAP7_75t_L g1424 ( .A1(n_626), .A2(n_639), .B1(n_1410), .B2(n_1417), .Y(n_1424) );
BUFx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_627), .Y(n_642) );
BUFx2_ASAP7_75t_L g697 ( .A(n_627), .Y(n_697) );
INVx2_ASAP7_75t_L g782 ( .A(n_629), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_629), .A2(n_823), .B1(n_824), .B2(n_826), .Y(n_822) );
OAI22xp33_ASAP7_75t_SL g1080 ( .A1(n_629), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_629), .A2(n_636), .B1(n_1326), .B2(n_1327), .Y(n_1325) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx5_ASAP7_75t_L g684 ( .A(n_630), .Y(n_684) );
INVx2_ASAP7_75t_SL g687 ( .A(n_630), .Y(n_687) );
INVx2_ASAP7_75t_SL g1135 ( .A(n_630), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1374 ( .A(n_630), .Y(n_1374) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_631), .A2(n_635), .B1(n_878), .B2(n_879), .Y(n_877) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g636 ( .A(n_632), .Y(n_636) );
CKINVDCx8_ASAP7_75t_R g685 ( .A(n_632), .Y(n_685) );
INVx3_ASAP7_75t_L g982 ( .A(n_632), .Y(n_982) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g825 ( .A(n_633), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_635), .A2(n_688), .B1(n_1215), .B2(n_1222), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_635), .A2(n_688), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_636), .A2(n_687), .B1(n_881), .B2(n_882), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g811 ( .A1(n_639), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_639), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_639), .A2(n_949), .B1(n_974), .B2(n_975), .Y(n_973) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_639), .A2(n_814), .B1(n_985), .B2(n_986), .Y(n_984) );
OAI22xp5_ASAP7_75t_SL g1328 ( .A1(n_639), .A2(n_875), .B1(n_1329), .B2(n_1330), .Y(n_1328) );
OAI22xp33_ASAP7_75t_L g1419 ( .A1(n_639), .A2(n_875), .B1(n_1409), .B2(n_1416), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_640), .A2(n_772), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g726 ( .A(n_641), .Y(n_726) );
INVx2_ASAP7_75t_L g949 ( .A(n_641), .Y(n_949) );
INVx1_ASAP7_75t_L g1117 ( .A(n_641), .Y(n_1117) );
INVx1_ASAP7_75t_L g1501 ( .A(n_641), .Y(n_1501) );
INVx4_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx3_ASAP7_75t_L g775 ( .A(n_642), .Y(n_775) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_642), .Y(n_814) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_642), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1795 ( .A(n_642), .B(n_1752), .Y(n_1795) );
OA21x2_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_740), .B(n_802), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_644), .A2(n_740), .B(n_802), .Y(n_803) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g802 ( .A(n_645), .B(n_741), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_698), .C(n_719), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_675), .Y(n_647) );
OAI33xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .A3(n_656), .B1(n_660), .B2(n_667), .B3(n_671), .Y(n_648) );
OAI33xp33_ASAP7_75t_L g789 ( .A1(n_649), .A2(n_790), .A3(n_793), .B1(n_798), .B2(n_800), .B3(n_801), .Y(n_789) );
OAI33xp33_ASAP7_75t_L g1869 ( .A1(n_649), .A2(n_800), .A3(n_1870), .B1(n_1874), .B2(n_1877), .B3(n_1880), .Y(n_1869) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_651), .A2(n_664), .B1(n_678), .B2(n_681), .Y(n_677) );
INVx2_ASAP7_75t_SL g792 ( .A(n_652), .Y(n_792) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_653), .A2(n_666), .B1(n_678), .B2(n_695), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_654), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_654), .A2(n_771), .B1(n_787), .B2(n_791), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_654), .A2(n_779), .B1(n_784), .B2(n_791), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_654), .A2(n_672), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_654), .A2(n_672), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_654), .A2(n_672), .B1(n_1244), .B2(n_1248), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1485 ( .A1(n_654), .A2(n_672), .B1(n_1454), .B2(n_1459), .Y(n_1485) );
INVx6_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx5_ASAP7_75t_L g930 ( .A(n_655), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_657), .A2(n_673), .B1(n_684), .B2(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g1031 ( .A(n_658), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_658), .A2(n_755), .B1(n_1134), .B2(n_1139), .C(n_1162), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_659), .A2(n_674), .B1(n_687), .B2(n_688), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_661), .A2(n_665), .B1(n_1453), .B2(n_1458), .Y(n_1481) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx4_ASAP7_75t_L g1099 ( .A(n_662), .Y(n_1099) );
INVx4_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_665), .A2(n_1030), .B1(n_1032), .B2(n_1033), .Y(n_1029) );
OAI33xp33_ASAP7_75t_L g1021 ( .A1(n_667), .A2(n_1022), .A3(n_1023), .B1(n_1026), .B2(n_1029), .B3(n_1034), .Y(n_1021) );
OAI33xp33_ASAP7_75t_L g1096 ( .A1(n_667), .A2(n_1022), .A3(n_1097), .B1(n_1098), .B2(n_1100), .B3(n_1101), .Y(n_1096) );
OAI33xp33_ASAP7_75t_L g1252 ( .A1(n_667), .A2(n_1022), .A3(n_1253), .B1(n_1255), .B2(n_1256), .B3(n_1257), .Y(n_1252) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_668), .Y(n_800) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_672), .A2(n_1035), .B1(n_1036), .B2(n_1038), .Y(n_1034) );
OAI33xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .A3(n_683), .B1(n_686), .B2(n_689), .B3(n_694), .Y(n_675) );
OAI33xp33_ASAP7_75t_L g1074 ( .A1(n_676), .A2(n_1075), .A3(n_1080), .B1(n_1085), .B2(n_1090), .B3(n_1093), .Y(n_1074) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_678), .A2(n_1499), .B1(n_1500), .B2(n_1501), .Y(n_1498) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g1232 ( .A(n_680), .Y(n_1232) );
INVx1_ASAP7_75t_L g1886 ( .A(n_680), .Y(n_1886) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx3_ASAP7_75t_L g778 ( .A(n_684), .Y(n_778) );
INVx8_ASAP7_75t_L g1087 ( .A(n_684), .Y(n_1087) );
OAI22xp33_ASAP7_75t_SL g1420 ( .A1(n_684), .A2(n_819), .B1(n_1406), .B2(n_1413), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_685), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_685), .A2(n_929), .B1(n_936), .B2(n_966), .C(n_968), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_685), .A2(n_1086), .B1(n_1088), .B2(n_1089), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_685), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1245) );
OAI22xp33_ASAP7_75t_L g1888 ( .A1(n_685), .A2(n_959), .B1(n_1875), .B2(n_1881), .Y(n_1888) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_687), .A2(n_819), .B1(n_1335), .B2(n_1336), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_688), .A2(n_781), .B1(n_783), .B2(n_784), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_688), .A2(n_1027), .B1(n_1035), .B2(n_1043), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_688), .A2(n_1028), .B1(n_1038), .B2(n_1045), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_688), .A2(n_1214), .B1(n_1221), .B2(n_1228), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1451 ( .A1(n_688), .A2(n_1452), .B1(n_1453), .B2(n_1454), .C(n_1455), .Y(n_1451) );
OAI221xp5_ASAP7_75t_L g1457 ( .A1(n_688), .A2(n_959), .B1(n_1458), .B2(n_1459), .C(n_1460), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_688), .A2(n_1506), .B1(n_1507), .B2(n_1508), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g1768 ( .A1(n_688), .A2(n_1769), .B1(n_1770), .B2(n_1772), .Y(n_1768) );
OAI221xp5_ASAP7_75t_L g1776 ( .A1(n_688), .A2(n_781), .B1(n_1777), .B2(n_1778), .C(n_1779), .Y(n_1776) );
OAI22xp5_ASAP7_75t_L g1889 ( .A1(n_688), .A2(n_1452), .B1(n_1876), .B2(n_1882), .Y(n_1889) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_690), .Y(n_785) );
INVx2_ASAP7_75t_L g1462 ( .A(n_690), .Y(n_1462) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g1092 ( .A(n_691), .Y(n_1092) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g1758 ( .A(n_693), .Y(n_1758) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_695), .A2(n_772), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g1048 ( .A(n_697), .Y(n_1048) );
INVx1_ASAP7_75t_L g1062 ( .A(n_697), .Y(n_1062) );
OAI31xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .A3(n_712), .B(n_718), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g1877 ( .A1(n_703), .A2(n_991), .B1(n_1878), .B2(n_1879), .Y(n_1877) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_709), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_705), .A2(n_849), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_706), .A2(n_729), .B1(n_731), .B2(n_733), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_707), .A2(n_748), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g1865 ( .A(n_708), .Y(n_1865) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g756 ( .A(n_711), .Y(n_756) );
AOI211xp5_ASAP7_75t_L g1149 ( .A1(n_711), .A2(n_1150), .B(n_1153), .C(n_1154), .Y(n_1149) );
INVx3_ASAP7_75t_L g1193 ( .A(n_711), .Y(n_1193) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g761 ( .A(n_714), .Y(n_761) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1110 ( .A(n_716), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_716), .A2(n_1010), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
INVx1_ASAP7_75t_L g1434 ( .A(n_716), .Y(n_1434) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx2_ASAP7_75t_L g764 ( .A(n_717), .Y(n_764) );
INVx1_ASAP7_75t_L g853 ( .A(n_717), .Y(n_853) );
OAI31xp33_ASAP7_75t_L g751 ( .A1(n_718), .A2(n_752), .A3(n_760), .B(n_765), .Y(n_751) );
OAI31xp33_ASAP7_75t_L g1049 ( .A1(n_718), .A2(n_1050), .A3(n_1054), .B(n_1055), .Y(n_1049) );
OAI31xp33_ASAP7_75t_SL g1104 ( .A1(n_718), .A2(n_1105), .A3(n_1109), .B(n_1111), .Y(n_1104) );
OAI31xp33_ASAP7_75t_L g1488 ( .A1(n_718), .A2(n_1489), .A3(n_1490), .B(n_1495), .Y(n_1488) );
OAI31xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_725), .A3(n_734), .B(n_738), .Y(n_719) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g745 ( .A(n_724), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_724), .A2(n_1147), .B1(n_1148), .B2(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1437 ( .A(n_724), .Y(n_1437) );
INVx1_ASAP7_75t_L g1860 ( .A(n_724), .Y(n_1860) );
OAI22xp33_ASAP7_75t_L g1093 ( .A1(n_726), .A2(n_1077), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1230 ( .A1(n_726), .A2(n_1212), .B1(n_1218), .B2(n_1231), .Y(n_1230) );
NAND3xp33_ASAP7_75t_L g1398 ( .A(n_727), .B(n_1399), .C(n_1400), .Y(n_1398) );
NAND3xp33_ASAP7_75t_L g1438 ( .A(n_727), .B(n_1439), .C(n_1440), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_729), .A2(n_731), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_729), .A2(n_731), .B1(n_1052), .B2(n_1064), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_729), .A2(n_731), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
BUFx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx3_ASAP7_75t_L g1205 ( .A(n_730), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_731), .A2(n_1195), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_731), .A2(n_1205), .B1(n_1467), .B2(n_1474), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_731), .A2(n_1205), .B1(n_1493), .B2(n_1521), .Y(n_1520) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g1118 ( .A1(n_732), .A2(n_860), .B1(n_1107), .B2(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1175 ( .A(n_732), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_732), .A2(n_860), .B1(n_1429), .B2(n_1432), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1856 ( .A1(n_732), .A2(n_860), .B1(n_1857), .B2(n_1858), .Y(n_1856) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI31xp33_ASAP7_75t_L g743 ( .A1(n_738), .A2(n_744), .A3(n_746), .B(n_750), .Y(n_743) );
OAI31xp33_ASAP7_75t_L g1056 ( .A1(n_738), .A2(n_1057), .A3(n_1060), .B(n_1065), .Y(n_1056) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g945 ( .A1(n_739), .A2(n_946), .B(n_956), .Y(n_945) );
OAI31xp33_ASAP7_75t_L g1200 ( .A1(n_739), .A2(n_1201), .A3(n_1203), .B(n_1207), .Y(n_1200) );
OAI31xp33_ASAP7_75t_L g1470 ( .A1(n_739), .A2(n_1471), .A3(n_1472), .B(n_1475), .Y(n_1470) );
OAI31xp33_ASAP7_75t_L g1517 ( .A1(n_739), .A2(n_1518), .A3(n_1519), .B(n_1522), .Y(n_1517) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_751), .C(n_767), .Y(n_742) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g1166 ( .A1(n_755), .A2(n_1132), .B1(n_1144), .B2(n_1167), .C(n_1169), .Y(n_1166) );
BUFx2_ASAP7_75t_L g1491 ( .A(n_755), .Y(n_1491) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_758), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_758), .A2(n_849), .B1(n_1347), .B2(n_1354), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1863 ( .A1(n_758), .A2(n_1857), .B1(n_1864), .B2(n_1865), .Y(n_1863) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_764), .Y(n_1198) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_789), .Y(n_767) );
OAI33xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .A3(n_776), .B1(n_780), .B2(n_785), .B3(n_786), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_769), .A2(n_785), .B1(n_957), .B2(n_965), .Y(n_956) );
OAI33xp33_ASAP7_75t_L g1039 ( .A1(n_769), .A2(n_785), .A3(n_1040), .B1(n_1042), .B2(n_1044), .B3(n_1046), .Y(n_1039) );
OAI33xp33_ASAP7_75t_L g1883 ( .A1(n_769), .A2(n_1462), .A3(n_1884), .B1(n_1888), .B2(n_1889), .B3(n_1890), .Y(n_1883) );
OAI22xp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_770) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_772), .A2(n_1024), .B1(n_1032), .B2(n_1041), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1046 ( .A1(n_772), .A2(n_1025), .B1(n_1033), .B2(n_1047), .Y(n_1046) );
OAI22xp33_ASAP7_75t_L g1225 ( .A1(n_772), .A2(n_1211), .B1(n_1217), .B2(n_1226), .Y(n_1225) );
OAI22xp33_ASAP7_75t_L g1238 ( .A1(n_772), .A2(n_1239), .B1(n_1240), .B2(n_1241), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1509 ( .A1(n_772), .A2(n_1143), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_773), .A2(n_788), .B1(n_794), .B2(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx3_ASAP7_75t_L g875 ( .A(n_775), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_777), .A2(n_783), .B1(n_794), .B2(n_796), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_778), .A2(n_1083), .B1(n_1243), .B2(n_1244), .Y(n_1242) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI33xp33_ASAP7_75t_L g1223 ( .A1(n_785), .A2(n_1224), .A3(n_1225), .B1(n_1227), .B2(n_1229), .B3(n_1230), .Y(n_1223) );
OAI33xp33_ASAP7_75t_L g1237 ( .A1(n_785), .A2(n_1224), .A3(n_1238), .B1(n_1242), .B2(n_1245), .B3(n_1249), .Y(n_1237) );
OAI22xp33_ASAP7_75t_L g1513 ( .A1(n_791), .A2(n_1254), .B1(n_1499), .B2(n_1510), .Y(n_1513) );
OAI221xp5_ASAP7_75t_L g1825 ( .A1(n_791), .A2(n_1774), .B1(n_1809), .B2(n_1826), .C(n_1827), .Y(n_1825) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_794), .A2(n_845), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
INVx4_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_797), .Y(n_799) );
INVx2_ASAP7_75t_L g837 ( .A(n_797), .Y(n_837) );
INVx2_ASAP7_75t_L g892 ( .A(n_797), .Y(n_892) );
INVx1_ASAP7_75t_L g932 ( .A(n_797), .Y(n_932) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_799), .A2(n_1081), .B1(n_1088), .B2(n_1099), .Y(n_1098) );
OAI22xp5_ASAP7_75t_SL g1160 ( .A1(n_800), .A2(n_831), .B1(n_1161), .B2(n_1166), .Y(n_1160) );
OA33x2_ASAP7_75t_L g1477 ( .A1(n_800), .A2(n_1022), .A3(n_1478), .B1(n_1481), .B2(n_1482), .B3(n_1485), .Y(n_1477) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_908), .Y(n_805) );
XNOR2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_869), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_843), .C(n_856), .Y(n_808) );
NOR2xp33_ASAP7_75t_SL g809 ( .A(n_810), .B(n_830), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_813), .A2(n_829), .B1(n_835), .B2(n_837), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g1128 ( .A1(n_814), .A2(n_1129), .B1(n_1130), .B2(n_1132), .Y(n_1128) );
INVx1_ASAP7_75t_L g1855 ( .A(n_814), .Y(n_1855) );
OAI22xp33_ASAP7_75t_L g1890 ( .A1(n_814), .A2(n_1873), .B1(n_1879), .B2(n_1885), .Y(n_1890) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_821), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_816), .A2(n_823), .B1(n_835), .B2(n_837), .Y(n_834) );
INVx2_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
INVx3_ASAP7_75t_L g980 ( .A(n_818), .Y(n_980) );
INVx2_ASAP7_75t_SL g1138 ( .A(n_818), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1750 ( .A(n_818), .B(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_820), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_821), .A2(n_826), .B1(n_833), .B2(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_824), .A2(n_966), .B1(n_977), .B2(n_978), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_824), .A2(n_1138), .B1(n_1139), .B2(n_1140), .Y(n_1137) );
BUFx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g1423 ( .A(n_825), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1786 ( .A(n_825), .B(n_1752), .Y(n_1786) );
OAI33xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .A3(n_834), .B1(n_838), .B2(n_839), .B3(n_842), .Y(n_830) );
OAI33xp33_ASAP7_75t_L g987 ( .A1(n_831), .A2(n_842), .A3(n_988), .B1(n_989), .B2(n_990), .B3(n_992), .Y(n_987) );
OAI33xp33_ASAP7_75t_L g1337 ( .A1(n_831), .A2(n_842), .A3(n_1338), .B1(n_1339), .B2(n_1341), .B3(n_1342), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_833), .A2(n_879), .B1(n_882), .B2(n_888), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_833), .A2(n_888), .B1(n_974), .B2(n_985), .Y(n_988) );
INVx2_ASAP7_75t_L g1810 ( .A(n_833), .Y(n_1810) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_835), .A2(n_837), .B1(n_1330), .B2(n_1333), .Y(n_1341) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g991 ( .A(n_836), .Y(n_991) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI31xp33_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_851), .A3(n_854), .B(n_855), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_845), .A2(n_891), .B1(n_977), .B2(n_981), .Y(n_989) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g1159 ( .A(n_852), .Y(n_1159) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_SL g923 ( .A(n_853), .B(n_924), .Y(n_923) );
OAI31xp33_ASAP7_75t_L g1191 ( .A1(n_855), .A2(n_1192), .A3(n_1197), .B(n_1199), .Y(n_1191) );
OAI31xp33_ASAP7_75t_SL g1350 ( .A1(n_855), .A2(n_1351), .A3(n_1352), .B(n_1355), .Y(n_1350) );
OAI31xp33_ASAP7_75t_L g1425 ( .A1(n_855), .A2(n_1426), .A3(n_1427), .B(n_1433), .Y(n_1425) );
OAI31xp33_ASAP7_75t_SL g1463 ( .A1(n_855), .A2(n_1464), .A3(n_1465), .B(n_1469), .Y(n_1463) );
OAI31xp33_ASAP7_75t_SL g856 ( .A1(n_857), .A2(n_858), .A3(n_867), .B(n_868), .Y(n_856) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g1764 ( .A(n_863), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_864), .B(n_1757), .Y(n_1756) );
INVx3_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OAI31xp33_ASAP7_75t_SL g901 ( .A1(n_868), .A2(n_902), .A3(n_903), .B(n_904), .Y(n_901) );
OAI21xp5_ASAP7_75t_L g994 ( .A1(n_868), .A2(n_995), .B(n_1001), .Y(n_994) );
OAI31xp33_ASAP7_75t_L g1343 ( .A1(n_868), .A2(n_1344), .A3(n_1345), .B(n_1349), .Y(n_1343) );
OAI21xp5_ASAP7_75t_L g1395 ( .A1(n_868), .A2(n_1396), .B(n_1398), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_894), .C(n_901), .Y(n_870) );
NOR2xp33_ASAP7_75t_SL g871 ( .A(n_872), .B(n_886), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_876), .A2(n_885), .B1(n_891), .B2(n_892), .Y(n_890) );
INVx2_ASAP7_75t_L g1168 ( .A(n_891), .Y(n_1168) );
XOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_969), .Y(n_908) );
OAI21xp5_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_943), .B(n_945), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_916), .B(n_1432), .Y(n_1431) );
OAI21xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_931), .B(n_935), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B1(n_929), .B2(n_930), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_928), .A2(n_930), .B1(n_1076), .B2(n_1094), .Y(n_1097) );
OAI22xp33_ASAP7_75t_L g1478 ( .A1(n_928), .A2(n_930), .B1(n_1479), .B2(n_1480), .Y(n_1478) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_930), .A2(n_1082), .B1(n_1089), .B2(n_1102), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g1870 ( .A1(n_930), .A2(n_1871), .B1(n_1872), .B2(n_1873), .Y(n_1870) );
OAI22xp5_ASAP7_75t_L g1880 ( .A1(n_930), .A2(n_1807), .B1(n_1881), .B2(n_1882), .Y(n_1880) );
OAI211xp5_ASAP7_75t_SL g935 ( .A1(n_936), .A2(n_937), .B(n_938), .C(n_941), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_937), .A2(n_1079), .B1(n_1095), .B2(n_1099), .Y(n_1100) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx3_ASAP7_75t_L g1828 ( .A(n_940), .Y(n_1828) );
INVx1_ASAP7_75t_L g1835 ( .A(n_943), .Y(n_1835) );
BUFx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NAND2xp5_ASAP7_75t_SL g946 ( .A(n_947), .B(n_953), .Y(n_946) );
INVx1_ASAP7_75t_L g1066 ( .A(n_954), .Y(n_1066) );
OAI211xp5_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_959), .B(n_961), .C(n_963), .Y(n_957) );
INVx2_ASAP7_75t_SL g959 ( .A(n_960), .Y(n_959) );
AND2x4_ASAP7_75t_L g1766 ( .A(n_962), .B(n_1757), .Y(n_1766) );
BUFx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx3_ASAP7_75t_L g1319 ( .A(n_967), .Y(n_1319) );
INVx1_ASAP7_75t_L g1771 ( .A(n_967), .Y(n_1771) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_994), .C(n_1004), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_972), .B(n_987), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1421 ( .A1(n_980), .A2(n_1407), .B1(n_1414), .B2(n_1422), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_982), .A2(n_1134), .B1(n_1135), .B2(n_1136), .Y(n_1133) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_1003), .A2(n_1157), .B1(n_1158), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1003), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_1003), .A2(n_1179), .B1(n_1388), .B2(n_1389), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1011), .B2(n_1012), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_1010), .A2(n_1157), .B1(n_1158), .B2(n_1159), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1016), .B1(n_1184), .B2(n_1523), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
XNOR2xp5_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1067), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
NAND3xp33_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1049), .C(n_1056), .Y(n_1019) );
NOR2xp33_ASAP7_75t_SL g1020 ( .A(n_1021), .B(n_1039), .Y(n_1020) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_1036), .A2(n_1220), .B1(n_1221), .B2(n_1222), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_1036), .A2(n_1220), .B1(n_1504), .B2(n_1508), .Y(n_1516) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1075 ( .A1(n_1047), .A2(n_1076), .B1(n_1077), .B2(n_1079), .Y(n_1075) );
INVxp67_ASAP7_75t_SL g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1048), .Y(n_1262) );
INVxp67_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1062), .Y(n_1887) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1124), .B1(n_1182), .B2(n_1183), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_1071), .Y(n_1182) );
NAND3xp33_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1104), .C(n_1112), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1096), .Y(n_1073) );
BUFx4f_ASAP7_75t_SL g1077 ( .A(n_1078), .Y(n_1077) );
INVx3_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1507 ( .A(n_1087), .Y(n_1507) );
OAI33xp33_ASAP7_75t_L g1126 ( .A1(n_1090), .A2(n_1127), .A3(n_1128), .B1(n_1133), .B2(n_1137), .B3(n_1141), .Y(n_1126) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
BUFx2_ASAP7_75t_L g1383 ( .A(n_1092), .Y(n_1383) );
OAI22xp33_ASAP7_75t_L g1253 ( .A1(n_1102), .A2(n_1239), .B1(n_1250), .B2(n_1254), .Y(n_1253) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1103), .Y(n_1220) );
INVx3_ASAP7_75t_L g1872 ( .A(n_1103), .Y(n_1872) );
OAI31xp33_ASAP7_75t_L g1112 ( .A1(n_1113), .A2(n_1116), .A3(n_1120), .B(n_1123), .Y(n_1112) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
OAI31xp33_ASAP7_75t_L g1258 ( .A1(n_1123), .A2(n_1259), .A3(n_1261), .B(n_1266), .Y(n_1258) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1124), .Y(n_1183) );
NOR4xp25_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1145), .C(n_1160), .D(n_1171), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_1127), .A2(n_1451), .B1(n_1457), .B2(n_1462), .Y(n_1450) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1135), .Y(n_1314) );
OAI22xp5_ASAP7_75t_L g1773 ( .A1(n_1143), .A2(n_1231), .B1(n_1774), .B2(n_1775), .Y(n_1773) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
BUFx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1834 ( .A(n_1165), .B(n_1805), .Y(n_1834) );
INVx3_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
AOI31xp33_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1176), .A3(n_1178), .B(n_1180), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1397 ( .A(n_1177), .Y(n_1397) );
INVx2_ASAP7_75t_L g1476 ( .A(n_1179), .Y(n_1476) );
CKINVDCx14_ASAP7_75t_R g1180 ( .A(n_1181), .Y(n_1180) );
OAI31xp33_ASAP7_75t_L g1851 ( .A1(n_1181), .A2(n_1852), .A3(n_1853), .B(n_1859), .Y(n_1851) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1184), .Y(n_1523) );
XNOR2xp5_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1357), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1187), .B1(n_1274), .B2(n_1356), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1189), .B1(n_1233), .B2(n_1234), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
NAND3xp33_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1200), .C(n_1208), .Y(n_1190) );
NAND3xp33_ASAP7_75t_L g1427 ( .A(n_1193), .B(n_1428), .C(n_1431), .Y(n_1427) );
NOR2xp33_ASAP7_75t_SL g1208 ( .A(n_1209), .B(n_1223), .Y(n_1208) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND3xp33_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1258), .C(n_1267), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1252), .Y(n_1236) );
OAI31xp33_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1269), .A3(n_1272), .B(n_1273), .Y(n_1267) );
OAI21xp5_ASAP7_75t_L g1385 ( .A1(n_1273), .A2(n_1386), .B(n_1394), .Y(n_1385) );
OAI31xp33_ASAP7_75t_L g1861 ( .A1(n_1273), .A2(n_1862), .A3(n_1866), .B(n_1867), .Y(n_1861) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1274), .Y(n_1356) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
XNOR2x1_ASAP7_75t_SL g1275 ( .A(n_1276), .B(n_1321), .Y(n_1275) );
NAND4xp75_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1292), .C(n_1300), .D(n_1312), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1291), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1290), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1289), .Y(n_1307) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1289), .Y(n_1309) );
AO21x1_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1294), .B(n_1299), .Y(n_1292) );
NAND3xp33_ASAP7_75t_L g1362 ( .A(n_1301), .B(n_1363), .C(n_1367), .Y(n_1362) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1301), .Y(n_1411) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
BUFx2_ASAP7_75t_L g1461 ( .A(n_1317), .Y(n_1461) );
INVx2_ASAP7_75t_L g1452 ( .A(n_1319), .Y(n_1452) );
AND3x1_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1343), .C(n_1350), .Y(n_1322) );
NOR2xp33_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1337), .Y(n_1323) );
XNOR2xp5_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1446), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_1359), .A2(n_1401), .B1(n_1444), .B2(n_1445), .Y(n_1358) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1359), .Y(n_1444) );
NAND3xp33_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1385), .C(n_1395), .Y(n_1360) );
AND4x1_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1369), .C(n_1372), .D(n_1381), .Y(n_1361) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
BUFx2_ASAP7_75t_L g1456 ( .A(n_1379), .Y(n_1456) );
NAND3xp33_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1383), .C(n_1384), .Y(n_1381) );
INVx3_ASAP7_75t_SL g1445 ( .A(n_1401), .Y(n_1445) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1402), .Y(n_1443) );
NAND3xp33_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1425), .C(n_1435), .Y(n_1402) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1418), .Y(n_1403) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
XNOR2x1_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1486), .Y(n_1446) );
NAND4xp75_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1463), .C(n_1470), .D(n_1477), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
AND3x1_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1496), .C(n_1517), .Y(n_1487) );
NOR2xp33_ASAP7_75t_SL g1496 ( .A(n_1497), .B(n_1512), .Y(n_1496) );
OAI221xp5_ASAP7_75t_L g1524 ( .A1(n_1525), .A2(n_1739), .B1(n_1741), .B2(n_1837), .C(n_1841), .Y(n_1524) );
AOI21xp5_ASAP7_75t_L g1525 ( .A1(n_1526), .A2(n_1665), .B(n_1713), .Y(n_1525) );
NAND5xp2_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1615), .C(n_1631), .D(n_1644), .E(n_1657), .Y(n_1526) );
AOI211xp5_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1559), .B(n_1574), .C(n_1599), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1545), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1529), .B(n_1626), .Y(n_1691) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_1530), .Y(n_1529) );
OR2x2_ASAP7_75t_L g1617 ( .A(n_1530), .B(n_1583), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1530), .B(n_1626), .Y(n_1625) );
AOI322xp5_ASAP7_75t_L g1644 ( .A1(n_1530), .A2(n_1601), .A3(n_1645), .B1(n_1649), .B2(n_1650), .C1(n_1654), .C2(n_1655), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1530), .B(n_1684), .Y(n_1683) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1530), .B(n_1701), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1729 ( .A(n_1530), .B(n_1591), .Y(n_1729) );
O2A1O1Ixp33_ASAP7_75t_SL g1735 ( .A1(n_1530), .A2(n_1585), .B(n_1600), .C(n_1685), .Y(n_1735) );
INVx4_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
INVx4_ASAP7_75t_L g1581 ( .A(n_1531), .Y(n_1581) );
NAND2xp5_ASAP7_75t_SL g1590 ( .A(n_1531), .B(n_1547), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1531), .B(n_1619), .Y(n_1618) );
NOR2xp33_ASAP7_75t_L g1634 ( .A(n_1531), .B(n_1566), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1653 ( .A(n_1531), .B(n_1547), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1654 ( .A(n_1531), .B(n_1552), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1680 ( .A(n_1531), .B(n_1660), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1531), .B(n_1620), .Y(n_1712) );
AOI321xp33_ASAP7_75t_R g1724 ( .A1(n_1531), .A2(n_1559), .A3(n_1618), .B1(n_1630), .B2(n_1649), .C(n_1725), .Y(n_1724) );
AND2x4_ASAP7_75t_SL g1531 ( .A(n_1532), .B(n_1540), .Y(n_1531) );
AND2x4_ASAP7_75t_L g1533 ( .A(n_1534), .B(n_1535), .Y(n_1533) );
AND2x6_ASAP7_75t_L g1538 ( .A(n_1534), .B(n_1539), .Y(n_1538) );
AND2x6_ASAP7_75t_L g1541 ( .A(n_1534), .B(n_1542), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1534), .B(n_1544), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1534), .B(n_1544), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1534), .B(n_1544), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1534), .B(n_1535), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1537), .Y(n_1535) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1538), .Y(n_1612) );
HB1xp67_ASAP7_75t_L g1894 ( .A(n_1539), .Y(n_1894) );
AOI221xp5_ASAP7_75t_L g1733 ( .A1(n_1545), .A2(n_1675), .B1(n_1698), .B2(n_1734), .C(n_1735), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1551), .Y(n_1545) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1546), .B(n_1552), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1546), .B(n_1620), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1685 ( .A(n_1546), .B(n_1585), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1715 ( .A(n_1546), .B(n_1664), .Y(n_1715) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1633 ( .A(n_1547), .B(n_1556), .Y(n_1633) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1547), .B(n_1553), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1547), .B(n_1591), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1547), .B(n_1643), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1547), .B(n_1621), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1732 ( .A(n_1547), .B(n_1621), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1549), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1548), .B(n_1549), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1551), .B(n_1625), .Y(n_1624) );
NAND3xp33_ASAP7_75t_L g1678 ( .A(n_1551), .B(n_1670), .C(n_1679), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_1551), .B(n_1677), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1551), .B(n_1589), .Y(n_1723) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
OR2x2_ASAP7_75t_L g1673 ( .A(n_1552), .B(n_1653), .Y(n_1673) );
OR2x2_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1556), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1553), .B(n_1586), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1553), .B(n_1556), .Y(n_1591) );
INVx2_ASAP7_75t_L g1621 ( .A(n_1553), .Y(n_1621) );
NAND2x1p5_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1555), .Y(n_1553) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1556), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1556), .B(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1556), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1702 ( .A(n_1556), .B(n_1584), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
AOI221xp5_ASAP7_75t_L g1714 ( .A1(n_1559), .A2(n_1604), .B1(n_1715), .B2(n_1716), .C(n_1717), .Y(n_1714) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
OR2x2_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1566), .Y(n_1560) );
AOI221xp5_ASAP7_75t_L g1615 ( .A1(n_1561), .A2(n_1601), .B1(n_1616), .B2(n_1618), .C(n_1622), .Y(n_1615) );
AOI221xp5_ASAP7_75t_L g1631 ( .A1(n_1561), .A2(n_1632), .B1(n_1634), .B2(n_1635), .C(n_1640), .Y(n_1631) );
OAI322xp33_ASAP7_75t_L g1689 ( .A1(n_1561), .A2(n_1584), .A3(n_1690), .B1(n_1692), .B2(n_1693), .C1(n_1694), .C2(n_1695), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1561), .B(n_1677), .Y(n_1711) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx3_ASAP7_75t_L g1577 ( .A(n_1562), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1562), .B(n_1594), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1562), .B(n_1570), .Y(n_1629) );
OR2x2_ASAP7_75t_L g1661 ( .A(n_1562), .B(n_1570), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1564), .Y(n_1562) );
AOI21xp33_ASAP7_75t_L g1738 ( .A1(n_1566), .A2(n_1617), .B(n_1638), .Y(n_1738) );
OR2x2_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1570), .Y(n_1566) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1567), .Y(n_1582) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1567), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
A2O1A1Ixp33_ASAP7_75t_L g1587 ( .A1(n_1570), .A2(n_1588), .B(n_1592), .C(n_1596), .Y(n_1587) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1570), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1570), .B(n_1577), .Y(n_1601) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_1570), .B(n_1598), .Y(n_1627) );
OAI22xp5_ASAP7_75t_L g1635 ( .A1(n_1570), .A2(n_1636), .B1(n_1637), .B2(n_1638), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1570), .B(n_1582), .Y(n_1649) );
INVx2_ASAP7_75t_L g1670 ( .A(n_1570), .Y(n_1670) );
INVx2_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
OR2x2_ASAP7_75t_L g1663 ( .A(n_1571), .B(n_1598), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1587), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1578), .Y(n_1575) );
CKINVDCx14_ASAP7_75t_R g1576 ( .A(n_1577), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1656 ( .A(n_1577), .B(n_1582), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1688 ( .A(n_1577), .B(n_1597), .Y(n_1688) );
OR2x2_ASAP7_75t_L g1693 ( .A(n_1577), .B(n_1582), .Y(n_1693) );
OR2x2_ASAP7_75t_L g1694 ( .A(n_1577), .B(n_1627), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1577), .B(n_1626), .Y(n_1698) );
O2A1O1Ixp33_ASAP7_75t_SL g1717 ( .A1(n_1577), .A2(n_1648), .B(n_1718), .C(n_1720), .Y(n_1717) );
OR2x2_ASAP7_75t_L g1731 ( .A(n_1577), .B(n_1663), .Y(n_1731) );
A2O1A1Ixp33_ASAP7_75t_R g1736 ( .A1(n_1577), .A2(n_1691), .B(n_1737), .C(n_1738), .Y(n_1736) );
AOI221xp5_ASAP7_75t_L g1666 ( .A1(n_1578), .A2(n_1601), .B1(n_1627), .B2(n_1667), .C(n_1672), .Y(n_1666) );
NOR2xp33_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1583), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
OAI21xp33_ASAP7_75t_L g1628 ( .A1(n_1580), .A2(n_1629), .B(n_1630), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1582), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1581), .B(n_1605), .Y(n_1604) );
NOR2x1_ASAP7_75t_L g1664 ( .A(n_1581), .B(n_1647), .Y(n_1664) );
NAND2x1_ASAP7_75t_L g1668 ( .A(n_1581), .B(n_1639), .Y(n_1668) );
CKINVDCx5p33_ASAP7_75t_R g1677 ( .A(n_1581), .Y(n_1677) );
NOR2xp33_ASAP7_75t_L g1719 ( .A(n_1581), .B(n_1594), .Y(n_1719) );
INVx2_ASAP7_75t_L g1660 ( .A(n_1582), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1582), .B(n_1677), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_1583), .B(n_1633), .Y(n_1632) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1585), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1584), .B(n_1620), .Y(n_1630) );
OR2x2_ASAP7_75t_L g1646 ( .A(n_1584), .B(n_1647), .Y(n_1646) );
AOI321xp33_ASAP7_75t_L g1708 ( .A1(n_1584), .A2(n_1606), .A3(n_1655), .B1(n_1709), .B2(n_1711), .C(n_1712), .Y(n_1708) );
OAI221xp5_ASAP7_75t_L g1599 ( .A1(n_1585), .A2(n_1600), .B1(n_1602), .B2(n_1603), .C(n_1606), .Y(n_1599) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1585), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1585), .B(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1588), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1591), .Y(n_1588) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1591), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1591), .B(n_1652), .Y(n_1651) );
OAI31xp33_ASAP7_75t_L g1657 ( .A1(n_1592), .A2(n_1658), .A3(n_1662), .B(n_1664), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1595), .Y(n_1592) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1593), .Y(n_1602) );
AOI221xp5_ASAP7_75t_L g1697 ( .A1(n_1593), .A2(n_1698), .B1(n_1699), .B2(n_1703), .C(n_1704), .Y(n_1697) );
OAI22xp5_ASAP7_75t_L g1667 ( .A1(n_1594), .A2(n_1668), .B1(n_1669), .B2(n_1671), .Y(n_1667) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1595), .Y(n_1707) );
OAI211xp5_ASAP7_75t_L g1622 ( .A1(n_1596), .A2(n_1623), .B(n_1624), .C(n_1628), .Y(n_1622) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1597), .B(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
NOR2xp33_ASAP7_75t_L g1721 ( .A(n_1598), .B(n_1722), .Y(n_1721) );
A2O1A1Ixp33_ASAP7_75t_L g1726 ( .A1(n_1598), .A2(n_1629), .B(n_1664), .C(n_1686), .Y(n_1726) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1601), .B(n_1676), .Y(n_1734) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVx2_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
OAI221xp5_ASAP7_75t_L g1609 ( .A1(n_1610), .A2(n_1611), .B1(n_1612), .B2(n_1613), .C(n_1614), .Y(n_1609) );
CKINVDCx20_ASAP7_75t_R g1740 ( .A(n_1612), .Y(n_1740) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1620), .B(n_1652), .Y(n_1671) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1620), .Y(n_1710) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1625), .Y(n_1636) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1625), .B(n_1642), .Y(n_1641) );
CKINVDCx5p33_ASAP7_75t_R g1626 ( .A(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1633), .Y(n_1737) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1637), .Y(n_1675) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVxp67_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1642), .Y(n_1648) );
NAND2xp5_ASAP7_75t_SL g1645 ( .A(n_1646), .B(n_1648), .Y(n_1645) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1646), .Y(n_1703) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
OAI211xp5_ASAP7_75t_L g1727 ( .A1(n_1652), .A2(n_1728), .B(n_1730), .C(n_1732), .Y(n_1727) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
OR2x2_ASAP7_75t_L g1659 ( .A(n_1660), .B(n_1661), .Y(n_1659) );
CKINVDCx5p33_ASAP7_75t_R g1662 ( .A(n_1663), .Y(n_1662) );
OAI211xp5_ASAP7_75t_L g1672 ( .A1(n_1663), .A2(n_1673), .B(n_1674), .C(n_1678), .Y(n_1672) );
NAND4xp25_ASAP7_75t_L g1665 ( .A(n_1666), .B(n_1681), .C(n_1697), .D(n_1708), .Y(n_1665) );
NAND3xp33_ASAP7_75t_L g1674 ( .A(n_1669), .B(n_1675), .C(n_1676), .Y(n_1674) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1673), .Y(n_1686) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
O2A1O1Ixp33_ASAP7_75t_L g1681 ( .A1(n_1682), .A2(n_1686), .B(n_1687), .C(n_1689), .Y(n_1681) );
INVxp67_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1693), .Y(n_1706) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1694), .Y(n_1716) );
CKINVDCx14_ASAP7_75t_R g1695 ( .A(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVxp67_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1707), .Y(n_1705) );
NAND4xp25_ASAP7_75t_L g1713 ( .A(n_1714), .B(n_1724), .C(n_1733), .D(n_1736), .Y(n_1713) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
NAND2xp5_ASAP7_75t_SL g1725 ( .A(n_1726), .B(n_1727), .Y(n_1725) );
INVxp67_ASAP7_75t_SL g1728 ( .A(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
CKINVDCx20_ASAP7_75t_R g1739 ( .A(n_1740), .Y(n_1739) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx2_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
AND3x2_ASAP7_75t_L g1745 ( .A(n_1746), .B(n_1783), .C(n_1799), .Y(n_1745) );
AOI211xp5_ASAP7_75t_SL g1746 ( .A1(n_1747), .A2(n_1748), .B(n_1754), .C(n_1767), .Y(n_1746) );
INVxp67_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx2_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1752), .Y(n_1782) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
AND2x4_ASAP7_75t_L g1762 ( .A(n_1757), .B(n_1763), .Y(n_1762) );
AND2x4_ASAP7_75t_L g1757 ( .A(n_1758), .B(n_1759), .Y(n_1757) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1758), .B(n_1788), .Y(n_1787) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
INVx2_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
INVx3_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
OAI221xp5_ASAP7_75t_L g1806 ( .A1(n_1772), .A2(n_1778), .B1(n_1807), .B2(n_1809), .C(n_1811), .Y(n_1806) );
INVxp67_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
AOI21xp5_ASAP7_75t_L g1783 ( .A1(n_1784), .A2(n_1790), .B(n_1791), .Y(n_1783) );
INVx8_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
AND2x4_ASAP7_75t_L g1785 ( .A(n_1786), .B(n_1787), .Y(n_1785) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1789), .Y(n_1824) );
AND2x4_ASAP7_75t_L g1792 ( .A(n_1793), .B(n_1795), .Y(n_1792) );
OR2x6_ASAP7_75t_L g1796 ( .A(n_1797), .B(n_1798), .Y(n_1796) );
OAI31xp33_ASAP7_75t_L g1799 ( .A1(n_1800), .A2(n_1817), .A3(n_1829), .B(n_1835), .Y(n_1799) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
INVx4_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
INVx2_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
INVx2_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
INVx2_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
INVxp67_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
HB1xp67_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
INVx2_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
NOR2x1_ASAP7_75t_L g1822 ( .A(n_1823), .B(n_1824), .Y(n_1822) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
BUFx6f_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
INVx3_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx2_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
BUFx3_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
BUFx2_ASAP7_75t_SL g1842 ( .A(n_1843), .Y(n_1842) );
BUFx3_ASAP7_75t_L g1843 ( .A(n_1844), .Y(n_1843) );
INVxp33_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
HB1xp67_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
INVx1_ASAP7_75t_L g1849 ( .A(n_1850), .Y(n_1849) );
NAND3xp33_ASAP7_75t_L g1850 ( .A(n_1851), .B(n_1861), .C(n_1868), .Y(n_1850) );
INVx2_ASAP7_75t_SL g1854 ( .A(n_1855), .Y(n_1854) );
NOR2xp33_ASAP7_75t_L g1868 ( .A(n_1869), .B(n_1883), .Y(n_1868) );
OAI22xp33_ASAP7_75t_L g1884 ( .A1(n_1871), .A2(n_1878), .B1(n_1885), .B2(n_1887), .Y(n_1884) );
INVx2_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
INVx2_ASAP7_75t_SL g1891 ( .A(n_1892), .Y(n_1891) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1893), .Y(n_1892) );
OAI21xp5_ASAP7_75t_L g1893 ( .A1(n_1894), .A2(n_1895), .B(n_1896), .Y(n_1893) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
endmodule