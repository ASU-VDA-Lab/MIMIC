module fake_jpeg_2473_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_81),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_67),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_69),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_66),
.B1(n_55),
.B2(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_59),
.B1(n_55),
.B2(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_94),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_53),
.B1(n_71),
.B2(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_101),
.Y(n_126)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_51),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_82),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_94),
.B1(n_66),
.B2(n_54),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_116),
.B1(n_125),
.B2(n_65),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_88),
.B1(n_66),
.B2(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_64),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_97),
.B1(n_111),
.B2(n_107),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_70),
.B(n_56),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_11),
.B(n_12),
.Y(n_156)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_68),
.B(n_60),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_60),
.C(n_73),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_124),
.C(n_128),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_73),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_54),
.B1(n_65),
.B2(n_80),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_3),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_4),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_27),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_139),
.Y(n_171)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_140),
.B1(n_13),
.B2(n_14),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_64),
.C(n_23),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_22),
.C(n_48),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_21),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_5),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_11),
.B(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_8),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_10),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_155),
.A2(n_156),
.B(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_159),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_115),
.B(n_31),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_164),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_32),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_166),
.B1(n_15),
.B2(n_16),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_28),
.B(n_45),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_144),
.C(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_175),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_136),
.B1(n_148),
.B2(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_137),
.B(n_145),
.C(n_15),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_160),
.B(n_168),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_13),
.C(n_14),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_180),
.B(n_170),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_159),
.B(n_167),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_178),
.B(n_177),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_184),
.B(n_174),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_187),
.B(n_189),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_161),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_190),
.A3(n_186),
.B1(n_185),
.B2(n_161),
.C1(n_34),
.C2(n_35),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_39),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_37),
.Y(n_195)
);

AOI31xp33_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_41),
.A3(n_19),
.B(n_20),
.Y(n_196)
);

OAI321xp33_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_24),
.A3(n_43),
.B1(n_50),
.B2(n_192),
.C(n_17),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_17),
.Y(n_198)
);


endmodule