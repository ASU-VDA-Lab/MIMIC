module fake_netlist_1_10204_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
AND3x2_ASAP7_75t_L g4 ( .A(n_0), .B(n_2), .C(n_1), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
AND2x2_ASAP7_75t_SL g7 ( .A(n_5), .B(n_4), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AOI221xp5_ASAP7_75t_SL g9 ( .A1(n_8), .A2(n_6), .B1(n_5), .B2(n_0), .C(n_1), .Y(n_9) );
A2O1A1Ixp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_2), .B(n_7), .C(n_8), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_10), .B(n_9), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_11), .B(n_2), .Y(n_12) );
endmodule