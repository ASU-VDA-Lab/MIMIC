module fake_jpeg_11430_n_641 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_641);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_641;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_576;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_0),
.B(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_73),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_11),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_63),
.B(n_117),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_27),
.B(n_9),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_30),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_75),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_9),
.C(n_16),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_85),
.A2(n_58),
.B(n_42),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_86),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_88),
.Y(n_148)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

AND2x4_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_9),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_43),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_21),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_91),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_101),
.Y(n_206)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_23),
.B(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_120),
.Y(n_141)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_20),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_118),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_109),
.Y(n_154)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_111),
.Y(n_204)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_23),
.B(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_26),
.B(n_13),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_26),
.B(n_13),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_34),
.B(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_18),
.Y(n_163)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_19),
.Y(n_125)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_36),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_135),
.B(n_140),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_43),
.B1(n_55),
.B2(n_20),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_137),
.A2(n_200),
.B1(n_57),
.B2(n_48),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_36),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_163),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_54),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_150),
.B(n_157),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_54),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_166),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_90),
.B(n_58),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_56),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_69),
.A2(n_43),
.B1(n_56),
.B2(n_50),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_172),
.A2(n_64),
.B1(n_94),
.B2(n_92),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_77),
.B(n_50),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_42),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_52),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_194),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_109),
.B(n_52),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_60),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_84),
.A2(n_89),
.B1(n_105),
.B2(n_108),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_193),
.B1(n_83),
.B2(n_79),
.Y(n_247)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_65),
.A2(n_24),
.B1(n_59),
.B2(n_46),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_96),
.B(n_39),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_66),
.B(n_59),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_76),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_67),
.A2(n_20),
.B1(n_60),
.B2(n_46),
.Y(n_200)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_209),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_24),
.B(n_116),
.C(n_74),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_210),
.B(n_237),
.Y(n_309)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_211),
.Y(n_322)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_128),
.Y(n_213)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_213),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_217),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_137),
.A2(n_86),
.B1(n_101),
.B2(n_100),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_218),
.A2(n_247),
.B1(n_266),
.B2(n_283),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_220),
.B(n_245),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_224),
.B(n_281),
.Y(n_291)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_230),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_231),
.A2(n_274),
.B1(n_148),
.B2(n_190),
.Y(n_290)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_232),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_233),
.B(n_250),
.Y(n_285)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_143),
.Y(n_235)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g237 ( 
.A1(n_159),
.A2(n_82),
.B1(n_88),
.B2(n_87),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_133),
.B(n_125),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_239),
.B(n_253),
.Y(n_345)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_240),
.Y(n_299)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_241),
.Y(n_328)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_243),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_201),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_134),
.Y(n_248)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

INVx3_ASAP7_75t_SL g249 ( 
.A(n_136),
.Y(n_249)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

INVx4_ASAP7_75t_SL g253 ( 
.A(n_204),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_152),
.Y(n_254)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_254),
.Y(n_339)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_256),
.Y(n_341)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_257),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_198),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_259),
.Y(n_316)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_134),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_260),
.A2(n_262),
.B1(n_272),
.B2(n_278),
.Y(n_327)
);

BUFx2_ASAP7_75t_SL g261 ( 
.A(n_154),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_261),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_271),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_132),
.B(n_141),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_267),
.B(n_269),
.Y(n_293)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_265),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_149),
.A2(n_68),
.B1(n_60),
.B2(n_57),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_138),
.B(n_60),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_268),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_130),
.B(n_60),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_270),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_154),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_146),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_273),
.B(n_275),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_202),
.A2(n_57),
.B1(n_48),
.B2(n_25),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_160),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_146),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_176),
.B(n_15),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_204),
.C(n_148),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_136),
.Y(n_278)
);

BUFx8_ASAP7_75t_L g279 ( 
.A(n_127),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_127),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_176),
.B(n_15),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_179),
.B(n_15),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_282),
.B(n_6),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_200),
.A2(n_57),
.B1(n_48),
.B2(n_25),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_250),
.A2(n_231),
.B1(n_228),
.B2(n_272),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_284),
.A2(n_331),
.B1(n_269),
.B2(n_278),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_279),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_279),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_218),
.A2(n_177),
.B1(n_196),
.B2(n_147),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_298),
.A2(n_313),
.B1(n_320),
.B2(n_335),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_221),
.A2(n_180),
.B1(n_179),
.B2(n_182),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_312),
.A2(n_216),
.B(n_222),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_221),
.A2(n_267),
.B1(n_239),
.B2(n_237),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_314),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_210),
.A2(n_206),
.B1(n_192),
.B2(n_164),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_317),
.A2(n_227),
.B1(n_213),
.B2(n_254),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_239),
.A2(n_237),
.B1(n_214),
.B2(n_215),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_277),
.A2(n_25),
.B(n_48),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_323),
.A2(n_238),
.B(n_268),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_329),
.Y(n_346)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_212),
.B(n_177),
.CI(n_192),
.CON(n_329),
.SN(n_329)
);

OAI22x1_ASAP7_75t_SL g331 ( 
.A1(n_274),
.A2(n_182),
.B1(n_206),
.B2(n_164),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_264),
.B(n_16),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_333),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_280),
.B(n_16),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_239),
.A2(n_196),
.B1(n_169),
.B2(n_147),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_219),
.B(n_160),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_249),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_347),
.A2(n_349),
.B1(n_359),
.B2(n_367),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_284),
.A2(n_169),
.B1(n_151),
.B2(n_158),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_380),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_352),
.A2(n_363),
.B(n_365),
.Y(n_434)
);

O2A1O1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_309),
.A2(n_253),
.B(n_229),
.C(n_270),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_354),
.A2(n_355),
.B(n_373),
.Y(n_399)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_234),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_240),
.C(n_211),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_287),
.C(n_304),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_357),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_361),
.B1(n_369),
.B2(n_375),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_296),
.A2(n_144),
.B1(n_265),
.B2(n_158),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_360),
.B(n_323),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_296),
.A2(n_144),
.B1(n_248),
.B2(n_230),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_345),
.A2(n_244),
.B1(n_260),
.B2(n_262),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_316),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_377),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_331),
.A2(n_241),
.B1(n_223),
.B2(n_217),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_320),
.A2(n_25),
.B1(n_19),
.B2(n_1),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_19),
.B(n_3),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_370),
.A2(n_387),
.B(n_325),
.Y(n_421)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_303),
.A2(n_2),
.B(n_18),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_379),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_313),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_298),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_376),
.A2(n_391),
.B1(n_375),
.B2(n_358),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_344),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_308),
.A2(n_6),
.B1(n_14),
.B2(n_16),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_378),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_291),
.B(n_14),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_14),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_18),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_390),
.Y(n_424)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_18),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_383),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_335),
.B(n_293),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g419 ( 
.A(n_384),
.B(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_285),
.A2(n_312),
.B(n_329),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_337),
.B(n_326),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_327),
.A2(n_307),
.B1(n_306),
.B2(n_326),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_297),
.B(n_341),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_302),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_307),
.A2(n_311),
.B1(n_328),
.B2(n_337),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_393),
.A2(n_305),
.B1(n_328),
.B2(n_325),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_398),
.B(n_411),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_402),
.B(n_405),
.C(n_407),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_341),
.C(n_287),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_286),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_359),
.A2(n_306),
.B1(n_334),
.B2(n_318),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_408),
.A2(n_430),
.B1(n_433),
.B2(n_386),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_292),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_415),
.A2(n_363),
.B1(n_365),
.B2(n_380),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_356),
.B(n_292),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_417),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_302),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_418),
.A2(n_358),
.B1(n_391),
.B2(n_361),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_419),
.A2(n_421),
.B(n_352),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_366),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_422),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_353),
.A2(n_318),
.B1(n_334),
.B2(n_315),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_425),
.A2(n_367),
.B1(n_363),
.B2(n_365),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_304),
.C(n_338),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_390),
.Y(n_445)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_429),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_347),
.A2(n_338),
.B1(n_340),
.B2(n_321),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_371),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_339),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_373),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_349),
.A2(n_321),
.B1(n_340),
.B2(n_300),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_435),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_394),
.A2(n_355),
.B(n_346),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_436),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_410),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_440),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_431),
.Y(n_440)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_428),
.Y(n_443)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_444),
.B(n_448),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_445),
.B(n_470),
.C(n_472),
.Y(n_488)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_423),
.Y(n_447)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_350),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_449),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_434),
.A2(n_355),
.B(n_348),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_454),
.Y(n_485)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_400),
.Y(n_451)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_396),
.B(n_392),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_388),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_406),
.B(n_388),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_465),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_460),
.B1(n_469),
.B2(n_399),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_357),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_471),
.B1(n_404),
.B2(n_425),
.Y(n_482)
);

OAI22x1_ASAP7_75t_SL g460 ( 
.A1(n_415),
.A2(n_354),
.B1(n_393),
.B2(n_381),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_394),
.A2(n_346),
.B(n_384),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_463),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_421),
.A2(n_354),
.B(n_384),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_464),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_406),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_466),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_395),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_440),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_353),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_413),
.A2(n_358),
.B1(n_369),
.B2(n_376),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_407),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_475),
.B(n_501),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_469),
.A2(n_409),
.B1(n_426),
.B2(n_430),
.Y(n_477)
);

XOR2x1_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_455),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_492),
.B1(n_496),
.B2(n_460),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_484),
.A2(n_450),
.B1(n_463),
.B2(n_436),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_454),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_500),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_499),
.C(n_503),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_471),
.A2(n_404),
.B1(n_409),
.B2(n_399),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_442),
.B(n_417),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_494),
.B(n_448),
.Y(n_521)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_459),
.A2(n_424),
.B1(n_405),
.B2(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_435),
.Y(n_497)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_442),
.B(n_416),
.C(n_398),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_453),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_438),
.B(n_424),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_457),
.B(n_429),
.Y(n_502)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_438),
.B(n_397),
.C(n_401),
.Y(n_503)
);

OA21x2_ASAP7_75t_SL g506 ( 
.A1(n_462),
.A2(n_397),
.B(n_434),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_506),
.A2(n_458),
.B(n_383),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_508),
.A2(n_477),
.B1(n_505),
.B2(n_487),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g509 ( 
.A(n_485),
.B(n_439),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_514),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_SL g510 ( 
.A(n_496),
.B(n_445),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_SL g553 ( 
.A(n_510),
.B(n_513),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_511),
.A2(n_524),
.B1(n_492),
.B2(n_505),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_470),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_535),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_495),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_499),
.C(n_494),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_517),
.B(n_518),
.C(n_525),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_501),
.C(n_483),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_521),
.B(n_526),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g522 ( 
.A(n_480),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_523),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_484),
.A2(n_467),
.B1(n_437),
.B2(n_452),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_483),
.B(n_468),
.C(n_466),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_474),
.B(n_444),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_527),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_383),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_529),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_485),
.B(n_383),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_497),
.Y(n_530)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_530),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_532),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_489),
.A2(n_491),
.B(n_493),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_490),
.B(n_351),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_370),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_464),
.C(n_441),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_502),
.C(n_478),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_478),
.B(n_461),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_SL g564 ( 
.A(n_541),
.B(n_559),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_558),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_480),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_547),
.B(n_549),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_479),
.B1(n_476),
.B2(n_408),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_512),
.B(n_482),
.C(n_490),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_473),
.C(n_504),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_554),
.C(n_555),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_523),
.B(n_351),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_551),
.B(n_560),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_504),
.Y(n_552)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_552),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_519),
.B(n_473),
.C(n_498),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_507),
.B(n_518),
.C(n_517),
.Y(n_555)
);

FAx1_ASAP7_75t_L g557 ( 
.A(n_511),
.B(n_524),
.CI(n_513),
.CON(n_557),
.SN(n_557)
);

AOI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_557),
.A2(n_456),
.B1(n_528),
.B2(n_476),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_507),
.B(n_498),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_486),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_486),
.Y(n_561)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_561),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_556),
.A2(n_525),
.B(n_536),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_565),
.B(n_568),
.C(n_570),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_508),
.C(n_535),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_573),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_481),
.Y(n_568)
);

MAJx2_ASAP7_75t_L g569 ( 
.A(n_549),
.B(n_509),
.C(n_515),
.Y(n_569)
);

XOR2x2_ASAP7_75t_SL g585 ( 
.A(n_569),
.B(n_575),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_550),
.B(n_481),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_509),
.C(n_516),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_538),
.B(n_529),
.C(n_520),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_576),
.Y(n_588)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_545),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_579),
.Y(n_596)
);

BUFx24_ASAP7_75t_SL g578 ( 
.A(n_544),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_578),
.B(n_538),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_537),
.B(n_479),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_546),
.A2(n_449),
.B1(n_447),
.B2(n_446),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_580),
.B(n_581),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_537),
.B(n_446),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_584),
.B(n_590),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_566),
.B(n_555),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_587),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_539),
.C(n_540),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_575),
.A2(n_557),
.B(n_553),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_591),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_562),
.B(n_368),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_573),
.A2(n_557),
.B(n_564),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_571),
.A2(n_539),
.B1(n_542),
.B2(n_558),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_597),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_451),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_594),
.A2(n_598),
.B(n_599),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_582),
.A2(n_542),
.B(n_441),
.Y(n_597)
);

AOI21x1_ASAP7_75t_SL g609 ( 
.A1(n_597),
.A2(n_412),
.B(n_401),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_574),
.B(n_428),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_567),
.B(n_389),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_389),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_600),
.A2(n_382),
.B(n_339),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_569),
.C(n_581),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_601),
.B(n_604),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_SL g604 ( 
.A(n_593),
.B(n_572),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_572),
.C(n_443),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_611),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_400),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_607),
.B(n_589),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_609),
.A2(n_614),
.B(n_378),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_414),
.C(n_412),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_585),
.C(n_289),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_596),
.B(n_414),
.C(n_385),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_612),
.B(n_613),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g614 ( 
.A(n_585),
.B(n_322),
.Y(n_614)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_603),
.A2(n_595),
.B(n_592),
.Y(n_617)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_617),
.Y(n_626)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_618),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_619),
.B(n_611),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_620),
.B(n_622),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_289),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_621),
.A2(n_608),
.B(n_300),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_605),
.B(n_288),
.Y(n_622)
);

OA21x2_ASAP7_75t_L g623 ( 
.A1(n_602),
.A2(n_609),
.B(n_612),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_623),
.B(n_602),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_625),
.A2(n_629),
.B(n_294),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_627),
.B(n_628),
.C(n_624),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_604),
.Y(n_629)
);

A2O1A1O1Ixp25_ASAP7_75t_L g632 ( 
.A1(n_625),
.A2(n_623),
.B(n_618),
.C(n_624),
.D(n_615),
.Y(n_632)
);

AOI31xp33_ASAP7_75t_L g636 ( 
.A1(n_632),
.A2(n_633),
.A3(n_634),
.B(n_626),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_631),
.B(n_288),
.C(n_301),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_635),
.A2(n_630),
.B(n_301),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_636),
.B(n_637),
.C(n_294),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_319),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_319),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_640),
.B(n_342),
.C(n_603),
.Y(n_641)
);


endmodule