module fake_jpeg_19533_n_272 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_41),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_52),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_21),
.B1(n_13),
.B2(n_29),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_41),
.B(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_21),
.B1(n_13),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_37),
.B1(n_40),
.B2(n_26),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_33),
.B(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_46),
.B1(n_44),
.B2(n_52),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_24),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_57),
.C(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_38),
.Y(n_63)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_68),
.B1(n_55),
.B2(n_57),
.Y(n_80)
);

OA21x2_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_41),
.B(n_42),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_51),
.B1(n_58),
.B2(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_35),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_77),
.B1(n_47),
.B2(n_50),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_74),
.B1(n_55),
.B2(n_48),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_37),
.B1(n_40),
.B2(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_92),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_82),
.B(n_87),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_51),
.B(n_54),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_22),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_75),
.B(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_56),
.B1(n_47),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_56),
.B1(n_55),
.B2(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_28),
.B1(n_41),
.B2(n_49),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_94),
.B1(n_68),
.B2(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_39),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_61),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_41),
.B1(n_30),
.B2(n_25),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_45),
.C(n_49),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_62),
.C(n_72),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_105),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_76),
.B1(n_65),
.B2(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_102),
.B1(n_117),
.B2(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_107),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_82),
.C(n_95),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_110),
.C(n_113),
.Y(n_118)
);

XNOR2x2_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_92),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_106),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_81),
.B(n_89),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_16),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_67),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_65),
.B1(n_27),
.B2(n_34),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_128),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_129),
.B1(n_14),
.B2(n_7),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_84),
.B1(n_91),
.B2(n_81),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_130),
.B1(n_139),
.B2(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_148)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_86),
.B(n_10),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_132),
.B(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_12),
.B1(n_23),
.B2(n_22),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_35),
.B1(n_59),
.B2(n_11),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_138),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_23),
.B(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_35),
.B1(n_59),
.B2(n_23),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_0),
.B1(n_1),
.B2(n_17),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_18),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_8),
.B(n_10),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_106),
.C(n_18),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_149),
.C(n_158),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_163),
.B1(n_141),
.B2(n_128),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_18),
.C(n_14),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_166),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_16),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_153),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_16),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_16),
.B1(n_19),
.B2(n_15),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_16),
.B(n_18),
.C(n_14),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_130),
.B(n_120),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_18),
.C(n_14),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_129),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_135),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_168),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_14),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_122),
.B(n_145),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_173),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_147),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_185),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_144),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_126),
.B1(n_127),
.B2(n_139),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_137),
.C(n_142),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_190),
.C(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_119),
.C(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_156),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_161),
.B1(n_191),
.B2(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_199),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_159),
.B1(n_146),
.B2(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_202),
.B1(n_201),
.B2(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_167),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_154),
.B(n_132),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_202),
.B(n_7),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_154),
.B(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_156),
.B1(n_158),
.B2(n_153),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_209),
.B1(n_184),
.B2(n_185),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_179),
.C(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_156),
.B1(n_17),
.B2(n_19),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_212),
.B1(n_6),
.B2(n_3),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_182),
.B1(n_181),
.B2(n_183),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_217),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_207),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_194),
.C(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_19),
.C(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_225),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_209),
.B(n_204),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_7),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_8),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_6),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_228),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_217),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_223),
.B(n_218),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_196),
.B(n_3),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_19),
.C(n_4),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_212),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_243),
.B(n_241),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_214),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_211),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_5),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_224),
.C(n_247),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_231),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_SL g260 ( 
.A(n_251),
.B(n_255),
.C(n_253),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_5),
.C(n_6),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_263),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_260),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_261),
.A2(n_256),
.B(n_9),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_8),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_259),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_268),
.B(n_265),
.C(n_9),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_262),
.C(n_9),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_9),
.C(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_270),
.B(n_0),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_10),
.Y(n_272)
);


endmodule