module real_jpeg_18435_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_0),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_0),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_0),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_0),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_0),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_0),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_1),
.Y(n_161)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_3),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_3),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_4),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_4),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_4),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_4),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_4),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_4),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_4),
.B(n_410),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_78),
.Y(n_77)
);

NAND2xp67_ASAP7_75t_SL g79 ( 
.A(n_6),
.B(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_9),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

NAND2x1_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_6),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_7),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_8),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_8),
.B(n_147),
.Y(n_146)
);

AND2x4_ASAP7_75t_SL g244 ( 
.A(n_8),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_8),
.B(n_255),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_8),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_8),
.B(n_143),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_9),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_9),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_9),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_9),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_9),
.B(n_143),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_9),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_9),
.B(n_385),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_11),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_11),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_11),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_11),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_11),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_11),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_11),
.B(n_294),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_12),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_12),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_14),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_15),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_15),
.B(n_35),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_15),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_15),
.B(n_255),
.Y(n_254)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_16),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_223),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_222),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_181),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_21),
.B(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.C(n_155),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_23),
.B(n_155),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_69),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_24),
.B(n_70),
.C(n_88),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.C(n_55),
.Y(n_24)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_25),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_28),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_33),
.Y(n_305)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_38),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_39),
.B(n_55),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_50),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_40),
.A2(n_50),
.B1(n_51),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_40),
.Y(n_265)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_46),
.B(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_49),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_50),
.B(n_323),
.C(n_327),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_50),
.A2(n_51),
.B1(n_323),
.B2(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_56),
.B(n_61),
.C(n_65),
.Y(n_169)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_61),
.A2(n_160),
.B1(n_166),
.B2(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_61),
.B(n_117),
.C(n_160),
.Y(n_217)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_62),
.Y(n_386)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_63),
.Y(n_365)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_88),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_79),
.C(n_83),
.Y(n_70)
);

XNOR2x1_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.C(n_77),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_77),
.Y(n_107)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_78),
.Y(n_252)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_78),
.Y(n_300)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_78),
.Y(n_363)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_78),
.Y(n_411)
);

AOI22x1_ASAP7_75t_SL g153 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_83),
.A2(n_84),
.B1(n_302),
.B2(n_303),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_84),
.B(n_297),
.C(n_302),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_87),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_89),
.B(n_91),
.C(n_98),
.Y(n_220)
);

OAI22x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_92),
.B(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_96),
.Y(n_326)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_103),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_128),
.C(n_151),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_105),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_115),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_106),
.B(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_108),
.A2(n_109),
.B1(n_115),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21x1_ASAP7_75t_SL g283 ( 
.A1(n_109),
.A2(n_284),
.B(n_291),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_110),
.Y(n_255)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_115),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_125),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_117),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_116),
.A2(n_117),
.B1(n_125),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_121),
.B(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_128),
.A2(n_151),
.B1(n_152),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_141),
.C(n_146),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_129),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_137),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_130),
.A2(n_137),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_130),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_130),
.B(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_134),
.B(n_280),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_161),
.Y(n_194)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_168),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_157),
.B(n_169),
.C(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_160),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_167),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_164),
.Y(n_358)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_175),
.C(n_197),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_212),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_220),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_217),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_266),
.B(n_440),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_225),
.B(n_227),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

XOR2x2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_260),
.C(n_263),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_248),
.C(n_256),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_239),
.B(n_249),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_244),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_240),
.A2(n_242),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_240),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_242),
.A2(n_320),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_242),
.B(n_388),
.C(n_392),
.Y(n_418)
);

XOR2x1_ASAP7_75t_SL g317 ( 
.A(n_244),
.B(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_250),
.B(n_254),
.Y(n_334)
);

NOR2x1_ASAP7_75t_R g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_257),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_337),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.C(n_309),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_271),
.B(n_275),
.Y(n_338)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.C(n_306),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_283),
.C(n_296),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_281),
.B(n_348),
.C(n_353),
.Y(n_375)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_297),
.B(n_427),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_298),
.B(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_298),
.A2(n_383),
.B1(n_384),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_312),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_335),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_313),
.B(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_316),
.B(n_335),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.C(n_333),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_317),
.B(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_322),
.B(n_334),
.Y(n_432)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2x2_ASAP7_75t_SL g376 ( 
.A(n_327),
.B(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_435),
.B(n_439),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_421),
.B(n_434),
.Y(n_341)
);

OAI21x1_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_379),
.B(n_420),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_368),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_368),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_354),
.C(n_360),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_346),
.B(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_354),
.A2(n_355),
.B1(n_360),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_356),
.B(n_359),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

AO22x1_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_364),
.B1(n_366),
.B2(n_367),
.Y(n_360)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_364),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_366),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_R g408 ( 
.A(n_367),
.B(n_409),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_374),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_369),
.B(n_375),
.C(n_376),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_372),
.C(n_373),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_414),
.B(n_419),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_396),
.B(n_413),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_387),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_408),
.B(n_412),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_406),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_406),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_SL g419 ( 
.A(n_415),
.B(n_418),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_433),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_SL g434 ( 
.A(n_422),
.B(n_433),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_430),
.B2(n_431),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_429),
.C(n_430),
.Y(n_436)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_436),
.B(n_437),
.Y(n_439)
);


endmodule