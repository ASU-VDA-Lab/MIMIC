module fake_aes_4208_n_557 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_557);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_557;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_47), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_12), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_43), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_18), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_38), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_32), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_57), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_29), .Y(n_87) );
NOR2xp33_ASAP7_75t_L g88 ( .A(n_54), .B(n_26), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_51), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_42), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_30), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_40), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_74), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_14), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_11), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_5), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_62), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_44), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_70), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_50), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_28), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_16), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_63), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_5), .B(n_22), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_10), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_55), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_76), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_65), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_102), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_99), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_80), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_102), .B(n_0), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_99), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_110), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_98), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_81), .B(n_3), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_85), .B(n_4), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_84), .B(n_6), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_108), .B(n_6), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
NOR2xp33_ASAP7_75t_R g132 ( .A(n_91), .B(n_45), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_79), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_95), .B(n_7), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_93), .B(n_7), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_113), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_79), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_135), .A2(n_129), .B1(n_130), .B2(n_119), .Y(n_139) );
NOR2x1p5_ASAP7_75t_L g140 ( .A(n_129), .B(n_112), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_115), .B(n_97), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_116), .B(n_105), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_135), .A2(n_96), .B1(n_93), .B2(n_112), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
INVxp67_ASAP7_75t_SL g148 ( .A(n_117), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_131), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_123), .B(n_101), .Y(n_150) );
INVx5_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
AND3x1_ASAP7_75t_L g153 ( .A(n_135), .B(n_86), .C(n_104), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_133), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_116), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_117), .B(n_94), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g158 ( .A(n_122), .B(n_94), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_122), .B(n_107), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_123), .B(n_103), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_129), .B(n_114), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_158), .B(n_132), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_153), .A2(n_130), .B1(n_120), .B2(n_124), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_159), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_154), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_148), .B(n_125), .Y(n_174) );
NOR2x2_ASAP7_75t_L g175 ( .A(n_154), .B(n_126), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_165), .B(n_130), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_139), .B(n_119), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_153), .A2(n_124), .B1(n_134), .B2(n_126), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_165), .B(n_138), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_150), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_158), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
BUFx12f_ASAP7_75t_L g187 ( .A(n_140), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_164), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_140), .A2(n_127), .B1(n_131), .B2(n_138), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_144), .A2(n_127), .B(n_138), .C(n_128), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_155), .B(n_104), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_155), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_189), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_193), .A2(n_157), .B(n_145), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_178), .B(n_139), .Y(n_204) );
BUFx2_ASAP7_75t_SL g205 ( .A(n_184), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_176), .A2(n_162), .B(n_144), .C(n_163), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_184), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
AOI22xp33_ASAP7_75t_SL g210 ( .A1(n_183), .A2(n_163), .B1(n_150), .B2(n_143), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_184), .B(n_150), .Y(n_211) );
AOI21x1_ASAP7_75t_L g212 ( .A1(n_197), .A2(n_163), .B(n_162), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
INVx8_ASAP7_75t_L g214 ( .A(n_187), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_184), .B(n_163), .Y(n_215) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_183), .B(n_190), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_191), .B(n_146), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_182), .B(n_143), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_187), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_189), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_168), .A2(n_146), .B1(n_143), .B2(n_145), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_142), .B(n_145), .C(n_118), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_171), .Y(n_224) );
NOR2xp33_ASAP7_75t_R g225 ( .A(n_178), .B(n_8), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_193), .A2(n_199), .B(n_169), .Y(n_226) );
NOR2xp33_ASAP7_75t_R g227 ( .A(n_182), .B(n_185), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_170), .B(n_151), .Y(n_229) );
INVx1_ASAP7_75t_SL g230 ( .A(n_186), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_194), .A2(n_136), .B1(n_121), .B2(n_118), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_168), .A2(n_179), .B1(n_167), .B2(n_180), .Y(n_233) );
INVx6_ASAP7_75t_L g234 ( .A(n_185), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_213), .A2(n_179), .B1(n_180), .B2(n_173), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_207), .A2(n_196), .B(n_192), .C(n_188), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_204), .B(n_185), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_223), .A2(n_192), .B(n_188), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_223), .A2(n_160), .B(n_152), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g243 ( .A1(n_224), .A2(n_175), .B1(n_219), .B2(n_210), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_215), .B(n_166), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_208), .B(n_173), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_217), .B(n_166), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_230), .A2(n_169), .B1(n_177), .B2(n_198), .Y(n_248) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_221), .A2(n_160), .B(n_152), .Y(n_249) );
BUFx2_ASAP7_75t_R g250 ( .A(n_205), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_212), .A2(n_200), .B(n_195), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_201), .A2(n_177), .B(n_109), .C(n_118), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g258 ( .A1(n_225), .A2(n_118), .B1(n_121), .B2(n_87), .Y(n_258) );
OR2x6_ASAP7_75t_L g259 ( .A(n_215), .B(n_121), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_198), .B(n_200), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_203), .Y(n_261) );
NOR2x1_ASAP7_75t_R g262 ( .A(n_214), .B(n_106), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_251), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_254), .B(n_220), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_250), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_241), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_241), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_238), .B(n_220), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_121), .B1(n_216), .B2(n_231), .C(n_211), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_256), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_251), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_251), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_236), .A2(n_202), .B(n_211), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
INVx4_ASAP7_75t_L g275 ( .A(n_251), .Y(n_275) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_249), .A2(n_152), .B(n_160), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_261), .B(n_222), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_261), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_246), .B(n_222), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_246), .A2(n_218), .B1(n_228), .B2(n_234), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_239), .B(n_222), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_235), .B(n_228), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_259), .B(n_218), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_253), .A2(n_218), .B1(n_234), .B2(n_227), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_271), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_269), .A2(n_258), .B1(n_257), .B2(n_259), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_270), .B(n_247), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_270), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_274), .B(n_240), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_274), .B(n_255), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_266), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_266), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_278), .B(n_255), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_278), .B(n_259), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_267), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_283), .B(n_257), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_279), .B(n_259), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_269), .A2(n_244), .B1(n_249), .B2(n_251), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_264), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_271), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_275), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_288), .B(n_279), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_306), .B(n_262), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_298), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_308), .B(n_281), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_308), .B(n_281), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_290), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_298), .B(n_276), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_293), .B(n_280), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_290), .B(n_276), .Y(n_317) );
OAI33xp33_ASAP7_75t_L g318 ( .A1(n_299), .A2(n_89), .A3(n_90), .B1(n_92), .B2(n_100), .B3(n_101), .Y(n_318) );
OAI211xp5_ASAP7_75t_SL g319 ( .A1(n_287), .A2(n_285), .B(n_89), .C(n_90), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_288), .B(n_268), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_293), .B(n_276), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_307), .B(n_275), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_300), .A2(n_280), .B1(n_268), .B2(n_284), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_295), .B(n_282), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_284), .B1(n_273), .B2(n_282), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_307), .B(n_275), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_305), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_296), .B(n_242), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g332 ( .A1(n_301), .A2(n_273), .B1(n_284), .B2(n_265), .C(n_236), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_296), .B(n_289), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_289), .B(n_242), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g335 ( .A1(n_301), .A2(n_284), .B1(n_92), .B2(n_103), .C(n_100), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_294), .B(n_242), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_307), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_297), .A2(n_284), .B1(n_244), .B2(n_277), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_333), .B(n_305), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
NAND2xp67_ASAP7_75t_L g342 ( .A(n_321), .B(n_292), .Y(n_342) );
NOR3xp33_ASAP7_75t_L g343 ( .A(n_310), .B(n_111), .C(n_292), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_333), .B(n_294), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_330), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_314), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
NAND4xp25_ASAP7_75t_L g349 ( .A(n_332), .B(n_302), .C(n_113), .D(n_114), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_320), .B(n_303), .Y(n_350) );
NAND4xp75_ASAP7_75t_L g351 ( .A(n_337), .B(n_291), .C(n_303), .D(n_263), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_327), .B(n_291), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_327), .B(n_275), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_313), .B(n_304), .Y(n_354) );
NAND4xp25_ASAP7_75t_L g355 ( .A(n_323), .B(n_88), .C(n_244), .D(n_277), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_313), .B(n_304), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_311), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_313), .B(n_304), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_339), .Y(n_360) );
AND3x1_ASAP7_75t_L g361 ( .A(n_323), .B(n_8), .C(n_9), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_324), .B(n_304), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_330), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_313), .B(n_304), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_328), .Y(n_369) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_322), .B(n_284), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_312), .B(n_304), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_312), .B(n_286), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_309), .B(n_286), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_322), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_335), .A2(n_245), .B(n_277), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_321), .B(n_286), .Y(n_378) );
NAND2xp33_ASAP7_75t_R g379 ( .A(n_326), .B(n_10), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_329), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_337), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_326), .B(n_286), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_316), .B(n_286), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_315), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_331), .B(n_286), .Y(n_385) );
AND2x4_ASAP7_75t_SL g386 ( .A(n_348), .B(n_326), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_368), .B(n_331), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_350), .B(n_317), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_385), .B(n_317), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_352), .B(n_316), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_341), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_384), .B(n_315), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_385), .B(n_336), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_361), .B(n_326), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_384), .B(n_325), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_357), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_372), .B(n_336), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_372), .B(n_334), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_373), .B(n_334), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_341), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_373), .B(n_338), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_355), .B(n_318), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_344), .B(n_263), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_346), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_344), .B(n_263), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_360), .B(n_363), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_340), .B(n_11), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_354), .B(n_272), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_358), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_354), .B(n_272), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_340), .B(n_12), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_362), .B(n_13), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_357), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_364), .Y(n_417) );
NOR2xp67_ASAP7_75t_L g418 ( .A(n_348), .B(n_13), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_362), .B(n_14), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_375), .B(n_15), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_342), .B(n_15), .Y(n_421) );
NOR2xp33_ASAP7_75t_SL g422 ( .A(n_351), .B(n_214), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_370), .Y(n_423) );
OAI21xp33_ASAP7_75t_SL g424 ( .A1(n_351), .A2(n_252), .B(n_319), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_345), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_342), .B(n_272), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_348), .B(n_271), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_376), .B(n_252), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_376), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_366), .B(n_245), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_358), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_365), .B(n_156), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_378), .B(n_245), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_376), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_356), .B(n_19), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_353), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_369), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_383), .B(n_156), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_404), .A2(n_343), .B1(n_349), .B2(n_381), .C(n_380), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_390), .B(n_356), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_401), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_388), .Y(n_444) );
OAI32xp33_ASAP7_75t_L g445 ( .A1(n_424), .A2(n_379), .A3(n_383), .B1(n_377), .B2(n_380), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g447 ( .A(n_423), .B(n_370), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_395), .A2(n_374), .B1(n_371), .B2(n_369), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_416), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_436), .B(n_374), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_389), .B(n_371), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_421), .B(n_367), .C(n_359), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_395), .A2(n_382), .B(n_364), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_437), .B(n_367), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_431), .Y(n_457) );
NAND2xp33_ASAP7_75t_L g458 ( .A(n_397), .B(n_359), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_425), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_390), .B(n_382), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_425), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_404), .A2(n_382), .B(n_229), .C(n_248), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_391), .B(n_156), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_398), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_398), .Y(n_465) );
AOI221x1_ASAP7_75t_L g466 ( .A1(n_410), .A2(n_156), .B1(n_260), .B2(n_195), .C(n_200), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_399), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_387), .B(n_147), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_399), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_422), .B(n_214), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_396), .B(n_403), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_394), .Y(n_472) );
AOI211x1_ASAP7_75t_L g473 ( .A1(n_414), .A2(n_229), .B(n_21), .C(n_23), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_394), .B(n_147), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_400), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_393), .B(n_151), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_388), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_386), .B(n_20), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_397), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_417), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_418), .A2(n_214), .B1(n_234), .B2(n_151), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_417), .B(n_25), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_415), .A2(n_195), .B(n_227), .C(n_34), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_471), .B(n_429), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_448), .A2(n_447), .B1(n_449), .B2(n_479), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_449), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_459), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_461), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_455), .B(n_429), .Y(n_489) );
AOI21xp33_ASAP7_75t_SL g490 ( .A1(n_445), .A2(n_434), .B(n_419), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_439), .B(n_434), .Y(n_491) );
XNOR2x1_ASAP7_75t_L g492 ( .A(n_475), .B(n_420), .Y(n_492) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_480), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_456), .B(n_408), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_464), .B(n_386), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_450), .Y(n_497) );
XOR2x2_ASAP7_75t_L g498 ( .A(n_470), .B(n_435), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_465), .B(n_405), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_454), .A2(n_426), .B1(n_411), .B2(n_413), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g501 ( .A1(n_441), .A2(n_428), .B1(n_407), .B2(n_427), .C1(n_432), .C2(n_151), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_458), .A2(n_427), .B1(n_428), .B2(n_407), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_478), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_469), .A2(n_428), .B1(n_427), .B2(n_433), .C(n_438), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_472), .B(n_452), .Y(n_506) );
OAI22xp5_ASAP7_75t_SL g507 ( .A1(n_473), .A2(n_430), .B1(n_31), .B2(n_35), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_478), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_440), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_460), .B(n_27), .Y(n_510) );
OAI21xp33_ASAP7_75t_SL g511 ( .A1(n_442), .A2(n_36), .B(n_37), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_443), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_490), .A2(n_481), .B(n_483), .C(n_462), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_495), .B(n_453), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_497), .Y(n_516) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_485), .A2(n_481), .B(n_476), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_L g518 ( .A1(n_489), .A2(n_457), .B(n_451), .C(n_463), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_511), .A2(n_507), .B(n_503), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_509), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_512), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_486), .Y(n_522) );
OAI322xp33_ASAP7_75t_L g523 ( .A1(n_486), .A2(n_476), .A3(n_474), .B1(n_468), .B2(n_482), .C1(n_477), .C2(n_444), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_503), .A2(n_466), .B1(n_151), .B2(n_48), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_508), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g526 ( .A1(n_501), .A2(n_151), .B(n_46), .C(n_49), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_498), .Y(n_527) );
OAI211xp5_ASAP7_75t_SL g528 ( .A1(n_505), .A2(n_39), .B(n_52), .C(n_53), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_513), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_502), .A2(n_56), .B(n_58), .C(n_59), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_494), .Y(n_531) );
NAND2xp33_ASAP7_75t_R g532 ( .A(n_519), .B(n_510), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_517), .A2(n_500), .B1(n_492), .B2(n_491), .C(n_496), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_527), .A2(n_484), .B1(n_504), .B2(n_488), .Y(n_534) );
AND4x1_ASAP7_75t_L g535 ( .A(n_519), .B(n_487), .C(n_506), .D(n_499), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_514), .A2(n_493), .B(n_61), .C(n_64), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_531), .B(n_151), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_518), .A2(n_60), .B(n_66), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_522), .Y(n_539) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_531), .A2(n_68), .B1(n_69), .B2(n_71), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_525), .A2(n_72), .B1(n_73), .B2(n_75), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_539), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_537), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_534), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_533), .B(n_516), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g546 ( .A1(n_536), .A2(n_538), .B(n_526), .C(n_532), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_542), .B(n_535), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_543), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_545), .A2(n_523), .B1(n_528), .B2(n_521), .Y(n_549) );
AOI21xp33_ASAP7_75t_SL g550 ( .A1(n_547), .A2(n_545), .B(n_544), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_548), .Y(n_551) );
OAI22xp5_ASAP7_75t_SL g552 ( .A1(n_551), .A2(n_549), .B1(n_546), .B2(n_541), .Y(n_552) );
INVx4_ASAP7_75t_L g553 ( .A(n_550), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_552), .A2(n_520), .B1(n_529), .B2(n_540), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_554), .A2(n_553), .B(n_530), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_524), .B1(n_515), .B2(n_526), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_556), .A2(n_515), .B1(n_77), .B2(n_78), .Y(n_557) );
endmodule