module real_aes_2485_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_0), .B(n_502), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_1), .A2(n_504), .B(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_2), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_3), .B(n_180), .Y(n_538) );
INVx1_ASAP7_75t_L g135 ( .A(n_4), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_5), .B(n_144), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_6), .B(n_180), .Y(n_526) );
INVx1_ASAP7_75t_L g190 ( .A(n_7), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_8), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_9), .Y(n_206) );
NAND2xp33_ASAP7_75t_L g559 ( .A(n_10), .B(n_177), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_11), .A2(n_492), .B1(n_819), .B2(n_820), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_11), .Y(n_819) );
INVx2_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
AOI221x1_ASAP7_75t_L g583 ( .A1(n_13), .A2(n_26), .B1(n_502), .B2(n_504), .C(n_584), .Y(n_583) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_15), .B(n_502), .Y(n_555) );
INVx1_ASAP7_75t_L g178 ( .A(n_16), .Y(n_178) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_17), .A2(n_166), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_18), .B(n_220), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_19), .B(n_180), .Y(n_515) );
AO21x1_ASAP7_75t_L g533 ( .A1(n_20), .A2(n_502), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_21), .B(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g119 ( .A(n_21), .Y(n_119) );
AOI221xp5_ASAP7_75t_L g111 ( .A1(n_22), .A2(n_112), .B1(n_793), .B2(n_794), .C(n_798), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g793 ( .A(n_22), .Y(n_793) );
INVx1_ASAP7_75t_L g175 ( .A(n_23), .Y(n_175) );
INVx1_ASAP7_75t_SL g250 ( .A(n_24), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_25), .B(n_155), .Y(n_154) );
AOI33xp33_ASAP7_75t_L g227 ( .A1(n_27), .A2(n_55), .A3(n_132), .B1(n_150), .B2(n_228), .B3(n_229), .Y(n_227) );
NAND2x1_ASAP7_75t_L g576 ( .A(n_28), .B(n_180), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_29), .Y(n_799) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_30), .B(n_177), .Y(n_525) );
INVx1_ASAP7_75t_L g199 ( .A(n_31), .Y(n_199) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_32), .A2(n_86), .B(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g145 ( .A(n_32), .B(n_86), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_33), .B(n_188), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_34), .B(n_177), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_35), .B(n_180), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_36), .B(n_177), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_37), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_38), .A2(n_504), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_39), .A2(n_100), .B1(n_109), .B2(n_821), .Y(n_99) );
AND2x2_ASAP7_75t_L g138 ( .A(n_40), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g149 ( .A(n_40), .Y(n_149) );
AND2x2_ASAP7_75t_L g164 ( .A(n_40), .B(n_135), .Y(n_164) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_41), .B(n_106), .C(n_108), .Y(n_105) );
OR2x6_ASAP7_75t_L g117 ( .A(n_41), .B(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_42), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_43), .B(n_502), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_44), .B(n_188), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_45), .A2(n_129), .B1(n_141), .B2(n_144), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_46), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_47), .B(n_155), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_48), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_49), .B(n_177), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_50), .B(n_166), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_51), .B(n_155), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_52), .A2(n_504), .B(n_524), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_53), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_54), .B(n_177), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_56), .B(n_155), .Y(n_218) );
INVx1_ASAP7_75t_L g133 ( .A(n_57), .Y(n_133) );
INVx1_ASAP7_75t_L g157 ( .A(n_57), .Y(n_157) );
AND2x2_ASAP7_75t_L g219 ( .A(n_58), .B(n_220), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g187 ( .A1(n_59), .A2(n_75), .B1(n_147), .B2(n_188), .C(n_189), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_60), .B(n_188), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_61), .B(n_180), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_62), .B(n_141), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g238 ( .A1(n_63), .A2(n_147), .B(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_64), .A2(n_504), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g171 ( .A(n_65), .Y(n_171) );
AO21x1_ASAP7_75t_L g535 ( .A1(n_66), .A2(n_504), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_67), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g217 ( .A(n_68), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_69), .B(n_502), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_70), .A2(n_147), .B(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g549 ( .A(n_71), .B(n_221), .Y(n_549) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
INVx1_ASAP7_75t_L g159 ( .A(n_72), .Y(n_159) );
AND2x2_ASAP7_75t_L g528 ( .A(n_73), .B(n_195), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_74), .B(n_188), .Y(n_230) );
AND2x2_ASAP7_75t_L g252 ( .A(n_76), .B(n_195), .Y(n_252) );
INVx1_ASAP7_75t_L g172 ( .A(n_77), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_78), .A2(n_147), .B(n_249), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_79), .A2(n_147), .B(n_153), .C(n_165), .Y(n_146) );
INVx1_ASAP7_75t_L g104 ( .A(n_80), .Y(n_104) );
AND2x2_ASAP7_75t_L g499 ( .A(n_81), .B(n_195), .Y(n_499) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_82), .B(n_195), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_83), .B(n_502), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_84), .A2(n_147), .B1(n_225), .B2(n_226), .Y(n_224) );
AND2x2_ASAP7_75t_L g534 ( .A(n_85), .B(n_144), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_87), .B(n_177), .Y(n_516) );
AND2x2_ASAP7_75t_L g579 ( .A(n_88), .B(n_195), .Y(n_579) );
INVx1_ASAP7_75t_L g240 ( .A(n_89), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_90), .B(n_180), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_91), .A2(n_504), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_92), .B(n_177), .Y(n_585) );
AND2x2_ASAP7_75t_L g231 ( .A(n_93), .B(n_195), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_94), .B(n_180), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_95), .A2(n_197), .B(n_198), .C(n_200), .Y(n_196) );
BUFx2_ASAP7_75t_SL g815 ( .A(n_96), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_97), .A2(n_504), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_98), .B(n_155), .Y(n_241) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g822 ( .A(n_101), .Y(n_822) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_104), .B(n_119), .Y(n_118) );
OR2x6_ASAP7_75t_SL g115 ( .A(n_108), .B(n_116), .Y(n_115) );
AND2x6_ASAP7_75t_SL g792 ( .A(n_108), .B(n_117), .Y(n_792) );
OR2x2_ASAP7_75t_L g802 ( .A(n_108), .B(n_117), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_108), .B(n_116), .Y(n_810) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_811), .B(n_816), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g110 ( .A(n_111), .B(n_803), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_120), .B1(n_492), .B2(n_791), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_114), .A2(n_120), .B1(n_492), .B2(n_796), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_426), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_349), .Y(n_121) );
NAND3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_296), .C(n_329), .Y(n_122) );
AOI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_253), .B(n_262), .C(n_286), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_182), .B(n_232), .Y(n_124) );
OR2x2_ASAP7_75t_L g306 ( .A(n_125), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g461 ( .A(n_125), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_126), .A2(n_352), .B1(n_356), .B2(n_358), .Y(n_351) );
AND2x2_ASAP7_75t_L g388 ( .A(n_126), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_167), .Y(n_126) );
INVx1_ASAP7_75t_L g285 ( .A(n_127), .Y(n_285) );
AND2x4_ASAP7_75t_L g302 ( .A(n_127), .B(n_283), .Y(n_302) );
INVx2_ASAP7_75t_L g324 ( .A(n_127), .Y(n_324) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_127), .Y(n_407) );
AND2x2_ASAP7_75t_L g478 ( .A(n_127), .B(n_235), .Y(n_478) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_146), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_136), .C(n_140), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g188 ( .A(n_131), .B(n_137), .Y(n_188) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
OR2x6_ASAP7_75t_L g162 ( .A(n_132), .B(n_151), .Y(n_162) );
INVxp33_ASAP7_75t_L g228 ( .A(n_132), .Y(n_228) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g152 ( .A(n_133), .B(n_135), .Y(n_152) );
AND2x4_ASAP7_75t_L g180 ( .A(n_133), .B(n_158), .Y(n_180) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g504 ( .A(n_138), .B(n_152), .Y(n_504) );
INVx2_ASAP7_75t_L g151 ( .A(n_139), .Y(n_151) );
AND2x6_ASAP7_75t_L g177 ( .A(n_139), .B(n_156), .Y(n_177) );
INVx4_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_141), .B(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx4f_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
AND2x4_ASAP7_75t_L g144 ( .A(n_143), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_143), .B(n_145), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_144), .B(n_163), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_144), .A2(n_238), .B(n_242), .Y(n_237) );
INVx1_ASAP7_75t_SL g511 ( .A(n_144), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_144), .B(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_144), .A2(n_555), .B(n_556), .Y(n_554) );
INVxp67_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NOR2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx1_ASAP7_75t_L g229 ( .A(n_150), .Y(n_229) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_160), .B(n_163), .Y(n_153) );
INVx1_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
AND2x4_ASAP7_75t_L g502 ( .A(n_155), .B(n_164), .Y(n_502) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_162), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_162), .A2(n_163), .B(n_190), .C(n_191), .Y(n_189) );
INVxp67_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_162), .A2(n_163), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_162), .A2(n_163), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_162), .A2(n_163), .B(n_250), .C(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_163), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_163), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_163), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_163), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_163), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_163), .A2(n_558), .B(n_559), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_163), .A2(n_576), .B(n_577), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_163), .A2(n_585), .B(n_586), .Y(n_584) );
INVx5_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_165), .A2(n_223), .B(n_231), .Y(n_222) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_165), .A2(n_223), .B(n_231), .Y(n_267) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_166), .A2(n_187), .B(n_192), .Y(n_186) );
AND2x2_ASAP7_75t_L g243 ( .A(n_167), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g272 ( .A(n_167), .Y(n_272) );
INVx3_ASAP7_75t_L g283 ( .A(n_167), .Y(n_283) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_174), .B(n_181), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_173), .B(n_199), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B1(n_178), .B2(n_179), .Y(n_174) );
INVxp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_182), .A2(n_473), .B1(n_475), .B2(n_477), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_182), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_210), .Y(n_183) );
INVx3_ASAP7_75t_L g256 ( .A(n_184), .Y(n_256) );
AND2x2_ASAP7_75t_L g264 ( .A(n_184), .B(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_184), .Y(n_294) );
NAND2x1_ASAP7_75t_SL g488 ( .A(n_184), .B(n_255), .Y(n_488) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_193), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g261 ( .A(n_186), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_186), .B(n_267), .Y(n_279) );
AND2x2_ASAP7_75t_L g292 ( .A(n_186), .B(n_193), .Y(n_292) );
AND2x4_ASAP7_75t_L g299 ( .A(n_186), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_186), .Y(n_348) );
INVxp67_ASAP7_75t_L g355 ( .A(n_186), .Y(n_355) );
INVx1_ASAP7_75t_L g360 ( .A(n_186), .Y(n_360) );
INVx1_ASAP7_75t_L g209 ( .A(n_188), .Y(n_209) );
INVx1_ASAP7_75t_L g259 ( .A(n_193), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_193), .B(n_269), .Y(n_278) );
INVx2_ASAP7_75t_L g346 ( .A(n_193), .Y(n_346) );
INVx1_ASAP7_75t_L g385 ( .A(n_193), .Y(n_385) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_201), .B2(n_202), .Y(n_194) );
INVx3_ASAP7_75t_L g202 ( .A(n_195), .Y(n_202) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_202), .A2(n_213), .B(n_219), .Y(n_212) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_202), .A2(n_213), .B(n_219), .Y(n_269) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_202), .A2(n_543), .B(n_549), .Y(n_542) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_202), .A2(n_543), .B(n_549), .Y(n_564) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_202), .A2(n_573), .B(n_579), .Y(n_572) );
AO21x2_ASAP7_75t_L g597 ( .A1(n_202), .A2(n_573), .B(n_579), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g315 ( .A(n_210), .B(n_292), .Y(n_315) );
AND2x2_ASAP7_75t_L g383 ( .A(n_210), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g397 ( .A(n_210), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_210), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_222), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_212), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g353 ( .A(n_212), .B(n_346), .Y(n_353) );
AND2x2_ASAP7_75t_L g444 ( .A(n_212), .B(n_266), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_220), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_220), .A2(n_501), .B(n_503), .Y(n_500) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_220), .A2(n_583), .B(n_587), .Y(n_582) );
OA21x2_ASAP7_75t_L g627 ( .A1(n_220), .A2(n_583), .B(n_587), .Y(n_627) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
INVx2_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
AND2x2_ASAP7_75t_L g345 ( .A(n_222), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_224), .B(n_230), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_243), .Y(n_233) );
AND2x2_ASAP7_75t_L g387 ( .A(n_234), .B(n_388), .Y(n_387) );
OR2x6_ASAP7_75t_L g446 ( .A(n_234), .B(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g276 ( .A(n_235), .Y(n_276) );
AND2x4_ASAP7_75t_L g284 ( .A(n_235), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g319 ( .A(n_235), .B(n_244), .Y(n_319) );
INVx2_ASAP7_75t_L g368 ( .A(n_235), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_235), .B(n_342), .Y(n_417) );
AND2x2_ASAP7_75t_L g454 ( .A(n_235), .B(n_272), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_235), .B(n_337), .Y(n_462) );
OR2x6_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AND2x2_ASAP7_75t_L g295 ( .A(n_243), .B(n_284), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_243), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_243), .B(n_322), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_243), .B(n_335), .Y(n_456) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_244), .Y(n_274) );
AND2x2_ASAP7_75t_L g282 ( .A(n_244), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
INVx2_ASAP7_75t_L g308 ( .A(n_244), .Y(n_308) );
INVx1_ASAP7_75t_L g341 ( .A(n_244), .Y(n_341) );
INVx1_ASAP7_75t_L g389 ( .A(n_244), .Y(n_389) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_252), .Y(n_244) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_245), .A2(n_522), .B(n_528), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_255), .B(n_258), .Y(n_331) );
OR2x2_ASAP7_75t_L g403 ( .A(n_255), .B(n_404), .Y(n_403) );
AND4x1_ASAP7_75t_SL g449 ( .A(n_255), .B(n_431), .C(n_450), .D(n_451), .Y(n_449) );
OR2x2_ASAP7_75t_L g473 ( .A(n_256), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g310 ( .A(n_259), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_259), .B(n_268), .Y(n_460) );
AND2x2_ASAP7_75t_L g485 ( .A(n_260), .B(n_345), .Y(n_485) );
OAI32xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_270), .A3(n_275), .B1(n_277), .B2(n_280), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g358 ( .A(n_265), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g458 ( .A(n_265), .B(n_412), .Y(n_458) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x2_ASAP7_75t_L g354 ( .A(n_266), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g440 ( .A(n_266), .Y(n_440) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_267), .B(n_269), .Y(n_474) );
INVx3_ASAP7_75t_L g291 ( .A(n_268), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_268), .B(n_396), .Y(n_469) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
AND2x2_ASAP7_75t_L g347 ( .A(n_269), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g481 ( .A(n_271), .Y(n_481) );
NAND2x1_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g321 ( .A(n_272), .Y(n_321) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_272), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_275), .B(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g313 ( .A(n_276), .B(n_281), .Y(n_313) );
AND2x4_ASAP7_75t_L g335 ( .A(n_276), .B(n_285), .Y(n_335) );
AND2x4_ASAP7_75t_SL g406 ( .A(n_276), .B(n_407), .Y(n_406) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_276), .B(n_357), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_277), .A2(n_400), .B1(n_403), .B2(n_405), .Y(n_399) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_SL g419 ( .A(n_278), .Y(n_419) );
INVx2_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_282), .B(n_288), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_282), .A2(n_418), .B1(n_421), .B2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g342 ( .A(n_283), .Y(n_342) );
AND2x2_ASAP7_75t_L g365 ( .A(n_283), .B(n_324), .Y(n_365) );
INVx2_ASAP7_75t_L g288 ( .A(n_284), .Y(n_288) );
OAI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_289), .B(n_293), .Y(n_286) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_290), .A2(n_362), .B1(n_366), .B2(n_367), .Y(n_361) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_291), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_291), .B(n_359), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_291), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NOR3xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_312), .C(n_316), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_306), .B2(n_309), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g326 ( .A(n_299), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g366 ( .A(n_299), .B(n_353), .Y(n_366) );
AND2x2_ASAP7_75t_L g418 ( .A(n_299), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g435 ( .A(n_299), .B(n_385), .Y(n_435) );
AND2x2_ASAP7_75t_L g490 ( .A(n_299), .B(n_384), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx4_ASAP7_75t_L g357 ( .A(n_302), .Y(n_357) );
AND2x2_ASAP7_75t_L g367 ( .A(n_302), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g372 ( .A(n_305), .Y(n_372) );
AND2x2_ASAP7_75t_L g381 ( .A(n_305), .B(n_365), .Y(n_381) );
INVx1_ASAP7_75t_L g416 ( .A(n_307), .Y(n_416) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_310), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_311), .B(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B(n_325), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_318), .B(n_357), .Y(n_466) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AOI21xp33_ASAP7_75t_SL g329 ( .A1(n_321), .A2(n_330), .B(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g476 ( .A(n_321), .B(n_335), .Y(n_476) );
AND2x4_ASAP7_75t_L g339 ( .A(n_322), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_SL g373 ( .A(n_322), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_322), .B(n_389), .Y(n_455) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_338), .B(n_343), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_335), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_335), .B(n_340), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_336), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g398 ( .A(n_336), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_336), .Y(n_402) );
AND2x2_ASAP7_75t_L g486 ( .A(n_336), .B(n_454), .Y(n_486) );
AND2x2_ASAP7_75t_L g489 ( .A(n_336), .B(n_406), .Y(n_489) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_SL g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_341), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g468 ( .A(n_345), .Y(n_468) );
AND2x2_ASAP7_75t_L g359 ( .A(n_346), .B(n_360), .Y(n_359) );
NAND4xp75_ASAP7_75t_L g349 ( .A(n_350), .B(n_369), .C(n_390), .D(n_408), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_361), .Y(n_350) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_353), .B(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_354), .B(n_419), .Y(n_425) );
NAND2xp5_ASAP7_75t_R g441 ( .A(n_357), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g491 ( .A(n_357), .Y(n_491) );
INVx2_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
BUFx3_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g447 ( .A(n_365), .Y(n_447) );
AND2x2_ASAP7_75t_L g401 ( .A(n_367), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g423 ( .A(n_368), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B(n_376), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_372), .B(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_373), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_375), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B1(n_382), .B2(n_386), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OA21x2_ASAP7_75t_L g391 ( .A1(n_384), .A2(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g412 ( .A(n_384), .Y(n_412) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g443 ( .A(n_385), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g451 ( .A(n_385), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_386), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g421 ( .A(n_389), .B(n_422), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_397), .B(n_399), .Y(n_390) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g438 ( .A(n_395), .B(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
INVx2_ASAP7_75t_SL g442 ( .A(n_406), .Y(n_442) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_420), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_413), .B1(n_415), .B2(n_418), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g471 ( .A(n_415), .Y(n_471) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_463), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_436), .C(n_448), .Y(n_427) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_441), .B1(n_443), .B2(n_445), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .C(n_459), .Y(n_448) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .B(n_457), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_482), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_472), .C(n_479), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_470), .B2(n_471), .Y(n_465) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_473), .B(n_478), .C(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B1(n_487), .B2(n_489), .C1(n_490), .C2(n_491), .Y(n_482) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g820 ( .A(n_492), .Y(n_820) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_676), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_631), .C(n_660), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_495), .B(n_604), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_529), .B1(n_550), .B2(n_561), .C(n_565), .Y(n_495) );
INVx3_ASAP7_75t_SL g721 ( .A(n_496), .Y(n_721) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_497), .B(n_508), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g567 ( .A(n_497), .B(n_520), .Y(n_567) );
INVx4_ASAP7_75t_L g602 ( .A(n_497), .Y(n_602) );
AND2x2_ASAP7_75t_L g624 ( .A(n_497), .B(n_521), .Y(n_624) );
AND2x2_ASAP7_75t_L g630 ( .A(n_497), .B(n_569), .Y(n_630) );
INVx5_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g599 ( .A(n_498), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_498), .B(n_520), .Y(n_675) );
AND2x2_ASAP7_75t_L g680 ( .A(n_498), .B(n_521), .Y(n_680) );
AND2x2_ASAP7_75t_L g692 ( .A(n_498), .B(n_553), .Y(n_692) );
NOR2x1_ASAP7_75t_SL g731 ( .A(n_498), .B(n_569), .Y(n_731) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g560 ( .A(n_508), .Y(n_560) );
AND2x2_ASAP7_75t_L g664 ( .A(n_508), .B(n_613), .Y(n_664) );
AND2x2_ASAP7_75t_L g761 ( .A(n_508), .B(n_692), .Y(n_761) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_520), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g593 ( .A(n_510), .Y(n_593) );
INVx2_ASAP7_75t_L g615 ( .A(n_510), .Y(n_615) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_511), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
AND2x2_ASAP7_75t_L g590 ( .A(n_520), .B(n_552), .Y(n_590) );
INVx2_ASAP7_75t_L g594 ( .A(n_520), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_520), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g693 ( .A(n_520), .B(n_658), .Y(n_693) );
OR2x2_ASAP7_75t_L g740 ( .A(n_520), .B(n_553), .Y(n_740) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_521), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
AND2x2_ASAP7_75t_L g737 ( .A(n_529), .B(n_618), .Y(n_737) );
AND2x2_ASAP7_75t_L g787 ( .A(n_529), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g663 ( .A(n_530), .B(n_607), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_541), .Y(n_530) );
AND2x2_ASAP7_75t_L g596 ( .A(n_531), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g626 ( .A(n_531), .B(n_627), .Y(n_626) );
AND2x4_ASAP7_75t_L g647 ( .A(n_531), .B(n_627), .Y(n_647) );
AND2x4_ASAP7_75t_L g682 ( .A(n_531), .B(n_670), .Y(n_682) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g563 ( .A(n_532), .Y(n_563) );
OAI21x1_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_535), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g540 ( .A(n_534), .Y(n_540) );
AND2x2_ASAP7_75t_L g609 ( .A(n_541), .B(n_562), .Y(n_609) );
AND2x2_ASAP7_75t_L g695 ( .A(n_541), .B(n_627), .Y(n_695) );
AND2x2_ASAP7_75t_L g706 ( .A(n_541), .B(n_571), .Y(n_706) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g570 ( .A(n_542), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g637 ( .A(n_542), .B(n_572), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_548), .Y(n_543) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_560), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_552), .B(n_602), .Y(n_659) );
AND2x2_ASAP7_75t_L g703 ( .A(n_552), .B(n_569), .Y(n_703) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_553), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g613 ( .A(n_553), .Y(n_613) );
BUFx3_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
AND2x2_ASAP7_75t_L g645 ( .A(n_553), .B(n_615), .Y(n_645) );
OAI322xp33_ASAP7_75t_L g565 ( .A1(n_560), .A2(n_566), .A3(n_570), .B1(n_580), .B2(n_588), .C1(n_595), .C2(n_600), .Y(n_565) );
INVx1_ASAP7_75t_L g726 ( .A(n_560), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_561), .B(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g639 ( .A(n_561), .B(n_581), .Y(n_639) );
INVx2_ASAP7_75t_L g684 ( .A(n_561), .Y(n_684) );
AND2x2_ASAP7_75t_L g700 ( .A(n_561), .B(n_642), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_561), .B(n_718), .Y(n_748) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_562), .B(n_627), .Y(n_651) );
OR2x2_ASAP7_75t_L g672 ( .A(n_562), .B(n_589), .Y(n_672) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g644 ( .A(n_563), .Y(n_644) );
INVx2_ASAP7_75t_L g589 ( .A(n_564), .Y(n_589) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_564), .Y(n_591) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g634 ( .A(n_567), .Y(n_634) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_568), .Y(n_654) );
INVx1_ASAP7_75t_L g752 ( .A(n_568), .Y(n_752) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_568), .Y(n_767) );
NAND2x1_ASAP7_75t_L g777 ( .A(n_570), .B(n_581), .Y(n_777) );
INVx1_ASAP7_75t_L g784 ( .A(n_570), .Y(n_784) );
BUFx2_ASAP7_75t_L g618 ( .A(n_571), .Y(n_618) );
AND2x2_ASAP7_75t_L g694 ( .A(n_571), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
INVxp67_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_580), .B(n_596), .C(n_598), .Y(n_595) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_SL g616 ( .A(n_581), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_581), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g768 ( .A(n_581), .B(n_717), .Y(n_768) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g670 ( .A(n_582), .Y(n_670) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_582), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_591), .B2(n_592), .Y(n_588) );
AND2x4_ASAP7_75t_SL g717 ( .A(n_589), .B(n_597), .Y(n_717) );
AND2x2_ASAP7_75t_L g730 ( .A(n_590), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_591), .Y(n_732) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_L g689 ( .A(n_593), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_593), .B(n_602), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_594), .B(n_612), .Y(n_611) );
AND3x2_ASAP7_75t_L g629 ( .A(n_594), .B(n_622), .C(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g653 ( .A(n_594), .Y(n_653) );
AND2x2_ASAP7_75t_L g766 ( .A(n_594), .B(n_767), .Y(n_766) );
BUFx2_ASAP7_75t_L g642 ( .A(n_597), .Y(n_642) );
INVx1_ASAP7_75t_L g720 ( .A(n_597), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_598), .B(n_621), .Y(n_759) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_599), .B(n_703), .Y(n_708) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g699 ( .A(n_602), .B(n_645), .Y(n_699) );
INVx1_ASAP7_75t_SL g650 ( .A(n_603), .Y(n_650) );
AND2x2_ASAP7_75t_L g758 ( .A(n_603), .B(n_670), .Y(n_758) );
AND2x2_ASAP7_75t_L g779 ( .A(n_603), .B(n_651), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_610), .B1(n_616), .B2(n_619), .C(n_625), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g771 ( .A(n_607), .Y(n_771) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_608), .A2(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g617 ( .A(n_609), .B(n_618), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g640 ( .A1(n_609), .A2(n_641), .B1(n_643), .B2(n_648), .C1(n_652), .C2(n_655), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_609), .B(n_758), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_610), .A2(n_639), .B1(n_662), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g646 ( .A(n_613), .Y(n_646) );
AND2x2_ASAP7_75t_L g765 ( .A(n_613), .B(n_731), .Y(n_765) );
OAI32xp33_ASAP7_75t_L g769 ( .A1(n_613), .A2(n_638), .A3(n_690), .B1(n_698), .B2(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g774 ( .A(n_613), .B(n_624), .Y(n_774) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g658 ( .A(n_615), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_616), .A2(n_666), .B(n_673), .Y(n_665) );
INVx1_ASAP7_75t_L g729 ( .A(n_618), .Y(n_729) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
AND2x2_ASAP7_75t_L g633 ( .A(n_621), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g641 ( .A(n_624), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g714 ( .A(n_624), .B(n_645), .Y(n_714) );
INVx1_ASAP7_75t_SL g785 ( .A(n_626), .Y(n_785) );
AND2x2_ASAP7_75t_L g719 ( .A(n_627), .B(n_720), .Y(n_719) );
OAI222xp33_ASAP7_75t_L g772 ( .A1(n_628), .A2(n_681), .B1(n_760), .B2(n_773), .C1(n_775), .C2(n_777), .Y(n_772) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g745 ( .A(n_630), .B(n_746), .Y(n_745) );
OAI21xp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_635), .B(n_640), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_634), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g713 ( .A(n_636), .Y(n_713) );
INVx1_ASAP7_75t_L g681 ( .A(n_637), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_637), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g735 ( .A(n_642), .Y(n_735) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_646), .B2(n_647), .Y(n_643) );
OAI322xp33_ASAP7_75t_L g755 ( .A1(n_644), .A2(n_705), .A3(n_708), .B1(n_756), .B2(n_757), .C1(n_759), .C2(n_760), .Y(n_755) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_645), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g674 ( .A(n_646), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_647), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g776 ( .A(n_647), .B(n_706), .Y(n_776) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g756 ( .A(n_650), .Y(n_756) );
INVx1_ASAP7_75t_SL g685 ( .A(n_651), .Y(n_685) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
OR2x2_ASAP7_75t_L g687 ( .A(n_659), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g725 ( .A(n_659), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g698 ( .A(n_669), .B(n_684), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_669), .B(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g728 ( .A(n_672), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_741), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_696), .C(n_709), .D(n_722), .Y(n_677) );
AOI322xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .A3(n_682), .B1(n_683), .B2(n_686), .C1(n_691), .C2(n_694), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g778 ( .A1(n_679), .A2(n_779), .B(n_780), .C(n_783), .Y(n_778) );
AND2x2_ASAP7_75t_L g790 ( .A(n_680), .B(n_767), .Y(n_790) );
INVx1_ASAP7_75t_L g712 ( .A(n_682), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_682), .B(n_717), .Y(n_754) );
NAND2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_690), .B(n_703), .Y(n_770) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B1(n_700), .B2(n_701), .C1(n_704), .C2(n_707), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_699), .A2(n_710), .B1(n_713), .B2(n_714), .C(n_715), .Y(n_709) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp33_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_718), .B(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_727), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g782 ( .A(n_731), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_736), .B(n_738), .Y(n_733) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g746 ( .A(n_740), .Y(n_746) );
OR2x2_ASAP7_75t_L g781 ( .A(n_740), .B(n_782), .Y(n_781) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_762), .C(n_778), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_755), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_747), .B(n_749), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_768), .B1(n_769), .B2(n_771), .C(n_772), .Y(n_762) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_777), .B(n_781), .Y(n_780) );
O2A1O1Ixp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B(n_786), .C(n_789), .Y(n_783) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_792), .Y(n_797) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx2_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVxp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_804), .A2(n_809), .B(n_818), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_813), .B(n_817), .Y(n_816) );
CKINVDCx11_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
CKINVDCx8_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
endmodule