module real_aes_10609_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
AOI22xp33_ASAP7_75t_SL g27 ( .A1(n_0), .A2(n_7), .B1(n_28), .B2(n_35), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_1), .Y(n_21) );
NOR4xp25_ASAP7_75t_SL g32 ( .A(n_1), .B(n_25), .C(n_33), .D(n_34), .Y(n_32) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_2), .B(n_12), .C(n_19), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_2), .B(n_9), .C(n_24), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_3), .B(n_6), .Y(n_20) );
NAND2xp33_ASAP7_75t_R g24 ( .A(n_4), .B(n_20), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_5), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g31 ( .A(n_8), .B(n_13), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g38 ( .A(n_8), .B(n_26), .Y(n_38) );
NAND2xp33_ASAP7_75t_SL g41 ( .A(n_8), .B(n_26), .Y(n_41) );
NAND2xp33_ASAP7_75t_R g45 ( .A(n_8), .B(n_13), .Y(n_45) );
AOI22xp33_ASAP7_75t_L g39 ( .A1(n_10), .A2(n_11), .B1(n_40), .B2(n_43), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_12), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_13), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g14 ( .A(n_15), .B(n_27), .C(n_39), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g15 ( .A(n_16), .B(n_26), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_17), .B(n_22), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_21), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g22 ( .A(n_23), .B(n_25), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_23), .Y(n_33) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_30), .Y(n_29) );
NAND2xp33_ASAP7_75t_R g30 ( .A(n_31), .B(n_32), .Y(n_30) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_32), .B(n_38), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_32), .Y(n_42) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
NOR2xp33_ASAP7_75t_R g40 ( .A(n_41), .B(n_42), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g44 ( .A(n_42), .B(n_45), .Y(n_44) );
HB1xp67_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
endmodule