module fake_jpeg_24591_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx2_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_33),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_27),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_44),
.B1(n_23),
.B2(n_29),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_20),
.B(n_18),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_21),
.B1(n_23),
.B2(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_87),
.Y(n_97)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_87),
.B1(n_31),
.B2(n_18),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_24),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_88),
.Y(n_108)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_52),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_93),
.Y(n_134)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_115),
.B1(n_73),
.B2(n_69),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_54),
.B1(n_55),
.B2(n_52),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_84),
.B1(n_90),
.B2(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_109),
.B1(n_84),
.B2(n_82),
.Y(n_137)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_21),
.Y(n_105)
);

NAND2x1_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_22),
.Y(n_138)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_83),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_15),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_39),
.B(n_58),
.C(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_17),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_124),
.B1(n_129),
.B2(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_126),
.B1(n_130),
.B2(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_31),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_36),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_99),
.C(n_32),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_35),
.B(n_34),
.C(n_36),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_68),
.B1(n_86),
.B2(n_85),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_24),
.B1(n_73),
.B2(n_56),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_62),
.B1(n_67),
.B2(n_82),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_140),
.B(n_65),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_112),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_32),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_105),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_106),
.B1(n_115),
.B2(n_91),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_23),
.B1(n_17),
.B2(n_19),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_102),
.C(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_102),
.C(n_35),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_155),
.C(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_162),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_36),
.C(n_114),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_118),
.A2(n_93),
.B1(n_107),
.B2(n_95),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_128),
.B1(n_125),
.B2(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_166),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_133),
.B(n_123),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_114),
.C(n_94),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_131),
.B(n_30),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_15),
.A3(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_190),
.B1(n_147),
.B2(n_145),
.Y(n_194)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_175),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_138),
.B(n_140),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_174),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_17),
.B1(n_65),
.B2(n_22),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_127),
.C(n_122),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_185),
.C(n_192),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_184),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_150),
.C(n_142),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_R g186 ( 
.A1(n_160),
.A2(n_132),
.B1(n_135),
.B2(n_122),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_147),
.B1(n_151),
.B2(n_148),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_26),
.B(n_19),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_132),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_22),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_89),
.B1(n_17),
.B2(n_26),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_25),
.B1(n_12),
.B2(n_11),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_111),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_195),
.B1(n_211),
.B2(n_216),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_155),
.C(n_154),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_203),
.C(n_206),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_22),
.C(n_25),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_22),
.C(n_25),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_25),
.C(n_26),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_214),
.C(n_177),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_14),
.B(n_13),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_25),
.C(n_1),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_228),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_220),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_192),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_208),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_196),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_235),
.B1(n_236),
.B2(n_211),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_193),
.C(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_189),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_226),
.A2(n_187),
.B1(n_195),
.B2(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_243),
.C(n_246),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_193),
.C(n_203),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_248),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_247),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_177),
.C(n_214),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_196),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_228),
.A2(n_187),
.B1(n_169),
.B2(n_210),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_223),
.C(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_231),
.C(n_224),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_174),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_168),
.B1(n_191),
.B2(n_171),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_253),
.B1(n_237),
.B2(n_219),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_175),
.B1(n_171),
.B2(n_168),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_204),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_190),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_227),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_270),
.C(n_242),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_268),
.B1(n_271),
.B2(n_244),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_222),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_263),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_230),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_220),
.CI(n_232),
.CON(n_264),
.SN(n_264)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_3),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_238),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_182),
.B1(n_12),
.B2(n_10),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_0),
.C(n_2),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_281),
.B1(n_284),
.B2(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_276),
.B(n_277),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_279),
.C(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_243),
.C(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_255),
.B(n_9),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_285),
.B(n_3),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_286),
.C(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_3),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_278),
.B(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_266),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_4),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_274),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_4),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_264),
.C(n_265),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_300),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_3),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_293),
.C(n_294),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_302),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_288),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_309),
.B(n_310),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_308),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_311),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_312),
.B1(n_298),
.B2(n_8),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_6),
.B(n_7),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_6),
.B(n_317),
.Y(n_320)
);


endmodule