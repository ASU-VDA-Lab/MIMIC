module fake_netlist_1_11599_n_28 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_10), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_7), .B(n_11), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_2), .B(n_3), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_13), .Y(n_19) );
INVx5_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
OA21x2_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_18), .B(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .B1(n_17), .B2(n_14), .C(n_16), .Y(n_23) );
NAND3xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_17), .C(n_14), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_14), .B1(n_1), .B2(n_2), .Y(n_25) );
OAI221xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_0), .B1(n_1), .B2(n_4), .C(n_5), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_24), .Y(n_27) );
XNOR2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_0), .Y(n_28) );
endmodule