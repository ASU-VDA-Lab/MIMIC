module fake_jpeg_30702_n_550 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_550);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_59),
.B(n_91),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_73),
.Y(n_133)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_9),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_86),
.Y(n_130)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_9),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_94),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_83),
.Y(n_149)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_9),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_33),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_9),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_30),
.B(n_11),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_35),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_19),
.Y(n_128)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_106),
.B(n_128),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_112),
.B(n_115),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_26),
.B1(n_21),
.B2(n_22),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_34),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_67),
.A2(n_26),
.B1(n_47),
.B2(n_19),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_122),
.A2(n_139),
.B1(n_142),
.B2(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_136),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_66),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_87),
.B1(n_61),
.B2(n_103),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_38),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_47),
.B1(n_19),
.B2(n_45),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_71),
.A2(n_19),
.B1(n_45),
.B2(n_20),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_73),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_143),
.B(n_50),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_65),
.B(n_21),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_41),
.B1(n_36),
.B2(n_22),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_176),
.B1(n_188),
.B2(n_190),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_92),
.B1(n_98),
.B2(n_96),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_171),
.A2(n_196),
.B1(n_210),
.B2(n_219),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_89),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_172),
.B(n_177),
.Y(n_236)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_90),
.B1(n_79),
.B2(n_82),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_120),
.B(n_52),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_163),
.Y(n_178)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_178),
.Y(n_279)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_107),
.A2(n_36),
.B1(n_41),
.B2(n_23),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_119),
.A2(n_20),
.B1(n_23),
.B2(n_38),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g281 ( 
.A1(n_183),
.A2(n_218),
.B1(n_224),
.B2(n_3),
.Y(n_281)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_116),
.A2(n_55),
.B1(n_57),
.B2(n_53),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_205),
.B1(n_217),
.B2(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_129),
.B1(n_142),
.B2(n_139),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_130),
.A2(n_54),
.B1(n_60),
.B2(n_69),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_163),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_193),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_144),
.A2(n_42),
.B(n_83),
.C(n_89),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_194),
.B(n_166),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_133),
.A2(n_45),
.B1(n_83),
.B2(n_42),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_202),
.Y(n_247)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_121),
.A2(n_134),
.B1(n_123),
.B2(n_168),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_208),
.B1(n_212),
.B2(n_149),
.Y(n_244)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_204),
.Y(n_255)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_135),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_116),
.A2(n_45),
.B1(n_42),
.B2(n_12),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_206),
.B(n_209),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_42),
.B1(n_50),
.B2(n_12),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_211),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_160),
.A2(n_42),
.B1(n_50),
.B2(n_11),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_11),
.B1(n_18),
.B2(n_17),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_230),
.B1(n_1),
.B2(n_2),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_216),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_125),
.A2(n_11),
.B1(n_18),
.B2(n_17),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_127),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_223),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_227),
.B1(n_228),
.B2(n_169),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_132),
.A2(n_8),
.B1(n_18),
.B2(n_17),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_149),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_226),
.B(n_229),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_138),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_127),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_172),
.A2(n_194),
.B(n_173),
.C(n_188),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_232),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_118),
.B1(n_117),
.B2(n_154),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_235),
.A2(n_261),
.B1(n_270),
.B2(n_274),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_244),
.A2(n_268),
.B1(n_201),
.B2(n_186),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_175),
.A2(n_147),
.B1(n_124),
.B2(n_166),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_248),
.A2(n_259),
.B(n_264),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_175),
.B(n_157),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_257),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_175),
.A2(n_105),
.B(n_162),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_177),
.C(n_212),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_180),
.B(n_118),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_264),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_170),
.A2(n_117),
.B1(n_162),
.B2(n_105),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_277),
.B1(n_278),
.B2(n_282),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_183),
.B(n_159),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_159),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_266),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_159),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_172),
.A2(n_50),
.B1(n_8),
.B2(n_13),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_172),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_218),
.B(n_1),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_3),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_207),
.B(n_8),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_193),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_202),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_177),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_195),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_281),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_223),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_236),
.Y(n_285)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_224),
.B1(n_214),
.B2(n_174),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_286),
.A2(n_290),
.B1(n_321),
.B2(n_324),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_289),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_248),
.A2(n_209),
.B1(n_210),
.B2(n_206),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_288),
.A2(n_315),
.B1(n_260),
.B2(n_243),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_247),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_239),
.B1(n_271),
.B2(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_293),
.Y(n_342)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_294),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_185),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_298),
.Y(n_331)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_182),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_309),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_236),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_308),
.Y(n_334)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_303),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_230),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_307),
.C(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_306),
.B(n_317),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_200),
.C(n_179),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_237),
.B(n_184),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_237),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_265),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_314),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_213),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_316),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_256),
.B(n_235),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_246),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_275),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_228),
.B1(n_227),
.B2(n_221),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_189),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_318),
.B(n_319),
.Y(n_361)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_239),
.A2(n_193),
.B1(n_178),
.B2(n_198),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_323),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_250),
.B(n_216),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_232),
.A2(n_181),
.B1(n_191),
.B2(n_192),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_276),
.A2(n_203),
.B1(n_204),
.B2(n_6),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_238),
.B1(n_269),
.B2(n_241),
.Y(n_332)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_328),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_6),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_234),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_258),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_332),
.A2(n_326),
.B(n_325),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_SL g337 ( 
.A(n_318),
.B(n_232),
.C(n_268),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_SL g383 ( 
.A(n_337),
.B(n_322),
.C(n_313),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_339),
.B(n_343),
.Y(n_392)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_233),
.B1(n_270),
.B2(n_244),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_341),
.A2(n_347),
.B1(n_353),
.B2(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_310),
.A2(n_233),
.B1(n_277),
.B2(n_275),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_351),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_298),
.B(n_273),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_346),
.B(n_369),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_290),
.A2(n_255),
.B1(n_242),
.B2(n_280),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_303),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_312),
.A2(n_280),
.B1(n_242),
.B2(n_241),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_316),
.A2(n_301),
.B1(n_328),
.B2(n_296),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_360),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_301),
.A2(n_231),
.B1(n_243),
.B2(n_241),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_308),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_359),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_296),
.A2(n_231),
.B1(n_245),
.B2(n_267),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_324),
.A2(n_245),
.B1(n_269),
.B2(n_267),
.Y(n_362)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_363),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_279),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_364),
.B(n_365),
.Y(n_402)
);

FAx1_ASAP7_75t_SL g365 ( 
.A(n_283),
.B(n_279),
.CI(n_258),
.CON(n_365),
.SN(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_321),
.A2(n_305),
.B1(n_320),
.B2(n_284),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_366),
.A2(n_370),
.B1(n_288),
.B2(n_322),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_304),
.B(n_283),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_368),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_299),
.A2(n_238),
.B1(n_240),
.B2(n_254),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_295),
.B(n_240),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_284),
.A2(n_311),
.B1(n_322),
.B2(n_314),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_285),
.C(n_302),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_387),
.C(n_392),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_354),
.A2(n_291),
.B(n_285),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_372),
.A2(n_364),
.B(n_338),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_291),
.B1(n_315),
.B2(n_299),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_378),
.B1(n_379),
.B2(n_388),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_341),
.A2(n_304),
.B1(n_302),
.B2(n_287),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_330),
.A2(n_289),
.B1(n_322),
.B2(n_293),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_381),
.Y(n_415)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_383),
.A2(n_405),
.B(n_333),
.Y(n_432)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_398),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_339),
.B(n_307),
.C(n_313),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_335),
.A2(n_306),
.B1(n_286),
.B2(n_327),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_391),
.B1(n_394),
.B2(n_351),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_335),
.A2(n_319),
.B1(n_317),
.B2(n_300),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_393),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_366),
.A2(n_292),
.B1(n_297),
.B2(n_238),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_348),
.Y(n_395)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_395),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_364),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_401),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_336),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_403),
.A2(n_336),
.B1(n_369),
.B2(n_331),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_404),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_SL g405 ( 
.A1(n_337),
.A2(n_303),
.B(n_279),
.C(n_329),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_406),
.B(n_407),
.C(n_424),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_339),
.C(n_343),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_376),
.A2(n_354),
.B1(n_330),
.B2(n_359),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_414),
.B1(n_418),
.B2(n_375),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_361),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_411),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_343),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_376),
.A2(n_330),
.B1(n_355),
.B2(n_347),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_367),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_425),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_375),
.A2(n_355),
.B1(n_356),
.B2(n_362),
.Y(n_418)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_384),
.A2(n_331),
.B1(n_346),
.B2(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_334),
.C(n_372),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_334),
.Y(n_425)
);

A2O1A1O1Ixp25_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_405),
.B(n_393),
.C(n_389),
.D(n_357),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_333),
.C(n_338),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_428),
.B(n_437),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_429),
.A2(n_436),
.B1(n_391),
.B2(n_401),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_365),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_402),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_432),
.Y(n_440)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_380),
.B(n_352),
.CI(n_365),
.CON(n_434),
.SN(n_434)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_380),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_402),
.A2(n_353),
.B(n_365),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_435),
.A2(n_405),
.B(n_399),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_373),
.A2(n_345),
.B1(n_360),
.B2(n_340),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_368),
.C(n_344),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_439),
.A2(n_448),
.B1(n_449),
.B2(n_436),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_461),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_443),
.A2(n_451),
.B1(n_457),
.B2(n_458),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_412),
.A2(n_385),
.B1(n_396),
.B2(n_384),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_444),
.Y(n_485)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_417),
.A2(n_388),
.B1(n_374),
.B2(n_394),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_374),
.B1(n_396),
.B2(n_398),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_409),
.Y(n_450)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_431),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_397),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_454),
.C(n_424),
.Y(n_468)
);

AO22x2_ASAP7_75t_L g453 ( 
.A1(n_432),
.A2(n_398),
.B1(n_381),
.B2(n_377),
.Y(n_453)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_397),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_417),
.A2(n_405),
.B(n_377),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_455),
.A2(n_405),
.B(n_415),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_390),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_459),
.A2(n_426),
.B1(n_437),
.B2(n_413),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_462),
.B(n_463),
.CI(n_464),
.CON(n_484),
.SN(n_484)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_433),
.B(n_357),
.C(n_395),
.Y(n_463)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_465),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_466),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_486),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_469),
.A2(n_472),
.B1(n_474),
.B2(n_481),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_456),
.C(n_406),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_475),
.C(n_477),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_445),
.A2(n_412),
.B1(n_429),
.B2(n_435),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_438),
.A2(n_427),
.B1(n_428),
.B2(n_408),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_456),
.C(n_447),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_449),
.A2(n_434),
.B1(n_418),
.B2(n_423),
.Y(n_476)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_407),
.C(n_441),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_411),
.C(n_430),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_479),
.B(n_482),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_448),
.A2(n_434),
.B1(n_426),
.B2(n_413),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_416),
.C(n_344),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_294),
.C(n_6),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_483),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_7),
.C(n_446),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_487),
.B(n_504),
.Y(n_515)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_455),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_496),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_458),
.Y(n_495)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_439),
.Y(n_496)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_471),
.Y(n_499)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_499),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_462),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_503),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_461),
.B1(n_464),
.B2(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_502),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_482),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_481),
.A2(n_443),
.B(n_453),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_492),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_496),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_470),
.C(n_475),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_506),
.A2(n_507),
.B(n_508),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_480),
.C(n_472),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_493),
.A2(n_478),
.B(n_471),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_469),
.C(n_474),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_514),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_489),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_467),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_484),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_502),
.B(n_488),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_522),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_506),
.A2(n_487),
.B(n_490),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_520),
.B(n_529),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_510),
.A2(n_466),
.B(n_497),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_527),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_518),
.A2(n_501),
.B1(n_490),
.B2(n_478),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_526),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_509),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_501),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_516),
.A2(n_476),
.B1(n_498),
.B2(n_504),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_484),
.C(n_512),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_532),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_525),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_527),
.A2(n_511),
.B1(n_507),
.B2(n_491),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_511),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_529),
.B(n_521),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_538),
.A2(n_539),
.B(n_540),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_534),
.B(n_533),
.Y(n_540)
);

OAI21x1_ASAP7_75t_SL g542 ( 
.A1(n_537),
.A2(n_522),
.B(n_530),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_523),
.B(n_528),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_541),
.A2(n_495),
.B(n_519),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_543),
.A2(n_544),
.B(n_484),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_513),
.C(n_486),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_513),
.C(n_483),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_453),
.C(n_7),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_453),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_549),
.B(n_7),
.Y(n_550)
);


endmodule