module fake_aes_6708_n_695 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_695, n_391);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_695;
output n_391;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_16), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_55), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_6), .Y(n_84) );
INVx1_ASAP7_75t_SL g85 ( .A(n_35), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_64), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_66), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_60), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_32), .Y(n_91) );
BUFx5_ASAP7_75t_L g92 ( .A(n_77), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_71), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_14), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_30), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_52), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_18), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_14), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_61), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_13), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_39), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_46), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_2), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_10), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_63), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_20), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_69), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_23), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_58), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_18), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_72), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_3), .Y(n_124) );
NOR2xp67_ASAP7_75t_L g125 ( .A(n_45), .B(n_10), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_0), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_21), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_5), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_8), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_101), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_105), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_118), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_82), .B(n_1), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_89), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_89), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_110), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_107), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_88), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_80), .B(n_1), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_126), .B(n_3), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_92), .B(n_4), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_102), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_82), .B(n_4), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_107), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_119), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_92), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_119), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_97), .B(n_5), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_84), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_92), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_103), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_94), .B(n_6), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_94), .B(n_7), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_108), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_109), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_111), .B(n_7), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_115), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_92), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_116), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_95), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_144), .B(n_111), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_135), .B(n_129), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_163), .B(n_129), .Y(n_181) );
CKINVDCx8_ASAP7_75t_R g182 ( .A(n_142), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_139), .B(n_128), .Y(n_183) );
AO22x2_ASAP7_75t_L g184 ( .A1(n_149), .A2(n_100), .B1(n_124), .B2(n_104), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_136), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_144), .B(n_95), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_139), .B(n_121), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_146), .B(n_127), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_131), .B(n_92), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_167), .B(n_98), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_132), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_146), .B(n_117), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_132), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_132), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_167), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_140), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_131), .B(n_125), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_147), .B(n_123), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_134), .B(n_120), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_138), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_142), .A2(n_112), .B1(n_106), .B2(n_114), .Y(n_218) );
AO22x2_ASAP7_75t_L g219 ( .A1(n_147), .A2(n_122), .B1(n_113), .B2(n_99), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_148), .B(n_106), .Y(n_220) );
AO22x2_ASAP7_75t_L g221 ( .A1(n_148), .A2(n_85), .B1(n_112), .B2(n_12), .Y(n_221) );
INVx1_ASAP7_75t_SL g222 ( .A(n_143), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_150), .B(n_92), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_141), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_132), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_150), .B(n_8), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_159), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_157), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_161), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_138), .Y(n_231) );
INVx5_ASAP7_75t_L g232 ( .A(n_133), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_152), .B(n_43), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_166), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_151), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_145), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_170), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_151), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_151), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_234), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_180), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_217), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_197), .Y(n_245) );
CKINVDCx6p67_ASAP7_75t_R g246 ( .A(n_222), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_234), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_231), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_199), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_175), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_179), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_206), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_194), .A2(n_145), .B(n_164), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_229), .B(n_235), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_229), .B(n_173), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_210), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
AND3x1_ASAP7_75t_SL g262 ( .A(n_181), .B(n_173), .C(n_171), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_207), .A2(n_145), .B(n_164), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_203), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_238), .B(n_156), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_203), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_226), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_208), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_177), .B(n_156), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_210), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_236), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_223), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_178), .B(n_137), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_213), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_177), .B(n_165), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_184), .A2(n_165), .B1(n_171), .B2(n_169), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_215), .B(n_169), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
NOR2xp33_ASAP7_75t_R g282 ( .A(n_182), .B(n_130), .Y(n_282) );
INVx5_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_183), .Y(n_284) );
INVx5_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
INVx5_ASAP7_75t_L g288 ( .A(n_232), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_183), .B(n_152), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_190), .B(n_168), .Y(n_290) );
BUFx10_ASAP7_75t_L g291 ( .A(n_228), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_196), .B(n_155), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_199), .Y(n_293) );
CKINVDCx8_ASAP7_75t_R g294 ( .A(n_209), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_215), .B(n_168), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_188), .B(n_153), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_184), .A2(n_153), .B1(n_154), .B2(n_172), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_185), .Y(n_298) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_190), .B(n_160), .Y(n_299) );
BUFx4f_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_198), .B(n_160), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_198), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_185), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_184), .A2(n_219), .B1(n_195), .B2(n_200), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_230), .B(n_172), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_195), .B(n_160), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_200), .B(n_164), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_227), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_211), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_211), .B(n_9), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_254), .B(n_219), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_267), .B(n_219), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_304), .B(n_212), .C(n_233), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_267), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_260), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_276), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_253), .A2(n_240), .B(n_239), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_276), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_256), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_260), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_263), .A2(n_196), .B(n_186), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_280), .B(n_212), .Y(n_324) );
AO31x2_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_233), .A3(n_193), .B(n_191), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_258), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_279), .A2(n_220), .B1(n_221), .B2(n_218), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
NAND2x2_ASAP7_75t_L g330 ( .A(n_294), .B(n_284), .Y(n_330) );
INVx8_ASAP7_75t_L g331 ( .A(n_310), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_278), .B(n_220), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_284), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_243), .Y(n_336) );
OA22x2_ASAP7_75t_L g337 ( .A1(n_272), .A2(n_225), .B1(n_221), .B2(n_214), .Y(n_337) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_300), .A2(n_221), .B1(n_214), .B2(n_186), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_246), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_295), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_252), .A2(n_255), .B(n_271), .C(n_296), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_306), .A2(n_250), .B(n_251), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_242), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_242), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_176), .B1(n_232), .B2(n_237), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_285), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_246), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_308), .B(n_176), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_258), .Y(n_351) );
INVxp33_ASAP7_75t_L g352 ( .A(n_274), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_244), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_286), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_285), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_285), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_275), .B(n_232), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_250), .A2(n_237), .B(n_192), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_248), .Y(n_359) );
INVxp33_ASAP7_75t_L g360 ( .A(n_282), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_310), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_289), .B(n_9), .Y(n_362) );
BUFx4f_ASAP7_75t_L g363 ( .A(n_310), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_278), .A2(n_193), .B1(n_192), .B2(n_191), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_300), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_354), .B(n_291), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_320), .B(n_251), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_343), .A2(n_307), .B(n_257), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_316), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_338), .A2(n_257), .B1(n_270), .B2(n_258), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_358), .A2(n_270), .B(n_292), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_361), .A2(n_281), .B1(n_248), .B2(n_290), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_328), .A2(n_262), .B1(n_309), .B2(n_301), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_352), .B(n_291), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_313), .A2(n_281), .B(n_299), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_313), .A2(n_292), .B(n_266), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_318), .A2(n_292), .B(n_245), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_315), .B(n_291), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_336), .B(n_247), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_365), .B(n_305), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_314), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_317), .B(n_241), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_361), .A2(n_247), .B1(n_241), .B2(n_264), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_314), .Y(n_384) );
AO21x2_ASAP7_75t_L g385 ( .A1(n_364), .A2(n_265), .B(n_245), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_327), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_322), .A2(n_261), .B1(n_264), .B2(n_288), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_294), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_323), .A2(n_268), .B(n_265), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_331), .Y(n_390) );
UNKNOWN g391 ( );
CKINVDCx11_ASAP7_75t_R g392 ( .A(n_339), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_336), .A2(n_287), .B(n_269), .C(n_268), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_319), .B(n_288), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_363), .B(n_288), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_337), .A2(n_266), .B(n_269), .Y(n_397) );
NOR2xp33_ASAP7_75t_R g398 ( .A(n_349), .B(n_288), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_344), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_396), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_388), .A2(n_363), .B1(n_332), .B2(n_331), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_396), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_370), .A2(n_312), .B1(n_331), .B2(n_311), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_362), .B1(n_347), .B2(n_359), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_392), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_364), .B(n_345), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_400), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_370), .A2(n_339), .B1(n_334), .B2(n_330), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_399), .B(n_324), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_388), .A2(n_353), .B1(n_326), .B2(n_321), .Y(n_411) );
OR2x6_ASAP7_75t_L g412 ( .A(n_400), .B(n_342), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_400), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_346), .B(n_325), .Y(n_414) );
AOI21x1_ASAP7_75t_L g415 ( .A1(n_368), .A2(n_287), .B(n_325), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_398), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_377), .A2(n_325), .B(n_357), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_378), .A2(n_333), .B1(n_335), .B2(n_340), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_367), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_367), .A2(n_355), .B1(n_356), .B2(n_314), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_378), .A2(n_350), .B1(n_355), .B2(n_356), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_298), .B(n_303), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_369), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_375), .A2(n_298), .B(n_303), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_391), .A2(n_350), .B1(n_356), .B2(n_348), .Y(n_428) );
OR2x6_ASAP7_75t_L g429 ( .A(n_372), .B(n_348), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_373), .A2(n_348), .B1(n_329), .B2(n_261), .C(n_283), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_429), .Y(n_431) );
NAND2xp33_ASAP7_75t_R g432 ( .A(n_429), .B(n_381), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_421), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_429), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_429), .Y(n_435) );
OAI211xp5_ASAP7_75t_L g436 ( .A1(n_409), .A2(n_373), .B(n_366), .C(n_374), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_421), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_421), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_413), .B(n_385), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_429), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_413), .B(n_379), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_420), .A2(n_382), .B1(n_379), .B2(n_383), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_415), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_409), .A2(n_387), .B(n_395), .C(n_393), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
NOR2xp33_ASAP7_75t_R g448 ( .A(n_406), .B(n_390), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_420), .B(n_385), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_412), .B(n_385), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_418), .A2(n_397), .B(n_368), .Y(n_451) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_418), .A2(n_397), .B(n_377), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_404), .B(n_385), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_404), .B(n_395), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_417), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_394), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_405), .A2(n_371), .B(n_389), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_407), .Y(n_461) );
BUFx4f_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_405), .A2(n_382), .B1(n_383), .B2(n_390), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_401), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_412), .B(n_394), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_411), .A2(n_401), .B1(n_403), .B2(n_426), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_440), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_440), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_443), .B(n_424), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_440), .B(n_407), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_439), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_448), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_441), .B(n_414), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_436), .A2(n_402), .B1(n_410), .B2(n_419), .C(n_428), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_441), .B(n_414), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_449), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_449), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_433), .B(n_414), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_457), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_464), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_433), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_437), .B(n_418), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_464), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_457), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_443), .B(n_410), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_457), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_443), .B(n_401), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_437), .B(n_403), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_437), .B(n_403), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_462), .A2(n_430), .B1(n_423), .B2(n_416), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_438), .B(n_417), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_462), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_464), .Y(n_496) );
OAI31xp33_ASAP7_75t_L g497 ( .A1(n_436), .A2(n_430), .A3(n_416), .B(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_465), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_465), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_466), .B(n_417), .Y(n_500) );
OAI33xp33_ASAP7_75t_L g501 ( .A1(n_463), .A2(n_12), .A3(n_13), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_438), .B(n_417), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_462), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_466), .A2(n_463), .B1(n_444), .B2(n_454), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
OAI33xp33_ASAP7_75t_L g506 ( .A1(n_444), .A2(n_15), .A3(n_17), .B1(n_19), .B2(n_394), .B3(n_386), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_442), .B(n_397), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_448), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_442), .B(n_384), .Y(n_509) );
INVxp67_ASAP7_75t_SL g510 ( .A(n_438), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_445), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_458), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_446), .A2(n_371), .B(n_380), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_450), .B(n_384), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_445), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_435), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_473), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_469), .B(n_454), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_511), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_501), .A2(n_460), .B1(n_458), .B2(n_455), .C(n_459), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_472), .Y(n_521) );
OR2x6_ASAP7_75t_L g522 ( .A(n_476), .B(n_435), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_508), .B(n_446), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_486), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_483), .B(n_462), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_490), .B(n_454), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_486), .Y(n_527) );
NAND2xp33_ASAP7_75t_SL g528 ( .A(n_476), .B(n_435), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_474), .B(n_450), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_488), .B(n_455), .Y(n_530) );
OAI332xp33_ASAP7_75t_L g531 ( .A1(n_472), .A2(n_453), .A3(n_460), .B1(n_461), .B2(n_434), .B3(n_447), .C1(n_445), .C2(n_19), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_477), .B(n_450), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_467), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_503), .B(n_442), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_486), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_513), .A2(n_459), .B(n_380), .Y(n_536) );
NAND2x1_ASAP7_75t_L g537 ( .A(n_503), .B(n_434), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_511), .Y(n_538) );
NAND4xp25_ASAP7_75t_L g539 ( .A(n_504), .B(n_453), .C(n_442), .D(n_432), .Y(n_539) );
NAND2x1_ASAP7_75t_L g540 ( .A(n_495), .B(n_434), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_491), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_515), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_514), .B(n_431), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_474), .B(n_453), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_478), .B(n_482), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_506), .B(n_456), .C(n_380), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_515), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_477), .B(n_461), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g549 ( .A(n_497), .B(n_431), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_475), .A2(n_432), .B1(n_456), .B2(n_461), .C(n_447), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_468), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_478), .B(n_452), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_504), .A2(n_380), .B1(n_456), .B2(n_381), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_482), .B(n_456), .Y(n_554) );
OAI211xp5_ASAP7_75t_SL g555 ( .A1(n_493), .A2(n_456), .B(n_447), .C(n_381), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_468), .Y(n_556) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_510), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_487), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_487), .B(n_451), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_489), .B(n_452), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_489), .B(n_451), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_498), .B(n_452), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_498), .B(n_452), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_499), .B(n_452), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_512), .B(n_201), .C(n_202), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_505), .B(n_452), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_471), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_492), .B(n_451), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_492), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_514), .B(n_451), .Y(n_570) );
AOI332xp33_ASAP7_75t_L g571 ( .A1(n_558), .A2(n_479), .A3(n_480), .B1(n_470), .B2(n_500), .B3(n_481), .C1(n_495), .C2(n_485), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_549), .A2(n_495), .B1(n_480), .B2(n_479), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_553), .A2(n_495), .B1(n_496), .B2(n_483), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_521), .Y(n_574) );
OAI321xp33_ASAP7_75t_L g575 ( .A1(n_539), .A2(n_470), .A3(n_485), .B1(n_481), .B2(n_494), .C(n_502), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_569), .Y(n_576) );
OAI22xp33_ASAP7_75t_SL g577 ( .A1(n_524), .A2(n_496), .B1(n_516), .B2(n_494), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g578 ( .A1(n_523), .A2(n_507), .B(n_496), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_517), .B(n_509), .Y(n_579) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_550), .A2(n_509), .B(n_451), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_546), .A2(n_502), .B1(n_484), .B2(n_471), .C(n_384), .Y(n_581) );
AOI32xp33_ASAP7_75t_L g582 ( .A1(n_528), .A2(n_507), .A3(n_509), .B1(n_484), .B2(n_384), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_536), .A2(n_427), .B1(n_425), .B2(n_202), .C(n_201), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_531), .B(n_509), .C(n_427), .Y(n_584) );
OAI21xp33_ASAP7_75t_SL g585 ( .A1(n_525), .A2(n_535), .B(n_522), .Y(n_585) );
OAI32xp33_ASAP7_75t_L g586 ( .A1(n_528), .A2(n_386), .A3(n_425), .B1(n_507), .B2(n_26), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_545), .B(n_507), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_524), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_529), .B(n_22), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_529), .B(n_24), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_530), .B(n_25), .Y(n_592) );
OAI222xp33_ASAP7_75t_L g593 ( .A1(n_522), .A2(n_389), .B1(n_283), .B2(n_273), .C1(n_288), .C2(n_40), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_557), .A2(n_329), .B1(n_283), .B2(n_273), .Y(n_594) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_519), .Y(n_595) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_525), .A2(n_27), .B(n_28), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_530), .A2(n_201), .B1(n_202), .B2(n_187), .C(n_189), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_522), .A2(n_329), .B1(n_283), .B2(n_273), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g599 ( .A(n_518), .B(n_37), .C(n_38), .D(n_42), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_526), .A2(n_201), .B1(n_189), .B2(n_187), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_552), .A2(n_570), .B(n_544), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_533), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_527), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_522), .A2(n_283), .B1(n_273), .B2(n_189), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_520), .A2(n_189), .B1(n_187), .B2(n_273), .C(n_259), .Y(n_605) );
AOI21xp33_ASAP7_75t_L g606 ( .A1(n_555), .A2(n_44), .B(n_47), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_559), .A2(n_48), .B(n_49), .C(n_50), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_551), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_534), .A2(n_187), .B1(n_277), .B2(n_259), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_570), .A2(n_293), .B1(n_277), .B2(n_259), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_535), .B(n_293), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_537), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g613 ( .A1(n_552), .A2(n_293), .B(n_277), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_532), .B(n_53), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_567), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_543), .B(n_54), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_544), .B(n_56), .Y(n_617) );
NOR2xp33_ASAP7_75t_SL g618 ( .A(n_585), .B(n_534), .Y(n_618) );
XNOR2xp5_ASAP7_75t_L g619 ( .A(n_588), .B(n_534), .Y(n_619) );
AOI211xp5_ASAP7_75t_SL g620 ( .A1(n_575), .A2(n_568), .B(n_561), .C(n_554), .Y(n_620) );
NAND2xp33_ASAP7_75t_SL g621 ( .A(n_589), .B(n_540), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_603), .B(n_562), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_576), .B(n_562), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_592), .A2(n_548), .B(n_534), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_571), .A2(n_556), .B(n_565), .C(n_566), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_586), .A2(n_567), .B(n_519), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_591), .B(n_566), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_602), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_611), .B(n_547), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_608), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_577), .B(n_547), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_587), .B(n_564), .Y(n_633) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_579), .B(n_564), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_601), .B(n_563), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_595), .B(n_563), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_615), .Y(n_637) );
NOR3xp33_ASAP7_75t_SL g638 ( .A(n_599), .B(n_57), .C(n_59), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_584), .B(n_560), .Y(n_639) );
INVxp33_ASAP7_75t_SL g640 ( .A(n_590), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_612), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_617), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_572), .B(n_542), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_573), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_593), .A2(n_538), .B(n_542), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_573), .Y(n_648) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_639), .B(n_580), .C(n_616), .D(n_606), .Y(n_649) );
NOR4xp75_ASAP7_75t_L g650 ( .A(n_632), .B(n_578), .C(n_605), .D(n_598), .Y(n_650) );
AOI21xp5_ASAP7_75t_SL g651 ( .A1(n_632), .A2(n_598), .B(n_604), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_618), .B(n_582), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_636), .B(n_538), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_641), .A2(n_580), .B1(n_594), .B2(n_604), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_645), .B(n_613), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_640), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_648), .B(n_594), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_620), .A2(n_583), .B1(n_606), .B2(n_596), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_621), .A2(n_607), .B(n_597), .C(n_609), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_635), .B(n_600), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_635), .A2(n_610), .B1(n_293), .B2(n_277), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_642), .B(n_68), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_619), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_622), .Y(n_664) );
AOI221x1_ASAP7_75t_L g665 ( .A1(n_621), .A2(n_293), .B1(n_277), .B2(n_259), .C(n_249), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_637), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_657), .B(n_641), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_651), .A2(n_633), .B1(n_626), .B2(n_628), .Y(n_668) );
AOI22x1_ASAP7_75t_L g669 ( .A1(n_656), .A2(n_646), .B1(n_630), .B2(n_627), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_655), .B(n_626), .Y(n_670) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_651), .B(n_629), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_660), .B(n_631), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_652), .A2(n_634), .B1(n_623), .B2(n_647), .Y(n_673) );
NOR2xp33_ASAP7_75t_R g674 ( .A(n_663), .B(n_643), .Y(n_674) );
NOR3xp33_ASAP7_75t_SL g675 ( .A(n_658), .B(n_649), .C(n_662), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_654), .B(n_644), .Y(n_676) );
OAI22xp33_ASAP7_75t_SL g677 ( .A1(n_664), .A2(n_630), .B1(n_638), .B2(n_625), .Y(n_677) );
XOR2xp5_ASAP7_75t_L g678 ( .A(n_658), .B(n_624), .Y(n_678) );
OAI321xp33_ASAP7_75t_L g679 ( .A1(n_659), .A2(n_638), .A3(n_74), .B1(n_76), .B2(n_78), .C(n_70), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_653), .A2(n_249), .A3(n_651), .B1(n_639), .B2(n_652), .C1(n_663), .C2(n_657), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_650), .B(n_661), .C(n_665), .Y(n_681) );
NOR4xp75_ASAP7_75t_L g682 ( .A(n_666), .B(n_652), .C(n_649), .D(n_639), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_674), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_680), .B(n_681), .C(n_671), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_675), .Y(n_685) );
NOR3xp33_ASAP7_75t_SL g686 ( .A(n_668), .B(n_679), .C(n_670), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_676), .B(n_667), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_687), .B(n_672), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_685), .B(n_683), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_684), .A2(n_675), .B1(n_678), .B2(n_673), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_688), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g692 ( .A(n_690), .B(n_682), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_691), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_692), .B1(n_689), .B2(n_686), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_677), .B(n_669), .Y(n_695) );
endmodule