module fake_jpeg_23673_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_40),
.B(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_24),
.B1(n_26),
.B2(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_32),
.B(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_38),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_65),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_29),
.B(n_30),
.C(n_34),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_36),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_80),
.B1(n_41),
.B2(n_35),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_30),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_86),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_50),
.C(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_95),
.B1(n_102),
.B2(n_58),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_19),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_100),
.Y(n_118)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_96),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_39),
.B1(n_34),
.B2(n_35),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_0),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_39),
.B1(n_41),
.B2(n_45),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_42),
.C(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_78),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_65),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_115),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_66),
.CON(n_110),
.SN(n_110)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_110),
.A2(n_126),
.B(n_74),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_58),
.B1(n_41),
.B2(n_82),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_111),
.C(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_65),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_125),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_67),
.B(n_80),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_62),
.B(n_47),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_99),
.B1(n_58),
.B2(n_45),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_89),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_151),
.C(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_124),
.B1(n_107),
.B2(n_57),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_145),
.B(n_149),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_120),
.B(n_114),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_109),
.B(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_61),
.C(n_77),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_155),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_118),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_169),
.C(n_178),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_159),
.B(n_160),
.Y(n_190)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_106),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_44),
.A3(n_48),
.B1(n_51),
.B2(n_33),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_126),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_165),
.B1(n_167),
.B2(n_24),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_134),
.B1(n_146),
.B2(n_136),
.Y(n_184)
);

OAI22x1_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_130),
.B1(n_117),
.B2(n_122),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_125),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_105),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_179),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_116),
.C(n_61),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_182),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_113),
.B1(n_57),
.B2(n_47),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_183),
.B1(n_132),
.B2(n_131),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_187),
.B1(n_189),
.B2(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_135),
.B1(n_141),
.B2(n_150),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_186),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_146),
.B1(n_150),
.B2(n_138),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_149),
.B1(n_141),
.B2(n_152),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_143),
.B(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_151),
.B1(n_137),
.B2(n_113),
.Y(n_194)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_137),
.C(n_116),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_178),
.C(n_168),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_208),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

XOR2x1_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_14),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_54),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_86),
.B(n_83),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_207),
.B1(n_176),
.B2(n_173),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_69),
.B1(n_24),
.B2(n_19),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_158),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_215),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_176),
.B1(n_164),
.B2(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_26),
.B1(n_14),
.B2(n_27),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_168),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_226),
.C(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_202),
.B1(n_200),
.B2(n_188),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_72),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_230),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_225),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_167),
.C(n_48),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_1),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_231),
.A2(n_236),
.B1(n_238),
.B2(n_21),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_187),
.B1(n_209),
.B2(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_240),
.C(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_228),
.B1(n_222),
.B2(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_194),
.B1(n_184),
.B2(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_201),
.C(n_97),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_201),
.C(n_69),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_76),
.B1(n_14),
.B2(n_26),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_76),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_51),
.C(n_44),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_248),
.B(n_227),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_52),
.C(n_54),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_214),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_211),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_261),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_241),
.B(n_20),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_211),
.C(n_13),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_264),
.C(n_267),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_250),
.B1(n_242),
.B2(n_246),
.Y(n_270)
);

NAND4xp25_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_52),
.C(n_33),
.D(n_37),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_17),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_25),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_236),
.B(n_11),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_33),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_37),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_238),
.B(n_249),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_274),
.B(n_275),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_276),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_281),
.B1(n_37),
.B2(n_2),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_240),
.B1(n_239),
.B2(n_233),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_273),
.A2(n_20),
.B1(n_16),
.B2(n_3),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_254),
.B(n_252),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_18),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_269),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_52),
.C(n_25),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_7),
.C(n_12),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_282),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_263),
.B(n_21),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_272),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_290),
.C(n_289),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_7),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_16),
.C(n_2),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_8),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_293),
.B(n_277),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_296),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_300),
.Y(n_308)
);

AOI211xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_6),
.B(n_12),
.C(n_11),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_10),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_6),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_290),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_286),
.A3(n_10),
.B1(n_4),
.B2(n_5),
.C1(n_3),
.C2(n_1),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_3),
.C(n_4),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_296),
.B(n_4),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_3),
.B(n_4),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_311),
.B(n_305),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_5),
.B(n_37),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule