module real_aes_16575_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1730;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_1749;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_1343;
wire n_465;
wire n_719;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_0), .A2(n_93), .B1(n_1001), .B2(n_1254), .C(n_1274), .Y(n_1273) );
AOI22xp33_ASAP7_75t_SL g1293 ( .A1(n_0), .A2(n_198), .B1(n_1294), .B2(n_1296), .Y(n_1293) );
INVx1_ASAP7_75t_L g884 ( .A(n_1), .Y(n_884) );
INVx1_ASAP7_75t_L g327 ( .A(n_2), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_2), .B(n_337), .Y(n_412) );
AND2x2_ASAP7_75t_L g598 ( .A(n_2), .B(n_211), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_2), .B(n_516), .Y(n_616) );
INVx1_ASAP7_75t_L g1222 ( .A(n_3), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1242 ( .A1(n_3), .A2(n_9), .B1(n_627), .B2(n_989), .Y(n_1242) );
INVx1_ASAP7_75t_L g1418 ( .A(n_4), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_4), .A2(n_73), .B1(n_942), .B2(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1178 ( .A(n_5), .Y(n_1178) );
INVx1_ASAP7_75t_L g1263 ( .A(n_6), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1300 ( .A1(n_6), .A2(n_80), .B1(n_909), .B2(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1407 ( .A(n_7), .Y(n_1407) );
INVx1_ASAP7_75t_L g693 ( .A(n_8), .Y(n_693) );
OA222x2_ASAP7_75t_L g717 ( .A1(n_8), .A2(n_120), .B1(n_144), .B2(n_718), .C1(n_720), .C2(n_726), .Y(n_717) );
INVx1_ASAP7_75t_L g1232 ( .A(n_9), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_10), .A2(n_285), .B1(n_753), .B2(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1689 ( .A(n_10), .Y(n_1689) );
OAI221xp5_ASAP7_75t_L g1311 ( .A1(n_11), .A2(n_302), .B1(n_695), .B2(n_942), .C(n_943), .Y(n_1311) );
OAI21xp33_ASAP7_75t_SL g1340 ( .A1(n_11), .A2(n_726), .B(n_754), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_12), .A2(n_79), .B1(n_878), .B2(n_1123), .C(n_1254), .Y(n_1253) );
AOI22xp33_ASAP7_75t_SL g1299 ( .A1(n_12), .A2(n_166), .B1(n_778), .B2(n_1292), .Y(n_1299) );
INVx2_ASAP7_75t_L g366 ( .A(n_13), .Y(n_366) );
INVx1_ASAP7_75t_L g883 ( .A(n_14), .Y(n_883) );
OAI322xp33_ASAP7_75t_L g887 ( .A1(n_14), .A2(n_538), .A3(n_888), .B1(n_893), .B2(n_894), .C1(n_897), .C2(n_903), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_15), .A2(n_18), .B1(n_1457), .B2(n_1464), .Y(n_1473) );
CKINVDCx5p33_ASAP7_75t_R g1737 ( .A(n_16), .Y(n_1737) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_17), .A2(n_148), .B1(n_673), .B2(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_17), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_19), .A2(n_196), .B1(n_736), .B2(n_875), .C(n_878), .Y(n_874) );
INVx1_ASAP7_75t_L g896 ( .A(n_19), .Y(n_896) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_20), .A2(n_247), .B1(n_920), .B2(n_923), .Y(n_1322) );
INVx1_ASAP7_75t_L g1339 ( .A(n_20), .Y(n_1339) );
INVx1_ASAP7_75t_L g985 ( .A(n_21), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_22), .A2(n_273), .B1(n_920), .B2(n_923), .Y(n_1179) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_22), .Y(n_1181) );
INVx1_ASAP7_75t_L g1376 ( .A(n_23), .Y(n_1376) );
AOI221xp5_ASAP7_75t_L g1391 ( .A1(n_23), .A2(n_118), .B1(n_926), .B2(n_1392), .C(n_1394), .Y(n_1391) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_24), .Y(n_322) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_24), .B(n_320), .Y(n_1458) );
OA22x2_ASAP7_75t_L g344 ( .A1(n_25), .A2(n_345), .B1(n_529), .B2(n_530), .Y(n_344) );
INVxp67_ASAP7_75t_L g530 ( .A(n_25), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_26), .A2(n_156), .B1(n_1457), .B2(n_1513), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_27), .A2(n_188), .B1(n_684), .B2(n_791), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_27), .A2(n_257), .B1(n_753), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_28), .A2(n_256), .B1(n_862), .B2(n_880), .Y(n_879) );
INVxp67_ASAP7_75t_L g891 ( .A(n_28), .Y(n_891) );
INVx1_ASAP7_75t_L g414 ( .A(n_29), .Y(n_414) );
INVx1_ASAP7_75t_L g1099 ( .A(n_30), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_30), .A2(n_56), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx1_ASAP7_75t_L g848 ( .A(n_31), .Y(n_848) );
OAI211xp5_ASAP7_75t_SL g981 ( .A1(n_32), .A2(n_982), .B(n_984), .C(n_987), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_32), .A2(n_232), .B1(n_607), .B2(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1171 ( .A(n_33), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_34), .A2(n_254), .B1(n_862), .B2(n_863), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_34), .A2(n_196), .B1(n_676), .B2(n_778), .Y(n_902) );
INVx1_ASAP7_75t_L g1382 ( .A(n_35), .Y(n_1382) );
OAI22xp33_ASAP7_75t_L g1389 ( .A1(n_35), .A2(n_43), .B1(n_942), .B2(n_943), .Y(n_1389) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_36), .A2(n_230), .B1(n_670), .B2(n_673), .Y(n_669) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_36), .Y(n_738) );
INVx1_ASAP7_75t_L g1678 ( .A(n_37), .Y(n_1678) );
INVx1_ASAP7_75t_L g938 ( .A(n_38), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g1724 ( .A1(n_39), .A2(n_940), .B1(n_1725), .B2(n_1728), .Y(n_1724) );
INVx1_ASAP7_75t_L g1742 ( .A(n_39), .Y(n_1742) );
INVx1_ASAP7_75t_L g935 ( .A(n_40), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_40), .A2(n_225), .B1(n_646), .B2(n_966), .C(n_967), .Y(n_965) );
INVx1_ASAP7_75t_L g1677 ( .A(n_41), .Y(n_1677) );
OAI221xp5_ASAP7_75t_L g994 ( .A1(n_42), .A2(n_102), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_994) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_42), .A2(n_102), .B1(n_1024), .B2(n_1026), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g1378 ( .A1(n_43), .A2(n_263), .B1(n_754), .B2(n_1148), .C(n_1202), .Y(n_1378) );
INVx1_ASAP7_75t_L g1157 ( .A(n_44), .Y(n_1157) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_45), .A2(n_215), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_45), .A2(n_304), .B1(n_561), .B2(n_778), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g1511 ( .A1(n_46), .A2(n_171), .B1(n_1464), .B2(n_1467), .Y(n_1511) );
AOI22xp5_ASAP7_75t_L g1482 ( .A1(n_47), .A2(n_291), .B1(n_1457), .B2(n_1461), .Y(n_1482) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_48), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_49), .A2(n_288), .B1(n_683), .B2(n_686), .C(n_1114), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_49), .A2(n_141), .B1(n_1121), .B2(n_1123), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g1164 ( .A1(n_50), .A2(n_686), .B(n_778), .Y(n_1164) );
INVxp67_ASAP7_75t_SL g1190 ( .A(n_50), .Y(n_1190) );
INVx1_ASAP7_75t_L g1221 ( .A(n_51), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_51), .A2(n_152), .B1(n_627), .B2(n_966), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_52), .A2(n_164), .B1(n_794), .B2(n_940), .Y(n_1095) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_52), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1371 ( .A(n_53), .Y(n_1371) );
AOI22xp5_ASAP7_75t_L g1512 ( .A1(n_54), .A2(n_268), .B1(n_1457), .B2(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1731 ( .A(n_55), .Y(n_1731) );
AOI22xp33_ASAP7_75t_L g1750 ( .A1(n_55), .A2(n_58), .B1(n_655), .B2(n_752), .Y(n_1750) );
INVx1_ASAP7_75t_L g1117 ( .A(n_56), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1463 ( .A1(n_57), .A2(n_109), .B1(n_1464), .B2(n_1467), .Y(n_1463) );
AOI221xp5_ASAP7_75t_L g1719 ( .A1(n_58), .A2(n_297), .B1(n_685), .B2(n_1297), .C(n_1720), .Y(n_1719) );
INVxp67_ASAP7_75t_SL g1380 ( .A(n_59), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_59), .A2(n_940), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
OAI221xp5_ASAP7_75t_L g1158 ( .A1(n_60), .A2(n_212), .B1(n_695), .B2(n_942), .C(n_943), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_60), .A2(n_273), .B1(n_754), .B2(n_1148), .C(n_1202), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_61), .A2(n_244), .B1(n_794), .B2(n_940), .Y(n_939) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_61), .Y(n_946) );
AOI21xp33_ASAP7_75t_L g1323 ( .A1(n_62), .A2(n_1324), .B(n_1327), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_62), .A2(n_94), .B1(n_1254), .B2(n_1351), .C(n_1352), .Y(n_1350) );
INVx1_ASAP7_75t_L g768 ( .A(n_63), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g1712 ( .A1(n_64), .A2(n_1713), .B1(n_1714), .B2(n_1715), .Y(n_1712) );
CKINVDCx5p33_ASAP7_75t_R g1713 ( .A(n_64), .Y(n_1713) );
INVx1_ASAP7_75t_L g1100 ( .A(n_65), .Y(n_1100) );
OAI21xp33_ASAP7_75t_L g1145 ( .A1(n_65), .A2(n_726), .B(n_754), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_66), .Y(n_907) );
INVx1_ASAP7_75t_L g870 ( .A(n_67), .Y(n_870) );
OAI211xp5_ASAP7_75t_L g908 ( .A1(n_67), .A2(n_909), .B(n_910), .C(n_913), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_68), .Y(n_779) );
INVx1_ASAP7_75t_L g1384 ( .A(n_69), .Y(n_1384) );
OAI222xp33_ASAP7_75t_L g1387 ( .A1(n_69), .A2(n_252), .B1(n_263), .B2(n_478), .C1(n_489), .C2(n_1048), .Y(n_1387) );
AOI21xp33_ASAP7_75t_L g1000 ( .A1(n_70), .A2(n_627), .B(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1010 ( .A(n_70), .Y(n_1010) );
XOR2x2_ASAP7_75t_L g1306 ( .A(n_71), .B(n_1307), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_72), .A2(n_270), .B1(n_580), .B2(n_584), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_72), .A2(n_294), .B1(n_625), .B2(n_627), .C(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g1412 ( .A(n_73), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_74), .A2(n_153), .B1(n_398), .B2(n_400), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_74), .A2(n_153), .B1(n_512), .B2(n_517), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_75), .A2(n_303), .B1(n_1464), .B2(n_1467), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_76), .Y(n_1105) );
INVx1_ASAP7_75t_L g453 ( .A(n_77), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_78), .A2(n_169), .B1(n_603), .B2(n_607), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_79), .A2(n_231), .B1(n_1291), .B2(n_1292), .Y(n_1290) );
INVx1_ASAP7_75t_L g1261 ( .A(n_80), .Y(n_1261) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_81), .A2(n_280), .B1(n_926), .B2(n_1054), .C(n_1056), .Y(n_1053) );
INVx1_ASAP7_75t_L g1086 ( .A(n_81), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_82), .A2(n_178), .B1(n_794), .B2(n_940), .Y(n_1312) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_82), .Y(n_1349) );
AOI22xp5_ASAP7_75t_SL g1490 ( .A1(n_83), .A2(n_182), .B1(n_1457), .B2(n_1461), .Y(n_1490) );
XNOR2xp5_ASAP7_75t_L g1665 ( .A(n_83), .B(n_1666), .Y(n_1665) );
AOI22xp33_ASAP7_75t_L g1707 ( .A1(n_83), .A2(n_1708), .B1(n_1711), .B2(n_1752), .Y(n_1707) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_84), .A2(n_100), .B1(n_683), .B2(n_684), .C(n_686), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_84), .A2(n_230), .B1(n_752), .B2(n_753), .Y(n_751) );
AOI222xp33_ASAP7_75t_L g1328 ( .A1(n_85), .A2(n_122), .B1(n_292), .B2(n_488), .C1(n_543), .C2(n_674), .Y(n_1328) );
INVx1_ASAP7_75t_L g1353 ( .A(n_85), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_86), .Y(n_1372) );
INVx1_ASAP7_75t_L g929 ( .A(n_87), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g958 ( .A1(n_87), .A2(n_163), .B1(n_959), .B2(n_960), .C(n_962), .Y(n_958) );
AOI21xp33_ASAP7_75t_L g1682 ( .A1(n_88), .A2(n_646), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1688 ( .A(n_88), .Y(n_1688) );
OAI22xp33_ASAP7_75t_L g1738 ( .A1(n_89), .A2(n_121), .B1(n_942), .B2(n_943), .Y(n_1738) );
OAI22xp5_ASAP7_75t_L g1751 ( .A1(n_89), .A2(n_250), .B1(n_1148), .B2(n_1202), .Y(n_1751) );
INVx1_ASAP7_75t_L g456 ( .A(n_90), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g1377 ( .A(n_91), .Y(n_1377) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_92), .A2(n_193), .B1(n_545), .B2(n_553), .C(n_559), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_92), .A2(n_612), .B(n_617), .C(n_630), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_93), .A2(n_235), .B1(n_788), .B2(n_791), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1314 ( .A1(n_94), .A2(n_187), .B1(n_1315), .B2(n_1317), .C(n_1319), .Y(n_1314) );
INVx1_ASAP7_75t_L g320 ( .A(n_95), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g1671 ( .A1(n_96), .A2(n_213), .B1(n_629), .B2(n_989), .C(n_1672), .Y(n_1671) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_96), .A2(n_145), .B1(n_561), .B2(n_778), .Y(n_1690) );
INVx1_ASAP7_75t_L g1727 ( .A(n_97), .Y(n_1727) );
AOI22xp33_ASAP7_75t_L g1747 ( .A1(n_97), .A2(n_297), .B1(n_724), .B2(n_752), .Y(n_1747) );
INVx1_ASAP7_75t_L g1381 ( .A(n_98), .Y(n_1381) );
INVx1_ASAP7_75t_L g1310 ( .A(n_99), .Y(n_1310) );
OAI21xp33_ASAP7_75t_L g1335 ( .A1(n_99), .A2(n_1336), .B(n_1337), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_100), .A2(n_129), .B1(n_734), .B2(n_736), .C(n_737), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_101), .A2(n_222), .B1(n_603), .B2(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g1230 ( .A(n_103), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_103), .A2(n_132), .B1(n_724), .B2(n_752), .Y(n_1243) );
XOR2x2_ASAP7_75t_L g1036 ( .A(n_104), .B(n_1037), .Y(n_1036) );
AOI22xp5_ASAP7_75t_L g1486 ( .A1(n_104), .A2(n_276), .B1(n_1461), .B2(n_1467), .Y(n_1486) );
CKINVDCx5p33_ASAP7_75t_R g1218 ( .A(n_105), .Y(n_1218) );
INVx1_ASAP7_75t_L g1051 ( .A(n_106), .Y(n_1051) );
INVx1_ASAP7_75t_L g1058 ( .A(n_107), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_108), .A2(n_201), .B1(n_753), .B2(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1013 ( .A(n_108), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1211 ( .A1(n_110), .A2(n_243), .B1(n_794), .B2(n_940), .C(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1246 ( .A(n_110), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_111), .A2(n_765), .B1(n_766), .B2(n_843), .Y(n_764) );
INVx1_ASAP7_75t_L g843 ( .A(n_111), .Y(n_843) );
INVx1_ASAP7_75t_L g1057 ( .A(n_112), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g1722 ( .A(n_113), .Y(n_1722) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_114), .A2(n_167), .B1(n_920), .B2(n_923), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_114), .A2(n_239), .B1(n_604), .B2(n_759), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g1416 ( .A1(n_115), .A2(n_217), .B1(n_753), .B2(n_1257), .Y(n_1416) );
AOI221xp5_ASAP7_75t_L g1434 ( .A1(n_115), .A2(n_290), .B1(n_683), .B2(n_686), .C(n_778), .Y(n_1434) );
INVx1_ASAP7_75t_L g867 ( .A(n_116), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_117), .A2(n_184), .B1(n_794), .B2(n_940), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_117), .Y(n_1065) );
INVx1_ASAP7_75t_L g1363 ( .A(n_118), .Y(n_1363) );
INVx1_ASAP7_75t_L g569 ( .A(n_119), .Y(n_569) );
INVx1_ASAP7_75t_L g710 ( .A(n_120), .Y(n_710) );
INVx1_ASAP7_75t_L g1743 ( .A(n_121), .Y(n_1743) );
INVx1_ASAP7_75t_L g1347 ( .A(n_122), .Y(n_1347) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_123), .A2(n_176), .B1(n_856), .B2(n_857), .C(n_860), .Y(n_855) );
INVxp67_ASAP7_75t_L g889 ( .A(n_123), .Y(n_889) );
OAI221xp5_ASAP7_75t_L g1679 ( .A1(n_124), .A2(n_299), .B1(n_995), .B2(n_996), .C(n_1680), .Y(n_1679) );
OAI22xp33_ASAP7_75t_L g1695 ( .A1(n_124), .A2(n_299), .B1(n_912), .B2(n_1026), .Y(n_1695) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_125), .A2(n_304), .B1(n_989), .B2(n_990), .C(n_991), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_125), .A2(n_215), .B1(n_778), .B2(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1106 ( .A(n_126), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g1126 ( .A1(n_126), .A2(n_135), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_127), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_127), .A2(n_214), .B1(n_625), .B2(n_646), .C(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g1214 ( .A(n_128), .Y(n_1214) );
OAI22xp5_ASAP7_75t_L g1240 ( .A1(n_128), .A2(n_284), .B1(n_604), .B2(n_759), .Y(n_1240) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_129), .A2(n_154), .B1(n_676), .B2(n_677), .C(n_678), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_130), .A2(n_163), .B1(n_926), .B2(n_932), .C(n_934), .Y(n_931) );
INVx1_ASAP7_75t_L g969 ( .A(n_130), .Y(n_969) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_131), .Y(n_773) );
OAI221xp5_ASAP7_75t_L g793 ( .A1(n_131), .A2(n_695), .B1(n_794), .B2(n_796), .C(n_804), .Y(n_793) );
INVx1_ASAP7_75t_L g1224 ( .A(n_132), .Y(n_1224) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_133), .A2(n_678), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g822 ( .A(n_133), .Y(n_822) );
INVx1_ASAP7_75t_L g803 ( .A(n_134), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_134), .A2(n_188), .B1(n_825), .B2(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g1112 ( .A(n_135), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_136), .A2(n_306), .B1(n_674), .B2(n_685), .Y(n_1174) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_136), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_137), .A2(n_239), .B1(n_695), .B2(n_942), .C(n_943), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_137), .Y(n_1063) );
INVx1_ASAP7_75t_L g601 ( .A(n_138), .Y(n_601) );
INVx1_ASAP7_75t_L g1733 ( .A(n_139), .Y(n_1733) );
INVx1_ASAP7_75t_L g1161 ( .A(n_140), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_141), .A2(n_261), .B1(n_678), .B2(n_1054), .C(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1523 ( .A(n_142), .Y(n_1523) );
AOI22xp5_ASAP7_75t_SL g1456 ( .A1(n_143), .A2(n_149), .B1(n_1457), .B2(n_1461), .Y(n_1456) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_144), .A2(n_147), .B1(n_577), .B2(n_703), .C(n_706), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g1684 ( .A1(n_145), .A2(n_267), .B1(n_655), .B2(n_993), .Y(n_1684) );
OAI211xp5_ASAP7_75t_L g1668 ( .A1(n_146), .A2(n_1669), .B(n_1670), .C(n_1676), .Y(n_1668) );
OAI22xp5_ASAP7_75t_L g1698 ( .A1(n_146), .A2(n_293), .B1(n_770), .B2(n_1031), .Y(n_1698) );
INVxp67_ASAP7_75t_SL g728 ( .A(n_147), .Y(n_728) );
INVxp33_ASAP7_75t_SL g739 ( .A(n_148), .Y(n_739) );
INVx2_ASAP7_75t_L g1460 ( .A(n_150), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_150), .B(n_258), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_150), .B(n_1466), .Y(n_1468) );
XNOR2xp5_ASAP7_75t_L g978 ( .A(n_151), .B(n_979), .Y(n_978) );
AOI22xp5_ASAP7_75t_SL g1471 ( .A1(n_151), .A2(n_216), .B1(n_1467), .B2(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1229 ( .A(n_152), .Y(n_1229) );
INVx1_ASAP7_75t_L g747 ( .A(n_154), .Y(n_747) );
INVx1_ASAP7_75t_L g1247 ( .A(n_155), .Y(n_1247) );
OAI21xp33_ASAP7_75t_L g1409 ( .A1(n_157), .A2(n_718), .B(n_1410), .Y(n_1409) );
OAI221xp5_ASAP7_75t_L g1438 ( .A1(n_157), .A2(n_242), .B1(n_807), .B2(n_1439), .C(n_1440), .Y(n_1438) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_158), .A2(n_271), .B1(n_1457), .B2(n_1472), .Y(n_1478) );
AOI22xp5_ASAP7_75t_L g1481 ( .A1(n_159), .A2(n_220), .B1(n_1464), .B2(n_1467), .Y(n_1481) );
INVx1_ASAP7_75t_L g1169 ( .A(n_160), .Y(n_1169) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_161), .A2(n_236), .B1(n_695), .B2(n_942), .C(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g976 ( .A(n_161), .Y(n_976) );
OAI21xp5_ASAP7_75t_SL g1093 ( .A1(n_162), .A2(n_713), .B(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1116 ( .A(n_162), .Y(n_1116) );
INVx1_ASAP7_75t_L g1139 ( .A(n_164), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1487 ( .A1(n_165), .A2(n_237), .B1(n_1457), .B2(n_1464), .Y(n_1487) );
INVxp67_ASAP7_75t_SL g1272 ( .A(n_166), .Y(n_1272) );
OAI211xp5_ASAP7_75t_L g1060 ( .A1(n_167), .A2(n_713), .B(n_1061), .C(n_1064), .Y(n_1060) );
INVx1_ASAP7_75t_L g708 ( .A(n_168), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_168), .A2(n_199), .B1(n_604), .B2(n_759), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g1251 ( .A1(n_169), .A2(n_653), .B(n_1252), .C(n_1260), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_170), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g1681 ( .A(n_172), .Y(n_1681) );
AOI22xp33_ASAP7_75t_SL g1415 ( .A1(n_173), .A2(n_274), .B1(n_877), .B2(n_966), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g1431 ( .A1(n_173), .A2(n_194), .B1(n_678), .B2(n_683), .C(n_1432), .Y(n_1431) );
INVx2_ASAP7_75t_L g350 ( .A(n_174), .Y(n_350) );
INVx1_ASAP7_75t_L g485 ( .A(n_174), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_174), .B(n_366), .Y(n_542) );
INVx1_ASAP7_75t_L g1029 ( .A(n_175), .Y(n_1029) );
INVxp67_ASAP7_75t_L g900 ( .A(n_176), .Y(n_900) );
OAI211xp5_ASAP7_75t_L g1096 ( .A1(n_177), .A2(n_695), .B(n_1097), .C(n_1098), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g1144 ( .A(n_177), .Y(n_1144) );
INVxp67_ASAP7_75t_SL g1331 ( .A(n_178), .Y(n_1331) );
INVx1_ASAP7_75t_L g1357 ( .A(n_179), .Y(n_1357) );
OAI221xp5_ASAP7_75t_SL g1266 ( .A1(n_180), .A2(n_259), .B1(n_1267), .B2(n_1268), .C(n_1269), .Y(n_1266) );
INVx1_ASAP7_75t_L g1284 ( .A(n_180), .Y(n_1284) );
INVx1_ASAP7_75t_L g1233 ( .A(n_181), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_181), .A2(n_278), .B1(n_864), .B2(n_993), .Y(n_1245) );
INVx1_ASAP7_75t_L g433 ( .A(n_183), .Y(n_433) );
INVxp67_ASAP7_75t_SL g1062 ( .A(n_184), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_185), .A2(n_289), .B1(n_1257), .B2(n_1258), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_185), .A2(n_217), .B1(n_778), .B2(n_1297), .Y(n_1430) );
BUFx3_ASAP7_75t_L g362 ( .A(n_186), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_187), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1320 ( .A(n_189), .Y(n_1320) );
INVx1_ASAP7_75t_L g1411 ( .A(n_190), .Y(n_1411) );
OAI221xp5_ASAP7_75t_L g1734 ( .A1(n_191), .A2(n_250), .B1(n_786), .B2(n_1735), .C(n_1736), .Y(n_1734) );
OAI211xp5_ASAP7_75t_L g1740 ( .A1(n_191), .A2(n_948), .B(n_1741), .C(n_1744), .Y(n_1740) );
CKINVDCx5p33_ASAP7_75t_R g1721 ( .A(n_192), .Y(n_1721) );
OAI221xp5_ASAP7_75t_SL g632 ( .A1(n_193), .A2(n_283), .B1(n_633), .B2(n_636), .C(n_640), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_194), .A2(n_290), .B1(n_1121), .B2(n_1274), .Y(n_1422) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_195), .A2(n_233), .B1(n_1464), .B2(n_1467), .Y(n_1477) );
XOR2xp5_ASAP7_75t_L g1248 ( .A(n_197), .B(n_1249), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_198), .A2(n_235), .B1(n_1256), .B2(n_1258), .Y(n_1255) );
INVx1_ASAP7_75t_L g691 ( .A(n_199), .Y(n_691) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_200), .A2(n_375), .B(n_382), .C(n_386), .Y(n_374) );
INVx1_ASAP7_75t_L g505 ( .A(n_200), .Y(n_505) );
INVx1_ASAP7_75t_L g1018 ( .A(n_201), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_202), .Y(n_1279) );
INVx1_ASAP7_75t_L g1177 ( .A(n_203), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_204), .Y(n_772) );
INVx1_ASAP7_75t_L g1049 ( .A(n_205), .Y(n_1049) );
INVx1_ASAP7_75t_L g396 ( .A(n_206), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g492 ( .A1(n_206), .A2(n_493), .B(n_495), .C(n_500), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g1369 ( .A(n_207), .Y(n_1369) );
OAI211xp5_ASAP7_75t_L g1215 ( .A1(n_208), .A2(n_608), .B(n_695), .C(n_1216), .Y(n_1215) );
INVxp33_ASAP7_75t_SL g1239 ( .A(n_208), .Y(n_1239) );
INVx1_ASAP7_75t_L g1040 ( .A(n_209), .Y(n_1040) );
INVx1_ASAP7_75t_L g986 ( .A(n_210), .Y(n_986) );
BUFx3_ASAP7_75t_L g337 ( .A(n_211), .Y(n_337) );
INVx1_ASAP7_75t_L g516 ( .A(n_211), .Y(n_516) );
INVxp67_ASAP7_75t_SL g1205 ( .A(n_212), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1693 ( .A1(n_213), .A2(n_267), .B1(n_778), .B2(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g574 ( .A(n_214), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_218), .B(n_839), .Y(n_838) );
OAI322xp33_ASAP7_75t_SL g562 ( .A1(n_219), .A2(n_458), .A3(n_563), .B1(n_568), .B2(n_573), .C1(n_585), .C2(n_588), .Y(n_562) );
OAI22xp33_ASAP7_75t_SL g649 ( .A1(n_219), .A2(n_222), .B1(n_650), .B2(n_653), .Y(n_649) );
INVxp67_ASAP7_75t_SL g1403 ( .A(n_220), .Y(n_1403) );
INVx1_ASAP7_75t_L g781 ( .A(n_221), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g1729 ( .A(n_223), .Y(n_1729) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_224), .A2(n_287), .B1(n_580), .B2(n_926), .C(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g963 ( .A(n_224), .Y(n_963) );
INVx1_ASAP7_75t_L g928 ( .A(n_225), .Y(n_928) );
INVx1_ASAP7_75t_L g578 ( .A(n_226), .Y(n_578) );
XOR2xp5_ASAP7_75t_L g915 ( .A(n_227), .B(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g1321 ( .A(n_228), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_229), .Y(n_799) );
INVxp67_ASAP7_75t_SL g1270 ( .A(n_231), .Y(n_1270) );
OAI22xp5_ASAP7_75t_SL g532 ( .A1(n_233), .A2(n_533), .B1(n_534), .B2(n_660), .Y(n_532) );
INVx1_ASAP7_75t_L g660 ( .A(n_233), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_233), .A2(n_533), .B1(n_534), .B2(n_660), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g1044 ( .A1(n_234), .A2(n_683), .B(n_1045), .C(n_1047), .Y(n_1044) );
INVx1_ASAP7_75t_L g1080 ( .A(n_234), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_236), .Y(n_951) );
INVx1_ASAP7_75t_L g364 ( .A(n_238), .Y(n_364) );
INVx1_ASAP7_75t_L g380 ( .A(n_238), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g1366 ( .A(n_240), .Y(n_1366) );
INVx1_ASAP7_75t_L g1419 ( .A(n_241), .Y(n_1419) );
INVxp67_ASAP7_75t_SL g1443 ( .A(n_242), .Y(n_1443) );
INVxp67_ASAP7_75t_SL g1237 ( .A(n_243), .Y(n_1237) );
INVx1_ASAP7_75t_L g957 ( .A(n_244), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_245), .A2(n_277), .B1(n_920), .B2(n_923), .Y(n_919) );
INVx1_ASAP7_75t_L g952 ( .A(n_245), .Y(n_952) );
INVx1_ASAP7_75t_L g438 ( .A(n_246), .Y(n_438) );
INVxp67_ASAP7_75t_SL g1334 ( .A(n_247), .Y(n_1334) );
AOI21xp33_ASAP7_75t_L g1173 ( .A1(n_248), .A2(n_471), .B(n_678), .Y(n_1173) );
INVxp67_ASAP7_75t_L g1193 ( .A(n_248), .Y(n_1193) );
INVx1_ASAP7_75t_L g442 ( .A(n_249), .Y(n_442) );
INVx1_ASAP7_75t_L g707 ( .A(n_251), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_251), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g1399 ( .A(n_252), .Y(n_1399) );
INVx1_ASAP7_75t_L g419 ( .A(n_253), .Y(n_419) );
INVxp33_ASAP7_75t_L g895 ( .A(n_254), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_255), .Y(n_998) );
INVx1_ASAP7_75t_L g901 ( .A(n_256), .Y(n_901) );
INVx1_ASAP7_75t_L g808 ( .A(n_257), .Y(n_808) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_258), .B(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1466 ( .A(n_258), .Y(n_1466) );
INVx1_ASAP7_75t_L g1286 ( .A(n_259), .Y(n_1286) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_260), .A2(n_311), .B1(n_358), .B2(n_367), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_260), .A2(n_311), .B1(n_329), .B2(n_521), .Y(n_520) );
AOI221xp5_ASAP7_75t_SL g1131 ( .A1(n_261), .A2(n_262), .B1(n_1123), .B2(n_1132), .C(n_1133), .Y(n_1131) );
INVx1_ASAP7_75t_L g1111 ( .A(n_262), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_264), .A2(n_1091), .B1(n_1092), .B2(n_1149), .Y(n_1090) );
INVx1_ASAP7_75t_L g1149 ( .A(n_264), .Y(n_1149) );
INVx1_ASAP7_75t_L g1525 ( .A(n_265), .Y(n_1525) );
XOR2x2_ASAP7_75t_L g1153 ( .A(n_266), .B(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1046 ( .A(n_269), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_270), .Y(n_644) );
INVx1_ASAP7_75t_L g782 ( .A(n_272), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g828 ( .A1(n_272), .A2(n_726), .B1(n_829), .B2(n_834), .C(n_835), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_274), .A2(n_289), .B1(n_1297), .B2(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g873 ( .A(n_275), .Y(n_873) );
INVxp67_ASAP7_75t_SL g972 ( .A(n_277), .Y(n_972) );
INVx1_ASAP7_75t_L g1226 ( .A(n_278), .Y(n_1226) );
INVx1_ASAP7_75t_L g392 ( .A(n_279), .Y(n_392) );
INVx1_ASAP7_75t_L g1073 ( .A(n_280), .Y(n_1073) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_281), .Y(n_333) );
INVx1_ASAP7_75t_L g1166 ( .A(n_282), .Y(n_1166) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_283), .Y(n_536) );
INVx1_ASAP7_75t_L g1217 ( .A(n_284), .Y(n_1217) );
INVx1_ASAP7_75t_L g1692 ( .A(n_285), .Y(n_1692) );
CKINVDCx5p33_ASAP7_75t_R g1726 ( .A(n_286), .Y(n_1726) );
INVx1_ASAP7_75t_L g968 ( .A(n_287), .Y(n_968) );
INVx1_ASAP7_75t_L g1135 ( .A(n_288), .Y(n_1135) );
AOI21xp33_ASAP7_75t_L g1348 ( .A1(n_292), .A2(n_856), .B(n_1069), .Y(n_1348) );
INVx1_ASAP7_75t_L g572 ( .A(n_294), .Y(n_572) );
INVx1_ASAP7_75t_L g1697 ( .A(n_295), .Y(n_1697) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_296), .Y(n_1364) );
INVx1_ASAP7_75t_L g762 ( .A(n_298), .Y(n_762) );
INVx1_ASAP7_75t_L g355 ( .A(n_300), .Y(n_355) );
INVx2_ASAP7_75t_L g411 ( .A(n_300), .Y(n_411) );
INVx1_ASAP7_75t_L g484 ( .A(n_300), .Y(n_484) );
INVx1_ASAP7_75t_L g936 ( .A(n_301), .Y(n_936) );
INVx1_ASAP7_75t_L g1338 ( .A(n_302), .Y(n_1338) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_305), .Y(n_784) );
INVxp67_ASAP7_75t_SL g1188 ( .A(n_306), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_307), .Y(n_852) );
OAI21xp33_ASAP7_75t_SL g1209 ( .A1(n_308), .A2(n_713), .B(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1213 ( .A(n_308), .Y(n_1213) );
INVx1_ASAP7_75t_L g567 ( .A(n_309), .Y(n_567) );
INVx1_ASAP7_75t_L g427 ( .A(n_310), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_338), .B(n_1449), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g1706 ( .A(n_317), .B(n_326), .Y(n_1706) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g1710 ( .A(n_319), .B(n_322), .Y(n_1710) );
INVx1_ASAP7_75t_L g1754 ( .A(n_319), .Y(n_1754) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g1756 ( .A(n_322), .B(n_1754), .Y(n_1756) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g526 ( .A(n_326), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g448 ( .A(n_327), .B(n_337), .Y(n_448) );
AND2x4_ASAP7_75t_L g648 ( .A(n_327), .B(n_336), .Y(n_648) );
AND2x4_ASAP7_75t_SL g1705 ( .A(n_328), .B(n_1706), .Y(n_1705) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_330), .B(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g418 ( .A(n_330), .Y(n_418) );
OR2x6_ASAP7_75t_L g514 ( .A(n_330), .B(n_515), .Y(n_514) );
BUFx4f_ASAP7_75t_L g1346 ( .A(n_330), .Y(n_1346) );
INVxp67_ASAP7_75t_L g1375 ( .A(n_330), .Y(n_1375) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx4f_ASAP7_75t_L g452 ( .A(n_331), .Y(n_452) );
INVx3_ASAP7_75t_L g620 ( .A(n_331), .Y(n_620) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g425 ( .A(n_333), .Y(n_425) );
INVx2_ASAP7_75t_L g432 ( .A(n_333), .Y(n_432) );
NAND2x1_ASAP7_75t_L g436 ( .A(n_333), .B(n_334), .Y(n_436) );
AND2x2_ASAP7_75t_L g499 ( .A(n_333), .B(n_334), .Y(n_499) );
INVx1_ASAP7_75t_L g510 ( .A(n_333), .Y(n_510) );
AND2x2_ASAP7_75t_L g523 ( .A(n_333), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_334), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g431 ( .A(n_334), .B(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g504 ( .A(n_334), .Y(n_504) );
INVx2_ASAP7_75t_L g524 ( .A(n_334), .Y(n_524) );
INVx1_ASAP7_75t_L g600 ( .A(n_334), .Y(n_600) );
AND2x2_ASAP7_75t_L g656 ( .A(n_334), .B(n_425), .Y(n_656) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g497 ( .A(n_336), .Y(n_497) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g503 ( .A(n_337), .Y(n_503) );
AND2x4_ASAP7_75t_L g508 ( .A(n_337), .B(n_509), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_1304), .B2(n_1448), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
XNOR2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_844), .Y(n_340) );
XNOR2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_663), .Y(n_341) );
AOI22x1_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_531), .B2(n_661), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g529 ( .A(n_345), .Y(n_529) );
OAI211xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_356), .B(n_405), .C(n_491), .Y(n_345) );
CKINVDCx14_ASAP7_75t_R g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp33_ASAP7_75t_SL g461 ( .A(n_350), .B(n_366), .Y(n_461) );
INVx1_ASAP7_75t_L g552 ( .A(n_350), .Y(n_552) );
AND2x2_ASAP7_75t_L g930 ( .A(n_350), .B(n_390), .Y(n_930) );
AND3x4_ASAP7_75t_L g1289 ( .A(n_350), .B(n_390), .C(n_812), .Y(n_1289) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g447 ( .A(n_353), .Y(n_447) );
OR2x2_ASAP7_75t_L g460 ( .A(n_353), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g541 ( .A(n_353), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_SL g1083 ( .A(n_353), .B(n_448), .Y(n_1083) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g528 ( .A(n_354), .Y(n_528) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR3xp33_ASAP7_75t_SL g356 ( .A(n_357), .B(n_374), .C(n_397), .Y(n_356) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_365), .Y(n_360) );
OR2x4_ASAP7_75t_L g399 ( .A(n_361), .B(n_369), .Y(n_399) );
BUFx3_ASAP7_75t_L g465 ( .A(n_361), .Y(n_465) );
INVx2_ASAP7_75t_L g488 ( .A(n_361), .Y(n_488) );
BUFx4f_ASAP7_75t_L g802 ( .A(n_361), .Y(n_802) );
BUFx3_ASAP7_75t_L g1048 ( .A(n_361), .Y(n_1048) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_L g373 ( .A(n_362), .Y(n_373) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_362), .Y(n_381) );
AND2x4_ASAP7_75t_L g384 ( .A(n_362), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_362), .B(n_380), .Y(n_404) );
INVx1_ASAP7_75t_L g583 ( .A(n_363), .Y(n_583) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g372 ( .A(n_364), .Y(n_372) );
INVx1_ASAP7_75t_L g369 ( .A(n_365), .Y(n_369) );
AND2x4_ASAP7_75t_L g383 ( .A(n_365), .B(n_384), .Y(n_383) );
OR2x6_ASAP7_75t_L g402 ( .A(n_365), .B(n_403), .Y(n_402) );
NAND3x1_ASAP7_75t_L g482 ( .A(n_365), .B(n_483), .C(n_485), .Y(n_482) );
AND2x4_ASAP7_75t_L g551 ( .A(n_365), .B(n_552), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_365), .B(n_485), .Y(n_688) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g390 ( .A(n_366), .Y(n_390) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_370), .Y(n_899) );
BUFx6f_ASAP7_75t_L g1017 ( .A(n_370), .Y(n_1017) );
INVx2_ASAP7_75t_L g1055 ( .A(n_370), .Y(n_1055) );
INVx1_ASAP7_75t_L g1316 ( .A(n_370), .Y(n_1316) );
INVx2_ASAP7_75t_L g1439 ( .A(n_370), .Y(n_1439) );
INVx2_ASAP7_75t_L g1723 ( .A(n_370), .Y(n_1723) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_371), .Y(n_471) );
INVx2_ASAP7_75t_L g478 ( .A(n_371), .Y(n_478) );
BUFx8_ASAP7_75t_L g543 ( .A(n_371), .Y(n_543) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AND2x4_ASAP7_75t_L g582 ( .A(n_373), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x6_ASAP7_75t_L g695 ( .A(n_377), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g1326 ( .A(n_377), .Y(n_1326) );
OAI221xp5_ASAP7_75t_L g1725 ( .A1(n_377), .A2(n_687), .B1(n_802), .B2(n_1726), .C(n_1727), .Y(n_1725) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_378), .Y(n_468) );
BUFx3_ASAP7_75t_L g571 ( .A(n_378), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
BUFx2_ASAP7_75t_L g395 ( .A(n_379), .Y(n_395) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g385 ( .A(n_380), .Y(n_385) );
BUFx2_ASAP7_75t_L g391 ( .A(n_381), .Y(n_391) );
INVx2_ASAP7_75t_L g548 ( .A(n_381), .Y(n_548) );
AND2x4_ASAP7_75t_L g674 ( .A(n_381), .B(n_558), .Y(n_674) );
CKINVDCx8_ASAP7_75t_R g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g561 ( .A(n_384), .Y(n_561) );
BUFx2_ASAP7_75t_L g584 ( .A(n_384), .Y(n_584) );
BUFx2_ASAP7_75t_L g676 ( .A(n_384), .Y(n_676) );
BUFx3_ASAP7_75t_L g683 ( .A(n_384), .Y(n_683) );
BUFx2_ASAP7_75t_L g709 ( .A(n_384), .Y(n_709) );
AND2x2_ASAP7_75t_L g924 ( .A(n_384), .B(n_922), .Y(n_924) );
INVx2_ASAP7_75t_L g1021 ( .A(n_384), .Y(n_1021) );
INVx1_ASAP7_75t_L g558 ( .A(n_385), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_392), .B1(n_393), .B2(n_396), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
AND2x4_ASAP7_75t_L g394 ( .A(n_389), .B(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_392), .A2(n_501), .B1(n_505), .B2(n_506), .Y(n_500) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx3_ASAP7_75t_L g479 ( .A(n_403), .Y(n_479) );
INVx1_ASAP7_75t_L g705 ( .A(n_403), .Y(n_705) );
BUFx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g474 ( .A(n_404), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_457), .Y(n_405) );
OAI33xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_413), .A3(n_426), .B1(n_437), .B2(n_443), .B3(n_449), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_407), .A2(n_743), .B(n_754), .Y(n_742) );
INVx1_ASAP7_75t_L g1137 ( .A(n_407), .Y(n_1137) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx4_ASAP7_75t_L g818 ( .A(n_409), .Y(n_818) );
AOI222xp33_ASAP7_75t_L g953 ( .A1(n_409), .A2(n_741), .B1(n_954), .B2(n_957), .C1(n_958), .C2(n_965), .Y(n_953) );
INVx2_ASAP7_75t_L g1069 ( .A(n_409), .Y(n_1069) );
INVx2_ASAP7_75t_L g1186 ( .A(n_409), .Y(n_1186) );
AOI31xp33_ASAP7_75t_L g1414 ( .A1(n_409), .A2(n_977), .A3(n_1415), .B(n_1416), .Y(n_1414) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g659 ( .A(n_410), .Y(n_659) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_411), .B(n_598), .Y(n_757) );
INVx2_ASAP7_75t_L g812 ( .A(n_411), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_419), .B2(n_420), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_414), .A2(n_438), .B1(n_463), .B2(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_417), .A2(n_968), .B1(n_969), .B2(n_970), .Y(n_967) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_419), .A2(n_442), .B1(n_487), .B2(n_489), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_420), .A2(n_1321), .B1(n_1346), .B2(n_1347), .Y(n_1345) );
INVx5_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx6_ASAP7_75t_L g740 ( .A(n_421), .Y(n_740) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g455 ( .A(n_422), .Y(n_455) );
INVx4_ASAP7_75t_L g623 ( .A(n_422), .Y(n_623) );
INVx2_ASAP7_75t_SL g970 ( .A(n_422), .Y(n_970) );
INVx2_ASAP7_75t_L g1076 ( .A(n_422), .Y(n_1076) );
INVx1_ASAP7_75t_L g1271 ( .A(n_422), .Y(n_1271) );
INVx8_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g519 ( .A(n_423), .B(n_503), .Y(n_519) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_423), .Y(n_1191) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_433), .B2(n_434), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_427), .A2(n_453), .B1(n_470), .B2(n_472), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_428), .A2(n_438), .B1(n_439), .B2(n_442), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_428), .A2(n_784), .B1(n_799), .B2(n_830), .C(n_831), .Y(n_829) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g1071 ( .A(n_429), .Y(n_1071) );
INVx4_ASAP7_75t_L g1368 ( .A(n_429), .Y(n_1368) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g746 ( .A(n_431), .Y(n_746) );
INVx2_ASAP7_75t_L g821 ( .A(n_431), .Y(n_821) );
INVx1_ASAP7_75t_L g1195 ( .A(n_431), .Y(n_1195) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_431), .Y(n_1197) );
AND2x2_ASAP7_75t_L g599 ( .A(n_432), .B(n_600), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_433), .A2(n_456), .B1(n_476), .B2(n_479), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g1196 ( .A1(n_434), .A2(n_1161), .B1(n_1171), .B2(n_1197), .Y(n_1196) );
OAI221xp5_ASAP7_75t_L g1748 ( .A1(n_434), .A2(n_1721), .B1(n_1726), .B2(n_1749), .C(n_1750), .Y(n_1748) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx4_ASAP7_75t_L g749 ( .A(n_435), .Y(n_749) );
OR2x6_ASAP7_75t_L g754 ( .A(n_435), .B(n_755), .Y(n_754) );
BUFx4f_ASAP7_75t_L g823 ( .A(n_435), .Y(n_823) );
BUFx4f_ASAP7_75t_L g830 ( .A(n_435), .Y(n_830) );
BUFx4f_ASAP7_75t_L g999 ( .A(n_435), .Y(n_999) );
BUFx4f_ASAP7_75t_L g1072 ( .A(n_435), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g441 ( .A(n_436), .Y(n_441) );
OAI211xp5_ASAP7_75t_L g1680 ( .A1(n_439), .A2(n_1681), .B(n_1682), .C(n_1684), .Y(n_1680) );
INVx5_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g494 ( .A(n_441), .Y(n_494) );
OR2x2_ASAP7_75t_L g726 ( .A(n_441), .B(n_723), .Y(n_726) );
OR2x2_ASAP7_75t_L g975 ( .A(n_441), .B(n_723), .Y(n_975) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g1745 ( .A1(n_445), .A2(n_1186), .B1(n_1746), .B2(n_1748), .Y(n_1745) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
AND2x4_ASAP7_75t_L g741 ( .A(n_446), .B(n_448), .Y(n_741) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx4_ASAP7_75t_L g629 ( .A(n_448), .Y(n_629) );
INVx4_ASAP7_75t_L g991 ( .A(n_448), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B1(n_454), .B2(n_456), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g1075 ( .A(n_451), .Y(n_1075) );
INVx2_ASAP7_75t_L g1134 ( .A(n_451), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g643 ( .A(n_452), .Y(n_643) );
INVx4_ASAP7_75t_L g964 ( .A(n_452), .Y(n_964) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI33xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_462), .A3(n_469), .B1(n_475), .B2(n_480), .B3(n_486), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx8_ASAP7_75t_L g893 ( .A(n_460), .Y(n_893) );
BUFx2_ASAP7_75t_L g678 ( .A(n_461), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_463), .A2(n_569), .B1(n_570), .B2(n_572), .Y(n_568) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_465), .A2(n_571), .B1(n_687), .B2(n_1057), .C(n_1058), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_465), .A2(n_687), .B1(n_1162), .B2(n_1229), .C(n_1230), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1396 ( .A1(n_465), .A2(n_571), .B1(n_687), .B2(n_1364), .C(n_1372), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g1220 ( .A1(n_467), .A2(n_930), .B1(n_1009), .B2(n_1221), .C(n_1222), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g490 ( .A(n_468), .Y(n_490) );
OR2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_541), .Y(n_606) );
INVx4_ASAP7_75t_L g1163 ( .A(n_468), .Y(n_1163) );
OAI221xp5_ASAP7_75t_L g1720 ( .A1(n_468), .A2(n_930), .B1(n_1721), .B2(n_1722), .C(n_1723), .Y(n_1720) );
INVx2_ASAP7_75t_L g677 ( .A(n_470), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g927 ( .A1(n_470), .A2(n_571), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_927) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g577 ( .A(n_471), .Y(n_577) );
INVx2_ASAP7_75t_SL g681 ( .A(n_471), .Y(n_681) );
INVx5_ASAP7_75t_L g1433 ( .A(n_471), .Y(n_1433) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
CKINVDCx8_ASAP7_75t_R g807 ( .A(n_473), .Y(n_807) );
INVx1_ASAP7_75t_L g1050 ( .A(n_473), .Y(n_1050) );
INVx3_ASAP7_75t_L g1227 ( .A(n_473), .Y(n_1227) );
INVx3_ASAP7_75t_L g1730 ( .A(n_473), .Y(n_1730) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g595 ( .A(n_474), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g1394 ( .A1(n_476), .A2(n_571), .B1(n_930), .B2(n_1369), .C(n_1371), .Y(n_1394) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g1735 ( .A(n_477), .Y(n_1735) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g566 ( .A(n_478), .Y(n_566) );
OR2x6_ASAP7_75t_SL g794 ( .A(n_478), .B(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_478), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_479), .A2(n_564), .B1(n_565), .B2(n_567), .Y(n_563) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_479), .A2(n_574), .B1(n_575), .B2(n_578), .C(n_579), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_479), .A2(n_898), .B1(n_900), .B2(n_901), .C(n_902), .Y(n_897) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g1022 ( .A(n_481), .Y(n_1022) );
AOI33xp33_ASAP7_75t_L g1287 ( .A1(n_481), .A2(n_1288), .A3(n_1290), .B1(n_1293), .B2(n_1298), .B3(n_1299), .Y(n_1287) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g587 ( .A(n_482), .Y(n_587) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_484), .B(n_616), .Y(n_723) );
OR2x2_ASAP7_75t_L g588 ( .A(n_487), .B(n_589), .Y(n_588) );
OR2x6_ASAP7_75t_L g909 ( .A(n_487), .B(n_589), .Y(n_909) );
INVx2_ASAP7_75t_SL g1104 ( .A(n_487), .Y(n_1104) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g1225 ( .A(n_488), .Y(n_1225) );
OAI22xp33_ASAP7_75t_L g894 ( .A1(n_489), .A2(n_800), .B1(n_895), .B2(n_896), .Y(n_894) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g786 ( .A(n_490), .Y(n_786) );
INVx3_ASAP7_75t_L g1172 ( .A(n_490), .Y(n_1172) );
OAI31xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_511), .A3(n_520), .B(n_525), .Y(n_491) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_494), .A2(n_1166), .B1(n_1193), .B2(n_1194), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_494), .A2(n_1078), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x4_ASAP7_75t_SL g615 ( .A(n_498), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g626 ( .A(n_498), .Y(n_626) );
AND2x6_ASAP7_75t_L g631 ( .A(n_498), .B(n_598), .Y(n_631) );
BUFx3_ASAP7_75t_L g736 ( .A(n_498), .Y(n_736) );
BUFx3_ASAP7_75t_L g856 ( .A(n_498), .Y(n_856) );
BUFx3_ASAP7_75t_L g966 ( .A(n_498), .Y(n_966) );
BUFx3_ASAP7_75t_L g989 ( .A(n_498), .Y(n_989) );
BUFx6f_ASAP7_75t_L g1125 ( .A(n_498), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g1276 ( .A(n_499), .Y(n_1276) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g638 ( .A(n_504), .Y(n_638) );
INVx1_ASAP7_75t_L g761 ( .A(n_504), .Y(n_761) );
BUFx2_ASAP7_75t_L g866 ( .A(n_504), .Y(n_866) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_509), .B(n_598), .Y(n_605) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g522 ( .A(n_515), .B(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_523), .Y(n_628) );
BUFx3_ASAP7_75t_L g646 ( .A(n_523), .Y(n_646) );
INVx2_ASAP7_75t_L g735 ( .A(n_523), .Y(n_735) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g604 ( .A(n_528), .B(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g609 ( .A(n_528), .Y(n_609) );
INVx1_ASAP7_75t_L g715 ( .A(n_528), .Y(n_715) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_528), .B(n_605), .Y(n_1148) );
INVxp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND3x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_591), .C(n_610), .Y(n_534) );
AOI211xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_537), .B(n_544), .C(n_562), .Y(n_535) );
INVxp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_539), .A2(n_985), .B1(n_986), .B2(n_1033), .Y(n_1032) );
INVx2_ASAP7_75t_L g1301 ( .A(n_539), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g1699 ( .A1(n_539), .A2(n_1677), .B1(n_1678), .B2(n_1700), .Y(n_1699) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_540), .B(n_1034), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1700 ( .A(n_540), .B(n_1034), .Y(n_1700) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
OR2x2_ASAP7_75t_L g594 ( .A(n_541), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g701 ( .A(n_542), .Y(n_701) );
INVx1_ASAP7_75t_L g922 ( .A(n_542), .Y(n_922) );
INVx3_ASAP7_75t_L g789 ( .A(n_543), .Y(n_789) );
INVx2_ASAP7_75t_SL g805 ( .A(n_543), .Y(n_805) );
INVx2_ASAP7_75t_SL g933 ( .A(n_543), .Y(n_933) );
INVx3_ASAP7_75t_L g1009 ( .A(n_543), .Y(n_1009) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x6_ASAP7_75t_L g690 ( .A(n_547), .B(n_551), .Y(n_690) );
NAND2x1_ASAP7_75t_L g912 ( .A(n_547), .B(n_549), .Y(n_912) );
AND2x4_ASAP7_75t_SL g1025 ( .A(n_547), .B(n_549), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_547), .B(n_549), .Y(n_1285) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g554 ( .A(n_549), .B(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g560 ( .A(n_549), .B(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_SL g1027 ( .A(n_549), .B(n_555), .Y(n_1027) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
OR2x2_ASAP7_75t_L g596 ( .A(n_550), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g955 ( .A(n_550), .Y(n_955) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_551), .B(n_582), .Y(n_608) );
AND2x2_ASAP7_75t_L g692 ( .A(n_551), .B(n_557), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_551), .Y(n_696) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_554), .A2(n_867), .B1(n_873), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_554), .A2(n_1284), .B1(n_1285), .B2(n_1286), .Y(n_1283) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g913 ( .A(n_560), .Y(n_913) );
NOR3xp33_ASAP7_75t_L g1006 ( .A(n_560), .B(n_1007), .C(n_1023), .Y(n_1006) );
NOR3xp33_ASAP7_75t_L g1685 ( .A(n_560), .B(n_1686), .C(n_1695), .Y(n_1685) );
BUFx2_ASAP7_75t_L g1292 ( .A(n_561), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_561), .A2(n_1407), .B1(n_1419), .B2(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g890 ( .A(n_566), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_567), .A2(n_578), .B1(n_618), .B2(n_621), .C(n_624), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_569), .A2(n_621), .B1(n_641), .B2(n_644), .C(n_645), .Y(n_640) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g798 ( .A(n_571), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_571), .A2(n_687), .B1(n_802), .B2(n_935), .C(n_936), .Y(n_934) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g1728 ( .A1(n_577), .A2(n_1729), .B1(n_1730), .B2(n_1731), .Y(n_1728) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_580), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_706) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx8_ASAP7_75t_L g778 ( .A(n_581), .Y(n_778) );
INVx2_ASAP7_75t_L g1034 ( .A(n_581), .Y(n_1034) );
INVx3_ASAP7_75t_L g1441 ( .A(n_581), .Y(n_1441) );
INVx8_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx3_ASAP7_75t_L g672 ( .A(n_582), .Y(n_672) );
BUFx3_ASAP7_75t_L g685 ( .A(n_582), .Y(n_685) );
AND2x2_ASAP7_75t_L g921 ( .A(n_582), .B(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g904 ( .A(n_587), .Y(n_904) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_601), .B(n_602), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_592), .A2(n_884), .B1(n_906), .B2(n_907), .C(n_908), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g1028 ( .A1(n_592), .A2(n_1029), .B(n_1030), .Y(n_1028) );
AOI21xp5_ASAP7_75t_L g1278 ( .A1(n_592), .A2(n_1279), .B(n_1280), .Y(n_1278) );
AOI21xp5_ASAP7_75t_L g1696 ( .A1(n_592), .A2(n_1697), .B(n_1698), .Y(n_1696) );
INVx8_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
BUFx3_ASAP7_75t_L g892 ( .A(n_595), .Y(n_892) );
INVx1_ASAP7_75t_L g1168 ( .A(n_595), .Y(n_1168) );
INVx1_ASAP7_75t_L g719 ( .A(n_596), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_596), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g956 ( .A(n_597), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g639 ( .A(n_598), .Y(n_639) );
AND2x2_ASAP7_75t_L g865 ( .A(n_598), .B(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g652 ( .A(n_599), .B(n_616), .Y(n_652) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_599), .Y(n_752) );
INVx3_ASAP7_75t_L g826 ( .A(n_599), .Y(n_826) );
INVx2_ASAP7_75t_L g851 ( .A(n_603), .Y(n_851) );
AND2x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx2_ASAP7_75t_SL g837 ( .A(n_604), .Y(n_837) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_604), .B(n_606), .Y(n_1031) );
INVx3_ASAP7_75t_L g906 ( .A(n_607), .Y(n_906) );
OR2x6_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g711 ( .A(n_608), .Y(n_711) );
OR2x2_ASAP7_75t_L g770 ( .A(n_608), .B(n_609), .Y(n_770) );
OAI31xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_632), .A3(n_649), .B(n_657), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g995 ( .A(n_613), .Y(n_995) );
INVx2_ASAP7_75t_L g1267 ( .A(n_613), .Y(n_1267) );
INVx4_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g872 ( .A(n_615), .Y(n_872) );
AND2x4_ASAP7_75t_L g635 ( .A(n_616), .B(n_628), .Y(n_635) );
AND2x4_ASAP7_75t_L g654 ( .A(n_616), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g731 ( .A(n_616), .B(n_628), .Y(n_731) );
AND2x2_ASAP7_75t_L g983 ( .A(n_616), .B(n_724), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_618), .A2(n_1169), .B1(n_1191), .B2(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
BUFx3_ASAP7_75t_L g1085 ( .A(n_620), .Y(n_1085) );
BUFx6f_ASAP7_75t_L g1189 ( .A(n_620), .Y(n_1189) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_623), .A2(n_936), .B1(n_963), .B2(n_964), .Y(n_962) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g959 ( .A(n_626), .Y(n_959) );
BUFx3_ASAP7_75t_L g1343 ( .A(n_627), .Y(n_1343) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g859 ( .A(n_628), .Y(n_859) );
INVx1_ASAP7_75t_L g1673 ( .A(n_628), .Y(n_1673) );
HB1xp67_ASAP7_75t_SL g878 ( .A(n_629), .Y(n_878) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_631), .A2(n_872), .B1(n_873), .B2(n_874), .C(n_879), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g987 ( .A1(n_631), .A2(n_988), .B(n_992), .Y(n_987) );
AOI21xp5_ASAP7_75t_L g1252 ( .A1(n_631), .A2(n_1253), .B(n_1255), .Y(n_1252) );
AOI21xp5_ASAP7_75t_L g1670 ( .A1(n_631), .A2(n_1671), .B(n_1674), .Y(n_1670) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx6f_ASAP7_75t_L g882 ( .A(n_635), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_635), .A2(n_651), .B1(n_985), .B2(n_986), .Y(n_984) );
INVx1_ASAP7_75t_L g1265 ( .A(n_635), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1676 ( .A1(n_635), .A2(n_652), .B1(n_1677), .B2(n_1678), .Y(n_1676) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g996 ( .A(n_637), .Y(n_996) );
NOR2x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_643), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g961 ( .A(n_646), .Y(n_961) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_646), .Y(n_1254) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g860 ( .A(n_648), .Y(n_860) );
INVx2_ASAP7_75t_L g1001 ( .A(n_648), .Y(n_1001) );
INVx1_ASAP7_75t_L g1683 ( .A(n_648), .Y(n_1683) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
HB1xp67_ASAP7_75t_L g1262 ( .A(n_651), .Y(n_1262) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g714 ( .A(n_652), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g869 ( .A(n_652), .Y(n_869) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_654), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
INVx2_ASAP7_75t_SL g1669 ( .A(n_654), .Y(n_1669) );
BUFx2_ASAP7_75t_L g827 ( .A(n_655), .Y(n_827) );
INVx1_ASAP7_75t_L g1259 ( .A(n_655), .Y(n_1259) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g725 ( .A(n_656), .Y(n_725) );
BUFx3_ASAP7_75t_L g753 ( .A(n_656), .Y(n_753) );
BUFx3_ASAP7_75t_L g864 ( .A(n_656), .Y(n_864) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_658), .A2(n_667), .B(n_712), .Y(n_666) );
INVx2_ASAP7_75t_L g944 ( .A(n_658), .Y(n_944) );
OAI31xp33_ASAP7_75t_SL g1094 ( .A1(n_658), .A2(n_1095), .A3(n_1096), .B(n_1101), .Y(n_1094) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_659), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
XNOR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_764), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_762), .B(n_763), .Y(n_664) );
AND3x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_716), .C(n_732), .Y(n_665) );
AOI31xp33_ASAP7_75t_L g763 ( .A1(n_666), .A2(n_716), .A3(n_732), .B(n_762), .Y(n_763) );
NAND3xp33_ASAP7_75t_SL g667 ( .A(n_668), .B(n_689), .C(n_697), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_675), .B1(n_679), .B2(n_682), .Y(n_668) );
BUFx2_ASAP7_75t_SL g1291 ( .A(n_670), .Y(n_1291) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g1319 ( .A1(n_671), .A2(n_792), .B1(n_930), .B2(n_1320), .C(n_1321), .Y(n_1319) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_672), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_672), .B(n_1737), .Y(n_1736) );
BUFx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx5_ASAP7_75t_L g792 ( .A(n_674), .Y(n_792) );
AND2x4_ASAP7_75t_L g842 ( .A(n_674), .B(n_701), .Y(n_842) );
BUFx3_ASAP7_75t_L g926 ( .A(n_674), .Y(n_926) );
BUFx12f_ASAP7_75t_L g1297 ( .A(n_674), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_676), .A2(n_772), .B1(n_778), .B2(n_779), .Y(n_777) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g1393 ( .A(n_685), .Y(n_1393) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g796 ( .A1(n_687), .A2(n_797), .B1(n_799), .B2(n_800), .C(n_803), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_687), .B(n_1328), .Y(n_1327) );
INVx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_692), .B2(n_693), .C(n_694), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_690), .A2(n_692), .B1(n_781), .B2(n_782), .Y(n_780) );
INVx4_ASAP7_75t_L g942 ( .A(n_690), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_690), .A2(n_692), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_690), .A2(n_692), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
INVx2_ASAP7_75t_L g943 ( .A(n_692), .Y(n_943) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_692), .Y(n_1428) );
NOR3xp33_ASAP7_75t_L g1390 ( .A(n_694), .B(n_1391), .C(n_1395), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1425 ( .A(n_694), .B(n_1426), .Y(n_1425) );
NOR3xp33_ASAP7_75t_L g1718 ( .A(n_694), .B(n_1719), .C(n_1724), .Y(n_1718) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B1(n_710), .B2(n_711), .Y(n_697) );
INVxp67_ASAP7_75t_L g776 ( .A(n_698), .Y(n_776) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g1388 ( .A(n_700), .Y(n_1388) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g795 ( .A(n_701), .Y(n_795) );
OAI21xp33_ASAP7_75t_L g1012 ( .A1(n_703), .A2(n_1013), .B(n_1014), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1687 ( .A1(n_703), .A2(n_805), .B1(n_1688), .B2(n_1689), .C(n_1690), .Y(n_1687) );
INVx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_709), .Y(n_1108) );
AOI211xp5_ASAP7_75t_SL g937 ( .A1(n_711), .A2(n_938), .B(n_939), .C(n_941), .Y(n_937) );
AOI211xp5_ASAP7_75t_L g1039 ( .A1(n_711), .A2(n_1040), .B(n_1041), .C(n_1042), .Y(n_1039) );
INVx2_ASAP7_75t_L g1097 ( .A(n_711), .Y(n_1097) );
AOI211xp5_ASAP7_75t_L g1156 ( .A1(n_711), .A2(n_1157), .B(n_1158), .C(n_1159), .Y(n_1156) );
AOI211xp5_ASAP7_75t_SL g1309 ( .A1(n_711), .A2(n_1310), .B(n_1311), .C(n_1312), .Y(n_1309) );
AOI221xp5_ASAP7_75t_L g1386 ( .A1(n_711), .A2(n_1381), .B1(n_1387), .B2(n_1388), .C(n_1389), .Y(n_1386) );
AOI221xp5_ASAP7_75t_L g1732 ( .A1(n_711), .A2(n_1388), .B1(n_1733), .B2(n_1734), .C(n_1738), .Y(n_1732) );
INVx1_ASAP7_75t_L g1182 ( .A(n_713), .Y(n_1182) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI222xp33_ASAP7_75t_L g767 ( .A1(n_714), .A2(n_730), .B1(n_768), .B2(n_769), .C1(n_772), .C2(n_773), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_714), .B(n_972), .Y(n_971) );
AOI211xp5_ASAP7_75t_L g1333 ( .A1(n_714), .A2(n_1334), .B(n_1335), .C(n_1340), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_714), .B(n_1384), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_714), .B(n_1407), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1739 ( .A(n_714), .B(n_1737), .Y(n_1739) );
AND2x4_ASAP7_75t_L g730 ( .A(n_715), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_727), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g771 ( .A(n_721), .Y(n_771) );
AOI222xp33_ASAP7_75t_L g950 ( .A1(n_721), .A2(n_836), .B1(n_837), .B2(n_938), .C1(n_951), .C2(n_952), .Y(n_950) );
AOI222xp33_ASAP7_75t_L g1061 ( .A1(n_721), .A2(n_954), .B1(n_974), .B2(n_1040), .C1(n_1062), .C2(n_1063), .Y(n_1061) );
AOI211xp5_ASAP7_75t_L g1143 ( .A1(n_721), .A2(n_1144), .B(n_1145), .C(n_1146), .Y(n_1143) );
AOI222xp33_ASAP7_75t_L g1204 ( .A1(n_721), .A2(n_954), .B1(n_974), .B2(n_1157), .C1(n_1178), .C2(n_1205), .Y(n_1204) );
AOI21xp33_ASAP7_75t_L g1238 ( .A1(n_721), .A2(n_1239), .B(n_1240), .Y(n_1238) );
INVx1_ASAP7_75t_L g1336 ( .A(n_721), .Y(n_1336) );
AOI222xp33_ASAP7_75t_L g1379 ( .A1(n_721), .A2(n_954), .B1(n_974), .B2(n_1380), .C1(n_1381), .C2(n_1382), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_721), .A2(n_974), .B1(n_1411), .B2(n_1412), .Y(n_1410) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
AOI332xp33_ASAP7_75t_L g1741 ( .A1(n_722), .A2(n_724), .A3(n_955), .B1(n_956), .B2(n_974), .B3(n_1733), .C1(n_1742), .C2(n_1743), .Y(n_1741) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g1004 ( .A(n_725), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g948 ( .A(n_730), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_730), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1141 ( .A(n_730), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_730), .B(n_1177), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_730), .B(n_1237), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_730), .B(n_1331), .Y(n_1330) );
NAND2xp33_ASAP7_75t_SL g1398 ( .A(n_730), .B(n_1399), .Y(n_1398) );
AOI211xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_741), .B(n_742), .C(n_758), .Y(n_732) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g877 ( .A(n_735), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_741), .Y(n_834) );
AOI322xp5_ASAP7_75t_L g1119 ( .A1(n_741), .A2(n_954), .A3(n_1120), .B1(n_1126), .B2(n_1130), .C1(n_1131), .C2(n_1137), .Y(n_1119) );
AOI332xp33_ASAP7_75t_L g1241 ( .A1(n_741), .A2(n_817), .A3(n_954), .B1(n_1242), .B2(n_1243), .B3(n_1244), .C1(n_1245), .C2(n_1246), .Y(n_1241) );
AOI322xp5_ASAP7_75t_L g1341 ( .A1(n_741), .A2(n_954), .A3(n_1342), .B1(n_1344), .B2(n_1348), .C1(n_1349), .C2(n_1350), .Y(n_1341) );
NAND3xp33_ASAP7_75t_L g1420 ( .A(n_741), .B(n_1421), .C(n_1422), .Y(n_1420) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_747), .B1(n_748), .B2(n_750), .C(n_751), .Y(n_743) );
INVx3_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g1746 ( .A1(n_746), .A2(n_823), .B1(n_1722), .B2(n_1729), .C(n_1747), .Y(n_1746) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g1081 ( .A(n_749), .Y(n_1081) );
INVx2_ASAP7_75t_L g1367 ( .A(n_749), .Y(n_1367) );
INVx3_ASAP7_75t_L g833 ( .A(n_752), .Y(n_833) );
BUFx6f_ASAP7_75t_L g1257 ( .A(n_752), .Y(n_1257) );
OAI21xp5_ASAP7_75t_SL g814 ( .A1(n_754), .A2(n_815), .B(n_819), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g977 ( .A(n_754), .Y(n_977) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2x2_ASAP7_75t_L g759 ( .A(n_756), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g836 ( .A(n_759), .Y(n_836) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_759), .Y(n_1147) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_759), .Y(n_1203) );
INVx2_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_774), .C(n_813), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_793), .B(n_809), .Y(n_774) );
OAI211xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B(n_780), .C(n_783), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_779), .A2(n_781), .B1(n_836), .B2(n_837), .Y(n_835) );
OAI211xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B(n_787), .C(n_790), .Y(n_783) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_789), .A2(n_1227), .B1(n_1366), .B2(n_1377), .Y(n_1397) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_794), .Y(n_1176) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g1691 ( .A1(n_805), .A2(n_807), .B1(n_1681), .B2(n_1692), .C(n_1693), .Y(n_1691) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_806), .A2(n_820), .B1(n_822), .B2(n_823), .C(n_824), .Y(n_819) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_807), .A2(n_998), .B1(n_1016), .B2(n_1018), .C(n_1019), .Y(n_1015) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g886 ( .A(n_810), .Y(n_886) );
A2O1A1Ixp33_ASAP7_75t_SL g1155 ( .A1(n_810), .A2(n_1156), .B(n_1175), .C(n_1180), .Y(n_1155) );
BUFx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_811), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1277 ( .A(n_811), .Y(n_1277) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI31xp33_ASAP7_75t_SL g1210 ( .A1(n_812), .A2(n_1211), .A3(n_1215), .B(n_1219), .Y(n_1210) );
INVx2_ASAP7_75t_SL g1329 ( .A(n_812), .Y(n_1329) );
AOI22xp33_ASAP7_75t_SL g1423 ( .A1(n_812), .A2(n_947), .B1(n_1424), .B2(n_1443), .Y(n_1423) );
NOR3xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_828), .C(n_838), .Y(n_813) );
INVxp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_821), .Y(n_1079) );
INVx2_ASAP7_75t_L g1749 ( .A(n_821), .Y(n_1749) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g862 ( .A(n_826), .Y(n_862) );
INVx2_ASAP7_75t_SL g993 ( .A(n_826), .Y(n_993) );
INVx1_ASAP7_75t_L g1003 ( .A(n_826), .Y(n_1003) );
INVx1_ASAP7_75t_L g1127 ( .A(n_826), .Y(n_1127) );
INVx2_ASAP7_75t_L g1675 ( .A(n_826), .Y(n_1675) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_836), .A2(n_837), .B1(n_1338), .B2(n_1339), .Y(n_1337) );
AOI22xp33_ASAP7_75t_SL g1417 ( .A1(n_836), .A2(n_837), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx3_ASAP7_75t_L g940 ( .A(n_842), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_842), .A2(n_1176), .B1(n_1177), .B2(n_1178), .C(n_1179), .Y(n_1175) );
XNOR2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_1088), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_1035), .B1(n_1036), .B2(n_1087), .Y(n_845) );
INVx1_ASAP7_75t_L g1087 ( .A(n_846), .Y(n_1087) );
XOR2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_914), .Y(n_846) );
XNOR2x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
AND2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_905), .Y(n_849) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_853), .B2(n_885), .C(n_887), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_871), .C(n_881), .Y(n_853) );
AOI222xp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_861), .B1(n_865), .B2(n_867), .C1(n_868), .C2(n_870), .Y(n_854) );
BUFx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g990 ( .A(n_859), .Y(n_990) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_864), .Y(n_880) );
INVx1_ASAP7_75t_SL g1129 ( .A(n_864), .Y(n_1129) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g1122 ( .A(n_877), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_877), .Y(n_1132) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g1102 ( .A1(n_892), .A2(n_1103), .B1(n_1105), .B2(n_1106), .C(n_1107), .Y(n_1102) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_892), .A2(n_1110), .B1(n_1111), .B2(n_1112), .C(n_1113), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_893), .Y(n_1011) );
OAI22xp5_ASAP7_75t_SL g1686 ( .A1(n_893), .A2(n_1022), .B1(n_1687), .B2(n_1691), .Y(n_1686) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g1110 ( .A(n_899), .Y(n_1110) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx2_ASAP7_75t_SL g1302 ( .A(n_913), .Y(n_1302) );
XNOR2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_978), .Y(n_914) );
OR2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_949), .Y(n_916) );
A2O1A1Ixp33_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_937), .B(n_944), .C(n_945), .Y(n_917) );
NOR3xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_925), .C(n_931), .Y(n_918) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_921), .A2(n_924), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g1212 ( .A1(n_921), .A2(n_924), .B1(n_1213), .B2(n_1214), .Y(n_1212) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
OAI21xp33_ASAP7_75t_L g1045 ( .A1(n_930), .A2(n_1009), .B(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_933), .A2(n_1166), .B1(n_1167), .B2(n_1169), .Y(n_1165) );
INVx1_ASAP7_75t_L g1059 ( .A(n_944), .Y(n_1059) );
A2O1A1Ixp33_ASAP7_75t_L g1385 ( .A1(n_944), .A2(n_1386), .B(n_1390), .C(n_1398), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
NAND4xp25_ASAP7_75t_L g949 ( .A(n_950), .B(n_953), .C(n_971), .D(n_973), .Y(n_949) );
AND2x4_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_970), .A2(n_1051), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_970), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_970), .A2(n_1346), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_970), .A2(n_1374), .B1(n_1376), .B2(n_1377), .Y(n_1373) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_974), .A2(n_976), .B(n_977), .Y(n_973) );
AOI21xp5_ASAP7_75t_L g1235 ( .A1(n_974), .A2(n_977), .B(n_1218), .Y(n_1235) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
OR3x1_ASAP7_75t_L g1066 ( .A(n_977), .B(n_1067), .C(n_1068), .Y(n_1066) );
NOR3xp33_ASAP7_75t_L g1744 ( .A(n_977), .B(n_1745), .C(n_1751), .Y(n_1744) );
AND4x1_ASAP7_75t_L g979 ( .A(n_980), .B(n_1006), .C(n_1028), .D(n_1032), .Y(n_979) );
OAI21xp33_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_994), .B(n_1005), .Y(n_980) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_996), .Y(n_1268) );
OAI211xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .B(n_1000), .C(n_1002), .Y(n_997) );
A2O1A1Ixp33_ASAP7_75t_L g1717 ( .A1(n_1005), .A2(n_1718), .B(n_1732), .C(n_1739), .Y(n_1717) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1012), .B1(n_1015), .B2(n_1022), .Y(n_1007) );
OAI21xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B(n_1011), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_1009), .A2(n_1167), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1009), .Y(n_1436) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g1694 ( .A(n_1021), .Y(n_1694) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
AOI211x1_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1059), .B(n_1060), .C(n_1066), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1043), .Y(n_1038) );
NOR3xp33_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1052), .C(n_1053), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_1046), .A2(n_1071), .B1(n_1072), .B2(n_1073), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_1049), .A2(n_1058), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_1057), .A2(n_1078), .B1(n_1080), .B2(n_1081), .Y(n_1077) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .A3(n_1074), .B1(n_1077), .B2(n_1082), .B3(n_1084), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_1076), .A2(n_1085), .B1(n_1320), .B2(n_1353), .Y(n_1352) );
INVx4_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OAI33xp33_ASAP7_75t_L g1361 ( .A1(n_1082), .A2(n_1186), .A3(n_1362), .B1(n_1365), .B2(n_1370), .B3(n_1373), .Y(n_1361) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1083), .Y(n_1200) );
OA22x2_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1150), .B1(n_1151), .B2(n_1303), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1090), .Y(n_1303) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
NOR2x1_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1118), .Y(n_1092) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1097), .Y(n_1442) );
NAND3xp33_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1109), .C(n_1115), .Y(n_1101) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
OAI22xp5_ASAP7_75t_SL g1133 ( .A1(n_1105), .A2(n_1134), .B1(n_1135), .B2(n_1136), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1138), .Y(n_1118) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1351 ( .A(n_1125), .Y(n_1351) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_1129), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g1269 ( .A1(n_1134), .A2(n_1270), .B1(n_1271), .B2(n_1272), .C(n_1273), .Y(n_1269) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1140), .B(n_1142), .Y(n_1138) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
XNOR2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1248), .Y(n_1151) );
XNOR2xp5_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1207), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1183), .Y(n_1154) );
OAI21xp33_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1165), .B(n_1170), .Y(n_1159) );
OAI21xp33_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1162), .B(n_1164), .Y(n_1160) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx2_ASAP7_75t_L g1318 ( .A(n_1163), .Y(n_1318) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
OAI211xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1172), .B(n_1173), .C(n_1174), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
NAND3xp33_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1204), .C(n_1206), .Y(n_1183) );
NOR2xp33_ASAP7_75t_SL g1184 ( .A(n_1185), .B(n_1201), .Y(n_1184) );
OAI33xp33_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1187), .A3(n_1192), .B1(n_1196), .B2(n_1198), .B3(n_1200), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1189), .B1(n_1190), .B2(n_1191), .Y(n_1187) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
XOR2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1247), .Y(n_1207) );
NOR2xp33_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1234), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_1220), .A2(n_1223), .B1(n_1228), .B2(n_1231), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B1(n_1226), .B2(n_1227), .Y(n_1223) );
NAND4xp25_ASAP7_75t_SL g1234 ( .A(n_1235), .B(n_1236), .C(n_1238), .D(n_1241), .Y(n_1234) );
NAND3xp33_ASAP7_75t_SL g1249 ( .A(n_1250), .B(n_1278), .C(n_1281), .Y(n_1249) );
OAI21xp33_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1266), .B(n_1277), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_1261), .A2(n_1262), .B1(n_1263), .B2(n_1264), .Y(n_1260) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
OAI21xp5_ASAP7_75t_L g1667 ( .A1(n_1277), .A2(n_1668), .B(n_1679), .Y(n_1667) );
NOR3xp33_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1300), .C(n_1302), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1287), .Y(n_1282) );
BUFx3_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
BUFx2_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVxp67_ASAP7_75t_SL g1448 ( .A(n_1304), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_1305), .A2(n_1354), .B1(n_1446), .B2(n_1447), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx2_ASAP7_75t_L g1446 ( .A(n_1306), .Y(n_1446) );
NOR2x1_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1332), .Y(n_1307) );
A2O1A1Ixp33_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1313), .B(n_1329), .C(n_1330), .Y(n_1308) );
NOR3xp33_ASAP7_75t_SL g1313 ( .A(n_1314), .B(n_1322), .C(n_1323), .Y(n_1313) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1341), .Y(n_1332) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1354), .Y(n_1447) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_1355), .A2(n_1400), .B1(n_1401), .B2(n_1445), .Y(n_1354) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1355), .Y(n_1445) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
XNOR2x1_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
NOR2x1_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1385), .Y(n_1358) );
NAND3xp33_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1379), .C(n_1383), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1378), .Y(n_1360) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1367), .B1(n_1368), .B2(n_1369), .Y(n_1365) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_1388), .A2(n_1411), .B1(n_1438), .B2(n_1442), .Y(n_1437) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
OAI21x1_ASAP7_75t_SL g1402 ( .A1(n_1403), .A2(n_1404), .B(n_1444), .Y(n_1402) );
NAND4xp25_ASAP7_75t_L g1444 ( .A(n_1403), .B(n_1406), .C(n_1408), .D(n_1423), .Y(n_1444) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
NAND3xp33_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1408), .C(n_1423), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1413), .Y(n_1408) );
NAND3xp33_ASAP7_75t_SL g1413 ( .A(n_1414), .B(n_1417), .C(n_1420), .Y(n_1413) );
NAND3xp33_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1429), .C(n_1437), .Y(n_1424) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1431), .B1(n_1434), .B2(n_1435), .Y(n_1429) );
INVx8_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
OAI221xp5_ASAP7_75t_SL g1449 ( .A1(n_1450), .A2(n_1660), .B1(n_1663), .B2(n_1701), .C(n_1707), .Y(n_1449) );
AND5x1_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1616), .C(n_1633), .D(n_1642), .E(n_1653), .Y(n_1450) );
OAI33xp33_ASAP7_75t_L g1451 ( .A1(n_1452), .A2(n_1544), .A3(n_1561), .B1(n_1570), .B2(n_1597), .B3(n_1611), .Y(n_1451) );
OAI211xp5_ASAP7_75t_SL g1452 ( .A1(n_1453), .A2(n_1474), .B(n_1491), .C(n_1534), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g1551 ( .A(n_1453), .Y(n_1551) );
OR2x2_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1469), .Y(n_1453) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_1454), .A2(n_1501), .B1(n_1504), .B2(n_1507), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1454), .B(n_1508), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_1454), .B(n_1470), .Y(n_1543) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1454), .Y(n_1554) );
INVx2_ASAP7_75t_L g1572 ( .A(n_1454), .Y(n_1572) );
OR2x2_ASAP7_75t_L g1586 ( .A(n_1454), .B(n_1510), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1454), .B(n_1509), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1454), .B(n_1510), .Y(n_1641) );
INVx2_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1455), .B(n_1469), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1463), .Y(n_1455) );
INVx2_ASAP7_75t_L g1662 ( .A(n_1457), .Y(n_1662) );
AND2x6_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1459), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1458), .B(n_1462), .Y(n_1461) );
AND2x4_ASAP7_75t_L g1464 ( .A(n_1458), .B(n_1465), .Y(n_1464) );
AND2x6_ASAP7_75t_L g1467 ( .A(n_1458), .B(n_1468), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1458), .B(n_1462), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1458), .B(n_1462), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1458), .B(n_1465), .Y(n_1522) );
OAI21xp5_ASAP7_75t_L g1753 ( .A1(n_1459), .A2(n_1754), .B(n_1755), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1460), .B(n_1466), .Y(n_1465) );
INVx2_ASAP7_75t_L g1524 ( .A(n_1467), .Y(n_1524) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1469), .Y(n_1515) );
NOR2xp33_ASAP7_75t_L g1629 ( .A(n_1469), .B(n_1556), .Y(n_1629) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1470), .Y(n_1508) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1473), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1479), .Y(n_1474) );
NOR2xp33_ASAP7_75t_L g1501 ( .A(n_1475), .B(n_1502), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_1475), .B(n_1537), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1475), .B(n_1551), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g1596 ( .A(n_1475), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1475), .B(n_1505), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1475), .B(n_1518), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1475), .B(n_1515), .Y(n_1645) );
INVx4_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
O2A1O1Ixp33_ASAP7_75t_L g1527 ( .A1(n_1476), .A2(n_1528), .B(n_1530), .C(n_1533), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1476), .B(n_1532), .Y(n_1531) );
INVx4_ASAP7_75t_L g1547 ( .A(n_1476), .Y(n_1547) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1476), .B(n_1550), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1476), .B(n_1497), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1476), .B(n_1545), .Y(n_1555) );
NAND2xp5_ASAP7_75t_SL g1560 ( .A(n_1476), .B(n_1497), .Y(n_1560) );
NOR2xp33_ASAP7_75t_L g1567 ( .A(n_1476), .B(n_1498), .Y(n_1567) );
NOR3xp33_ASAP7_75t_L g1589 ( .A(n_1476), .B(n_1586), .C(n_1590), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1476), .B(n_1539), .Y(n_1640) );
AND2x4_ASAP7_75t_SL g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
NOR2xp33_ASAP7_75t_L g1615 ( .A(n_1479), .B(n_1578), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1483), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1538 ( .A(n_1480), .B(n_1485), .Y(n_1538) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1480), .B(n_1584), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1480), .B(n_1532), .Y(n_1591) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1480), .B(n_1567), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1482), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1481), .B(n_1482), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1607 ( .A(n_1483), .B(n_1496), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1483), .B(n_1655), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1488), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_1485), .B(n_1488), .Y(n_1498) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1485), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1485), .B(n_1488), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1485), .B(n_1506), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1485), .B(n_1497), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1487), .Y(n_1485) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1488), .Y(n_1506) );
NAND2x1p5_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1490), .Y(n_1488) );
AOI211xp5_ASAP7_75t_L g1491 ( .A1(n_1492), .A2(n_1494), .B(n_1499), .C(n_1527), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1492), .B(n_1596), .Y(n_1595) );
CKINVDCx5p33_ASAP7_75t_R g1492 ( .A(n_1493), .Y(n_1492) );
OR2x2_ASAP7_75t_L g1659 ( .A(n_1493), .B(n_1509), .Y(n_1659) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
NOR2xp33_ASAP7_75t_L g1587 ( .A(n_1495), .B(n_1541), .Y(n_1587) );
OR2x2_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1498), .Y(n_1495) );
NOR2xp33_ASAP7_75t_L g1505 ( .A(n_1496), .B(n_1506), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1496), .B(n_1532), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1496), .B(n_1558), .Y(n_1593) );
A2O1A1Ixp33_ASAP7_75t_L g1653 ( .A1(n_1496), .A2(n_1654), .B(n_1656), .C(n_1658), .Y(n_1653) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_1497), .B(n_1503), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1497), .B(n_1518), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1497), .B(n_1503), .Y(n_1529) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1497), .B(n_1506), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1497), .B(n_1506), .Y(n_1626) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1498), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1619 ( .A(n_1498), .B(n_1553), .Y(n_1619) );
OAI221xp5_ASAP7_75t_SL g1499 ( .A1(n_1500), .A2(n_1509), .B1(n_1514), .B2(n_1516), .C(n_1519), .Y(n_1499) );
HB1xp67_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1507), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1533 ( .A(n_1508), .B(n_1509), .Y(n_1533) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1508), .Y(n_1545) );
OAI221xp5_ASAP7_75t_L g1561 ( .A1(n_1508), .A2(n_1554), .B1(n_1562), .B2(n_1566), .C(n_1568), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1508), .B(n_1578), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1508), .B(n_1547), .Y(n_1605) );
A2O1A1Ixp33_ASAP7_75t_L g1633 ( .A1(n_1508), .A2(n_1634), .B(n_1640), .C(n_1641), .Y(n_1633) );
OR2x2_ASAP7_75t_L g1514 ( .A(n_1509), .B(n_1515), .Y(n_1514) );
A2O1A1Ixp33_ASAP7_75t_L g1548 ( .A1(n_1509), .A2(n_1549), .B(n_1551), .C(n_1552), .Y(n_1548) );
CKINVDCx14_ASAP7_75t_R g1610 ( .A(n_1509), .Y(n_1610) );
INVx3_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1510), .Y(n_1542) );
AOI221xp5_ASAP7_75t_L g1616 ( .A1(n_1510), .A2(n_1545), .B1(n_1617), .B2(n_1620), .C(n_1627), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1510), .B(n_1554), .Y(n_1622) );
OAI21xp33_ASAP7_75t_L g1627 ( .A1(n_1510), .A2(n_1628), .B(n_1630), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1512), .Y(n_1510) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1515), .Y(n_1564) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NAND2x1_ASAP7_75t_L g1546 ( .A(n_1517), .B(n_1547), .Y(n_1546) );
OAI21xp33_ASAP7_75t_L g1630 ( .A1(n_1517), .A2(n_1631), .B(n_1632), .Y(n_1630) );
OAI321xp33_ASAP7_75t_L g1552 ( .A1(n_1518), .A2(n_1528), .A3(n_1553), .B1(n_1554), .B2(n_1555), .C(n_1556), .Y(n_1552) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1518), .Y(n_1584) );
OAI21xp5_ASAP7_75t_L g1592 ( .A1(n_1518), .A2(n_1593), .B(n_1594), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1518), .B(n_1559), .Y(n_1624) );
AOI211xp5_ASAP7_75t_L g1601 ( .A1(n_1519), .A2(n_1602), .B(n_1603), .C(n_1604), .Y(n_1601) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1520), .B(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
OAI221xp5_ASAP7_75t_L g1521 ( .A1(n_1522), .A2(n_1523), .B1(n_1524), .B2(n_1525), .C(n_1526), .Y(n_1521) );
NAND2xp5_ASAP7_75t_SL g1582 ( .A(n_1528), .B(n_1583), .Y(n_1582) );
O2A1O1Ixp33_ASAP7_75t_L g1597 ( .A1(n_1528), .A2(n_1598), .B(n_1601), .C(n_1608), .Y(n_1597) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1529), .B(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1532), .Y(n_1655) );
OAI322xp33_ASAP7_75t_L g1611 ( .A1(n_1533), .A2(n_1538), .A3(n_1542), .B1(n_1551), .B2(n_1612), .C1(n_1613), .C2(n_1614), .Y(n_1611) );
OAI21xp33_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1539), .B(n_1540), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
INVxp67_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
NOR2xp33_ASAP7_75t_L g1565 ( .A(n_1538), .B(n_1547), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1539), .B(n_1551), .Y(n_1580) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1539), .Y(n_1650) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
OR2x2_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1543), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1542), .B(n_1645), .Y(n_1644) );
OAI21xp33_ASAP7_75t_L g1544 ( .A1(n_1545), .A2(n_1546), .B(n_1548), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1613 ( .A(n_1545), .B(n_1586), .Y(n_1613) );
CKINVDCx5p33_ASAP7_75t_R g1578 ( .A(n_1547), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1551), .B(n_1596), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1573 ( .A(n_1554), .B(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1554), .Y(n_1602) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
AOI211xp5_ASAP7_75t_L g1571 ( .A1(n_1557), .A2(n_1572), .B(n_1573), .C(n_1579), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1649 ( .A(n_1557), .B(n_1564), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1559), .Y(n_1557) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVxp67_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1564), .B(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
O2A1O1Ixp33_ASAP7_75t_L g1642 ( .A1(n_1569), .A2(n_1643), .B(n_1646), .C(n_1648), .Y(n_1642) );
NAND4xp25_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1581), .C(n_1588), .D(n_1592), .Y(n_1570) );
INVxp33_ASAP7_75t_L g1631 ( .A(n_1574), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1577), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1576), .B(n_1596), .Y(n_1637) );
AOI31xp33_ASAP7_75t_L g1581 ( .A1(n_1578), .A2(n_1582), .A3(n_1585), .B(n_1587), .Y(n_1581) );
NOR2xp33_ASAP7_75t_L g1599 ( .A(n_1578), .B(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
CKINVDCx14_ASAP7_75t_R g1585 ( .A(n_1586), .Y(n_1585) );
OAI22xp5_ASAP7_75t_L g1620 ( .A1(n_1586), .A2(n_1621), .B1(n_1623), .B2(n_1625), .Y(n_1620) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1590), .B(n_1639), .Y(n_1647) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1593), .Y(n_1639) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVxp67_ASAP7_75t_SL g1598 ( .A(n_1599), .Y(n_1598) );
OAI22xp5_ASAP7_75t_L g1648 ( .A1(n_1602), .A2(n_1649), .B1(n_1650), .B2(n_1651), .Y(n_1648) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1603), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
CKINVDCx14_ASAP7_75t_R g1625 ( .A(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1639), .Y(n_1634) );
INVxp67_ASAP7_75t_SL g1635 ( .A(n_1636), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1638), .Y(n_1636) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVxp67_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
CKINVDCx20_ASAP7_75t_R g1660 ( .A(n_1661), .Y(n_1660) );
CKINVDCx20_ASAP7_75t_R g1661 ( .A(n_1662), .Y(n_1661) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
AND4x1_ASAP7_75t_L g1666 ( .A(n_1667), .B(n_1685), .C(n_1696), .D(n_1699), .Y(n_1666) );
INVx2_ASAP7_75t_SL g1672 ( .A(n_1673), .Y(n_1672) );
CKINVDCx20_ASAP7_75t_R g1701 ( .A(n_1702), .Y(n_1701) );
CKINVDCx20_ASAP7_75t_R g1702 ( .A(n_1703), .Y(n_1702) );
INVx3_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
BUFx3_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
HB1xp67_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
BUFx3_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVxp33_ASAP7_75t_SL g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
HB1xp67_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1740), .Y(n_1716) );
HB1xp67_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
endmodule