module real_jpeg_17882_n_20 (n_17, n_8, n_0, n_648, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_648;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_620;
wire n_332;
wire n_366;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_1),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_1),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g446 ( 
.A(n_1),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_3),
.B(n_171),
.Y(n_318)
);

OAI32xp33_ASAP7_75t_L g425 ( 
.A1(n_3),
.A2(n_52),
.A3(n_359),
.B1(n_426),
.B2(n_429),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_3),
.B(n_80),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_3),
.A2(n_84),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_3),
.A2(n_108),
.B1(n_534),
.B2(n_538),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_4),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_4),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_4),
.A2(n_40),
.B1(n_144),
.B2(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_4),
.A2(n_144),
.B1(n_232),
.B2(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_4),
.A2(n_144),
.B1(n_535),
.B2(n_536),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_5),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_5),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_6),
.A2(n_39),
.B1(n_162),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_6),
.A2(n_39),
.B1(n_417),
.B2(n_420),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_6),
.A2(n_39),
.B1(n_462),
.B2(n_465),
.Y(n_461)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_120),
.B1(n_125),
.B2(n_126),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_125),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_7),
.A2(n_125),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_7),
.A2(n_125),
.B1(n_260),
.B2(n_570),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_8),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_8),
.A2(n_193),
.B1(n_385),
.B2(n_389),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_8),
.A2(n_193),
.B1(n_588),
.B2(n_590),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_8),
.A2(n_193),
.B1(n_630),
.B2(n_631),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g314 ( 
.A(n_9),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_10),
.A2(n_165),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_10),
.A2(n_165),
.B1(n_231),
.B2(n_459),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_10),
.A2(n_165),
.B1(n_184),
.B2(n_518),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_12),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_12),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_12),
.A2(n_245),
.B1(n_265),
.B2(n_269),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_12),
.A2(n_245),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_12),
.A2(n_245),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_133),
.B1(n_136),
.B2(n_141),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_13),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_141),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_13),
.A2(n_141),
.B1(n_375),
.B2(n_377),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_13),
.A2(n_141),
.B1(n_570),
.B2(n_583),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_14),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_14),
.A2(n_75),
.B1(n_288),
.B2(n_291),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_14),
.A2(n_75),
.B1(n_350),
.B2(n_353),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_14),
.A2(n_75),
.B1(n_437),
.B2(n_440),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_16),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_16),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_16),
.A2(n_181),
.B1(n_331),
.B2(n_335),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_16),
.A2(n_181),
.B1(n_574),
.B2(n_577),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_16),
.A2(n_181),
.B1(n_619),
.B2(n_620),
.Y(n_618)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_17),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_17),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_17),
.Y(n_237)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_17),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_17),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g164 ( 
.A(n_19),
.Y(n_164)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_19),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_640),
.B(n_644),
.Y(n_24)
);

AO21x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_560),
.B(n_633),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_406),
.B(n_555),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_322),
.C(n_365),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_270),
.B(n_295),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_29),
.B(n_270),
.C(n_557),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_172),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_30),
.B(n_173),
.C(n_238),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_81),
.C(n_142),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_32),
.B(n_142),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_45),
.B1(n_70),
.B2(n_79),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_34),
.A2(n_80),
.B1(n_278),
.B2(n_282),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_45),
.A2(n_70),
.B1(n_79),
.B2(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_45),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_45),
.A2(n_79),
.B1(n_264),
.B2(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_45),
.A2(n_79),
.B1(n_303),
.B2(n_478),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_45),
.A2(n_79),
.B1(n_374),
.B2(n_573),
.Y(n_572)
);

OAI22x1_ASAP7_75t_SL g586 ( 
.A1(n_45),
.A2(n_79),
.B1(n_573),
.B2(n_587),
.Y(n_586)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_52),
.B(n_57),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_55),
.Y(n_589)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.Y(n_57)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_58),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_59),
.Y(n_211)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_59),
.Y(n_248)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_60),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_60),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_60),
.Y(n_510)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_74),
.Y(n_360)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_74),
.Y(n_381)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_74),
.Y(n_593)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_77),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_77),
.Y(n_281)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_80),
.A2(n_278),
.B1(n_282),
.B2(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_80),
.A2(n_282),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_80),
.A2(n_282),
.B(n_615),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_81),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_107),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_82),
.B(n_107),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_89),
.B1(n_96),
.B2(n_102),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_SL g284 ( 
.A1(n_83),
.A2(n_84),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_84),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_84),
.B(n_499),
.Y(n_498)
);

OAI21xp33_ASAP7_75t_SL g507 ( 
.A1(n_84),
.A2(n_498),
.B(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_84),
.B(n_530),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_84),
.B(n_197),
.Y(n_542)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_88),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_100),
.Y(n_268)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_101),
.Y(n_307)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_101),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_149),
.B(n_154),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_104),
.Y(n_401)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_118),
.B1(n_130),
.B2(n_132),
.Y(n_107)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_108),
.A2(n_132),
.B1(n_177),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_108),
.A2(n_190),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_108),
.A2(n_461),
.B1(n_467),
.B2(n_469),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_108),
.A2(n_342),
.B1(n_517),
.B2(n_534),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_111),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_112),
.Y(n_344)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_119),
.A2(n_175),
.B1(n_309),
.B2(n_315),
.Y(n_308)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_124),
.Y(n_520)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_127),
.Y(n_191)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_128),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_131),
.Y(n_468)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_140),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_148),
.B1(n_160),
.B2(n_171),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_143),
.A2(n_148),
.B1(n_171),
.B2(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_148),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_148),
.A2(n_171),
.B1(n_581),
.B2(n_582),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_148),
.A2(n_171),
.B(n_642),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_161),
.A2(n_256),
.B1(n_257),
.B2(n_262),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_164),
.Y(n_285)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_169),
.Y(n_352)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_169),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_170),
.Y(n_399)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_238),
.Y(n_172)
);

XNOR2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_194),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_174),
.A2(n_195),
.B(n_218),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_186),
.B2(n_189),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_175),
.A2(n_309),
.B1(n_436),
.B2(n_443),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_175),
.A2(n_516),
.B1(n_521),
.B2(n_522),
.Y(n_515)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_180),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_180),
.Y(n_535)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_188),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_218),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_208),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_196),
.A2(n_219),
.B1(n_287),
.B2(n_294),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_196),
.A2(n_219),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_196),
.A2(n_219),
.B1(n_453),
.B2(n_458),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_196),
.A2(n_219),
.B1(n_416),
.B2(n_458),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_196),
.A2(n_219),
.B1(n_453),
.B2(n_507),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g566 ( 
.A1(n_196),
.A2(n_219),
.B(n_384),
.Y(n_566)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_197),
.A2(n_229),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_197),
.A2(n_209),
.B1(n_241),
.B2(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_197),
.A2(n_241),
.B1(n_415),
.B2(n_422),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_202),
.Y(n_439)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_217),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_228),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_219),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_225),
.B2(n_227),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_225),
.Y(n_497)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_226),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_227),
.Y(n_230)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_227),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_236),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_236),
.Y(n_428)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_254),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_239),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_249),
.Y(n_239)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_263),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

OAI22x1_ASAP7_75t_L g348 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_349),
.Y(n_348)
);

OAI22x1_ASAP7_75t_L g395 ( 
.A1(n_256),
.A2(n_262),
.B1(n_349),
.B2(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_256),
.A2(n_262),
.B1(n_396),
.B2(n_569),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_256),
.A2(n_262),
.B1(n_617),
.B2(n_618),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_256),
.A2(n_262),
.B1(n_618),
.B2(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_263),
.B(n_325),
.C(n_326),
.Y(n_324)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_267),
.Y(n_577)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_275),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_271),
.A2(n_272),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_276),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.C(n_286),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_286),
.Y(n_298)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_279),
.Y(n_357)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_280),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_280),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_285),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_287),
.Y(n_422)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_288),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_319),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_296),
.B(n_319),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_297),
.B(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_299),
.B(n_300),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.C(n_318),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_301),
.B(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_308),
.B(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_310),
.Y(n_466)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_313),
.Y(n_464)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_314),
.Y(n_442)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_314),
.Y(n_504)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

A2O1A1O1Ixp25_ASAP7_75t_L g555 ( 
.A1(n_322),
.A2(n_365),
.B(n_556),
.C(n_558),
.D(n_559),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_364),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_323),
.B(n_364),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_346),
.B1(n_362),
.B2(n_363),
.Y(n_327)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_328),
.B(n_363),
.C(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_340),
.B1(n_341),
.B2(n_345),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_329),
.B(n_341),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_334),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_340),
.A2(n_341),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_340),
.A2(n_395),
.B1(n_403),
.B2(n_648),
.Y(n_603)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_361),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_361),
.C(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_353),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_404),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_366),
.B(n_404),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_367),
.B(n_606),
.C(n_607),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_391),
.Y(n_369)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_370),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_382),
.B(n_390),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_382),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_380),
.Y(n_576)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_387),
.Y(n_499)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_390),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_390),
.A2(n_599),
.B1(n_602),
.B2(n_610),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_391),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_402),
.B2(n_403),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_398),
.Y(n_631)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_401),
.Y(n_630)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_402),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_447),
.B(n_554),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_408),
.B(n_410),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_414),
.C(n_423),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_411),
.A2(n_412),
.B1(n_549),
.B2(n_550),
.Y(n_548)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_414),
.A2(n_423),
.B1(n_424),
.B2(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_414),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_434),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_425),
.A2(n_434),
.B1(n_435),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_425),
.Y(n_474)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_437),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_547),
.B(n_553),
.Y(n_447)
);

AOI21x1_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_485),
.B(n_546),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_472),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_450),
.B(n_472),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_460),
.C(n_470),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_451),
.A2(n_452),
.B1(n_470),
.B2(n_471),
.Y(n_512)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_460),
.B(n_512),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_467),
.Y(n_521)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_473),
.B(n_476),
.C(n_484),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_483),
.B2(n_484),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_513),
.B(n_545),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_511),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_487),
.B(n_511),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_505),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_488),
.A2(n_505),
.B1(n_506),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

OAI32xp33_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_491),
.A3(n_495),
.B1(n_498),
.B2(n_500),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_525),
.B(n_544),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_523),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_515),
.B(n_523),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_540),
.B(n_543),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_533),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_542),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_542),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g547 ( 
.A(n_548),
.B(n_552),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_552),
.Y(n_553)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_611),
.C(n_626),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_604),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_563),
.A2(n_636),
.B(n_637),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_SL g563 ( 
.A(n_564),
.B(n_598),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_564),
.B(n_598),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_578),
.Y(n_564)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_567),
.C(n_571),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_566),
.A2(n_586),
.B1(n_594),
.B2(n_595),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_566),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_566),
.B(n_572),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_580),
.C(n_595),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_567),
.A2(n_579),
.B1(n_596),
.B2(n_597),
.Y(n_578)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_567),
.A2(n_568),
.B1(n_600),
.B2(n_601),
.Y(n_599)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_569),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_579),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_579),
.B(n_596),
.C(n_625),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_585),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_583),
.Y(n_619)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_586),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_587),
.Y(n_615)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_602),
.C(n_603),
.Y(n_598)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_599),
.Y(n_610)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_600),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_603),
.B(n_609),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_608),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_605),
.B(n_608),
.Y(n_636)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

A2O1A1O1Ixp25_ASAP7_75t_L g634 ( 
.A1(n_612),
.A2(n_627),
.B(n_635),
.C(n_638),
.D(n_639),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_624),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_613),
.B(n_624),
.Y(n_638)
);

BUFx24_ASAP7_75t_SL g647 ( 
.A(n_613),
.Y(n_647)
);

FAx1_ASAP7_75t_SL g613 ( 
.A(n_614),
.B(n_616),
.CI(n_623),
.CON(n_613),
.SN(n_613)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_616),
.C(n_623),
.Y(n_632)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_628),
.B(n_632),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_632),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_641),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_641),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_629),
.Y(n_643)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g642 ( 
.A(n_643),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_645),
.Y(n_644)
);


endmodule