module fake_jpeg_9755_n_144 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_51),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_26),
.Y(n_59)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_67),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_38),
.C(n_18),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_63),
.Y(n_85)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_69),
.B1(n_45),
.B2(n_19),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_65),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_38),
.C(n_18),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_28),
.B1(n_29),
.B2(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_70),
.B1(n_25),
.B2(n_23),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_16),
.B1(n_20),
.B2(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_24),
.B1(n_20),
.B2(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_76),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_48),
.B1(n_53),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_53),
.B1(n_43),
.B2(n_25),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_87),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_86),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_58),
.B(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_55),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_1),
.C(n_2),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_63),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_96),
.C(n_74),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_57),
.B(n_64),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

XOR2x1_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_61),
.C(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_3),
.C(n_4),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_112),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_88),
.B(n_82),
.C(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_100),
.C(n_73),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_93),
.B(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_23),
.B1(n_81),
.B2(n_5),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_95),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_91),
.C(n_103),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_120),
.B(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_131)
);

XOR2x2_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_106),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_118),
.B1(n_122),
.B2(n_109),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_124),
.B(n_3),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.C(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_81),
.C(n_73),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_66),
.C(n_7),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_11),
.B(n_13),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_7),
.C(n_9),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_4),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_130),
.C(n_134),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_66),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_140),
.Y(n_144)
);


endmodule