module fake_aes_12517_n_724 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_724);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_724;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g108 ( .A(n_105), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_60), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_53), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_102), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_95), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_10), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_96), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_52), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_25), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_20), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_11), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_5), .B(n_85), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_97), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_9), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_33), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_9), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_45), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_61), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_35), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_87), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_59), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_38), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_0), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_30), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_37), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_29), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_84), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_76), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_24), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_70), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_68), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_79), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_47), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_43), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_73), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_2), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_148), .A2(n_48), .B(n_106), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_148), .B(n_0), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_148), .B(n_1), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_126), .B(n_1), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_109), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g160 ( .A1(n_121), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_128), .B(n_3), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_131), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_109), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_110), .B(n_27), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_119), .B(n_4), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_119), .B(n_5), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_113), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_120), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_112), .B(n_6), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_155), .B(n_120), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_158), .B(n_127), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_153), .B(n_127), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_169), .B(n_124), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_164), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_155), .A2(n_137), .B1(n_150), .B2(n_130), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_153), .B(n_149), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_164), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_153), .B(n_149), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_155), .Y(n_184) );
BUFx10_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_159), .B(n_113), .Y(n_186) );
INVx4_ASAP7_75t_SL g187 ( .A(n_156), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_159), .B(n_114), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_159), .B(n_114), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_164), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_156), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_163), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_187), .B(n_161), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_198), .B(n_163), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_182), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_178), .Y(n_202) );
NOR2x2_ASAP7_75t_L g203 ( .A(n_179), .B(n_162), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_187), .B(n_161), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_187), .B(n_172), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_198), .B(n_163), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
AND2x6_ASAP7_75t_SL g209 ( .A(n_176), .B(n_157), .Y(n_209) );
OR2x4_ASAP7_75t_L g210 ( .A(n_174), .B(n_167), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_187), .B(n_172), .Y(n_211) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_185), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_192), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_192), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_176), .B(n_169), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_185), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_194), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_179), .A2(n_172), .B1(n_166), .B2(n_157), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_173), .A2(n_168), .B(n_158), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_192), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_187), .B(n_172), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_198), .B(n_168), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_185), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_176), .Y(n_225) );
INVxp67_ASAP7_75t_L g226 ( .A(n_186), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_179), .A2(n_172), .B1(n_166), .B2(n_157), .Y(n_227) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_177), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_179), .A2(n_172), .B1(n_166), .B2(n_168), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_194), .B(n_162), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_191), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_187), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_202), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_212), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_202), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_226), .B(n_177), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_212), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_216), .B(n_184), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_201), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_225), .B(n_194), .Y(n_241) );
O2A1O1Ixp5_ASAP7_75t_L g242 ( .A1(n_206), .A2(n_173), .B(n_188), .C(n_174), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_200), .A2(n_197), .B(n_195), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_211), .A2(n_197), .B(n_195), .C(n_186), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_219), .A2(n_179), .B1(n_196), .B2(n_184), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_190), .B(n_189), .C(n_167), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_200), .A2(n_188), .B(n_196), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_212), .B(n_185), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_218), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_202), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_218), .B(n_194), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_201), .Y(n_253) );
OAI21xp33_ASAP7_75t_L g254 ( .A1(n_230), .A2(n_179), .B(n_177), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_220), .A2(n_188), .B(n_180), .C(n_177), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_219), .A2(n_196), .B1(n_194), .B2(n_180), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_210), .B(n_115), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
OAI22x1_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_165), .B1(n_160), .B2(n_140), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_210), .B(n_180), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_227), .B(n_185), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
AOI221x1_ASAP7_75t_L g263 ( .A1(n_220), .A2(n_171), .B1(n_142), .B2(n_135), .C(n_144), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_229), .B(n_180), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_240), .Y(n_265) );
INVxp33_ASAP7_75t_L g266 ( .A(n_257), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_246), .B(n_232), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_238), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_238), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_254), .A2(n_189), .B1(n_190), .B2(n_181), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_254), .A2(n_188), .B1(n_232), .B2(n_231), .Y(n_273) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_255), .A2(n_154), .B(n_171), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_253), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g277 ( .A1(n_239), .A2(n_207), .B(n_223), .C(n_181), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_263), .A2(n_154), .B(n_165), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_263), .B(n_175), .C(n_183), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_262), .A2(n_154), .B(n_171), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_238), .Y(n_282) );
CKINVDCx11_ASAP7_75t_R g283 ( .A(n_243), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_248), .A2(n_207), .B(n_223), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_259), .A2(n_210), .B1(n_160), .B2(n_133), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_243), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_272), .A2(n_236), .B(n_234), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_268), .B(n_261), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_266), .A2(n_259), .B1(n_261), .B2(n_260), .Y(n_292) );
AOI221xp5_ASAP7_75t_SL g293 ( .A1(n_277), .A2(n_247), .B1(n_245), .B2(n_244), .C(n_183), .Y(n_293) );
NOR2x1_ASAP7_75t_L g294 ( .A(n_277), .B(n_234), .Y(n_294) );
AOI21xp33_ASAP7_75t_L g295 ( .A1(n_272), .A2(n_273), .B(n_268), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_256), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_265), .B(n_235), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_267), .B(n_256), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_266), .A2(n_237), .B1(n_243), .B2(n_235), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_285), .A2(n_237), .B1(n_243), .B2(n_241), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_267), .B(n_236), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g302 ( .A1(n_285), .A2(n_203), .B1(n_165), .B2(n_251), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_273), .A2(n_242), .B(n_237), .C(n_264), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_275), .A2(n_264), .B1(n_250), .B2(n_258), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_275), .A2(n_276), .B1(n_287), .B2(n_283), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_276), .B(n_251), .Y(n_306) );
AOI22xp33_ASAP7_75t_SL g307 ( .A1(n_287), .A2(n_165), .B1(n_209), .B2(n_118), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_284), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_308), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_310), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_291), .B(n_274), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_301), .B(n_271), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
CKINVDCx14_ASAP7_75t_R g318 ( .A(n_298), .Y(n_318) );
BUFx6f_ASAP7_75t_SL g319 ( .A(n_297), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_291), .B(n_282), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_310), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_291), .B(n_269), .Y(n_322) );
AO31x2_ASAP7_75t_L g323 ( .A1(n_309), .A2(n_288), .A3(n_282), .B(n_175), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_301), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_306), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_306), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_309), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_310), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_298), .B(n_288), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_298), .B(n_288), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_308), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_296), .B(n_269), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_296), .B(n_274), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_295), .B(n_270), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_295), .B(n_274), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_314), .B(n_274), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_333), .B(n_292), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_333), .B(n_302), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_327), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_314), .B(n_274), .Y(n_343) );
AOI22xp33_ASAP7_75t_SL g344 ( .A1(n_318), .A2(n_302), .B1(n_297), .B2(n_307), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_321), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_324), .B(n_209), .Y(n_346) );
OAI33xp33_ASAP7_75t_L g347 ( .A1(n_311), .A2(n_140), .A3(n_134), .B1(n_152), .B2(n_143), .B3(n_147), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_314), .B(n_289), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_334), .B(n_289), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_321), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_319), .A2(n_297), .B1(n_307), .B2(n_270), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_328), .A2(n_284), .B(n_278), .Y(n_357) );
OAI31xp33_ASAP7_75t_L g358 ( .A1(n_325), .A2(n_300), .A3(n_305), .B(n_297), .Y(n_358) );
INVx5_ASAP7_75t_SL g359 ( .A(n_316), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_320), .A2(n_280), .B1(n_286), .B2(n_271), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_328), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_334), .B(n_271), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_334), .B(n_281), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_337), .B(n_281), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_337), .B(n_281), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_315), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_337), .B(n_281), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_325), .B(n_303), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_323), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_326), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_326), .B(n_271), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_329), .B(n_281), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_313), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_329), .B(n_165), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_313), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_323), .Y(n_380) );
NOR2x1p5_ASAP7_75t_L g381 ( .A(n_317), .B(n_286), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_341), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_341), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_376), .B(n_332), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_344), .B(n_331), .C(n_336), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_376), .B(n_332), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_376), .B(n_332), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_363), .B(n_330), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_345), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_347), .B(n_143), .C(n_134), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_368), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_368), .B(n_324), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_363), .B(n_330), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_365), .B(n_323), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_365), .B(n_323), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_363), .B(n_336), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_338), .B(n_317), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_338), .B(n_317), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_369), .B(n_331), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_373), .B(n_317), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_354), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_338), .B(n_343), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_344), .A2(n_280), .B(n_125), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_350), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_346), .B(n_152), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_343), .B(n_335), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_343), .B(n_335), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_373), .B(n_322), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_354), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_354), .Y(n_419) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_362), .B(n_316), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_351), .A2(n_136), .B(n_150), .Y(n_421) );
OAI33xp33_ASAP7_75t_L g422 ( .A1(n_339), .A2(n_138), .A3(n_116), .B1(n_147), .B2(n_146), .B3(n_144), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_372), .B(n_374), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_349), .B(n_316), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_339), .B(n_322), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_347), .B(n_112), .C(n_136), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_349), .B(n_316), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_366), .B(n_320), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_366), .B(n_313), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_349), .B(n_313), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_350), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_348), .B(n_366), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_348), .B(n_313), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_367), .B(n_313), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_367), .B(n_116), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_351), .B(n_6), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_372), .B(n_130), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_353), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_381), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_353), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_362), .Y(n_441) );
OR2x6_ASAP7_75t_L g442 ( .A(n_381), .B(n_319), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_367), .B(n_135), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_340), .B(n_7), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_375), .B(n_319), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_340), .A2(n_319), .B1(n_299), .B2(n_304), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_348), .B(n_137), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_353), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_418), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_395), .B(n_362), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_395), .B(n_362), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_447), .B(n_370), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_387), .A2(n_359), .B1(n_380), .B2(n_374), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_447), .B(n_370), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_388), .B(n_380), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_359), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_432), .B(n_370), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_428), .B(n_361), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_435), .B(n_356), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_382), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_387), .A2(n_358), .B(n_139), .C(n_138), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_432), .B(n_361), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_400), .B(n_359), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_382), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_441), .B(n_379), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_410), .B(n_364), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_403), .B(n_364), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_443), .B(n_371), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_442), .B(n_375), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_383), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_383), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_385), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_424), .B(n_427), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_424), .B(n_359), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_384), .B(n_379), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
NAND2x1_ASAP7_75t_L g479 ( .A(n_442), .B(n_364), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_419), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_385), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_427), .B(n_359), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_414), .B(n_371), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_389), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_389), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_386), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_390), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_414), .B(n_378), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_390), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_403), .B(n_359), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_386), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_391), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_410), .B(n_384), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_394), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_444), .B(n_7), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_415), .B(n_378), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_415), .B(n_378), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_404), .B(n_379), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_413), .A2(n_139), .B(n_142), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_391), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_398), .Y(n_502) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_437), .B(n_379), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_420), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_392), .B(n_377), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_398), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_394), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_406), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_396), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_406), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_425), .B(n_358), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_436), .B(n_146), .C(n_122), .D(n_170), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_396), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_407), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_417), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_392), .B(n_377), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_404), .B(n_377), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_422), .A2(n_360), .B(n_357), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_405), .B(n_357), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_416), .B(n_8), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_393), .B(n_8), .Y(n_521) );
OA211x2_ASAP7_75t_L g522 ( .A1(n_421), .A2(n_283), .B(n_11), .C(n_12), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_393), .B(n_10), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g524 ( .A1(n_445), .A2(n_170), .B(n_193), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_401), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_405), .B(n_12), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_399), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_417), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_437), .B(n_13), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_408), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_412), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_478), .B(n_401), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_449), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_524), .A2(n_442), .B1(n_439), .B2(n_445), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_511), .A2(n_439), .B1(n_411), .B2(n_397), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_525), .A2(n_402), .B(n_429), .Y(n_536) );
NAND2x2_ASAP7_75t_L g537 ( .A(n_479), .B(n_402), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_478), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_480), .B(n_433), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_480), .B(n_433), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_481), .B(n_442), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_462), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_513), .Y(n_543) );
OAI31xp33_ASAP7_75t_L g544 ( .A1(n_496), .A2(n_445), .A3(n_420), .B(n_426), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_513), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_496), .A2(n_446), .B1(n_430), .B2(n_434), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_464), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_463), .A2(n_430), .B(n_412), .C(n_438), .Y(n_548) );
AOI32xp33_ASAP7_75t_L g549 ( .A1(n_523), .A2(n_448), .A3(n_438), .B1(n_440), .B2(n_431), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_504), .A2(n_448), .B1(n_440), .B2(n_431), .Y(n_550) );
INVxp33_ASAP7_75t_L g551 ( .A(n_523), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_466), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_472), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_530), .B(n_14), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_482), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_471), .A2(n_170), .B(n_278), .C(n_286), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
OAI21xp33_ASAP7_75t_SL g560 ( .A1(n_494), .A2(n_278), .B(n_170), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_486), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_488), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_522), .A2(n_286), .B1(n_279), .B2(n_170), .Y(n_563) );
NAND2xp33_ASAP7_75t_R g564 ( .A(n_464), .B(n_14), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_490), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_500), .A2(n_293), .B(n_193), .C(n_279), .Y(n_567) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_457), .B(n_279), .Y(n_568) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_450), .B(n_15), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_477), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g571 ( .A1(n_454), .A2(n_279), .B(n_16), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_501), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_526), .A2(n_279), .B1(n_249), .B2(n_193), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_453), .Y(n_574) );
O2A1O1Ixp5_ASAP7_75t_L g575 ( .A1(n_456), .A2(n_193), .B(n_191), .C(n_199), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_520), .B(n_293), .C(n_279), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_456), .B(n_15), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_502), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_506), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_494), .B(n_16), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_487), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_453), .Y(n_582) );
AOI21xp5_ASAP7_75t_SL g583 ( .A1(n_461), .A2(n_279), .B(n_18), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_477), .Y(n_584) );
AOI32xp33_ASAP7_75t_L g585 ( .A1(n_465), .A2(n_17), .A3(n_18), .B1(n_19), .B2(n_20), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_477), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_458), .B(n_17), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_481), .B(n_19), .Y(n_588) );
AOI32xp33_ASAP7_75t_L g589 ( .A1(n_451), .A2(n_21), .A3(n_22), .B1(n_23), .B2(n_24), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_503), .A2(n_145), .B1(n_117), .B2(n_123), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_525), .A2(n_111), .B(n_129), .C(n_132), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_458), .B(n_21), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_512), .A2(n_151), .B1(n_141), .B2(n_205), .C(n_26), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_475), .B(n_22), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_468), .B(n_23), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_503), .A2(n_250), .B1(n_26), .B2(n_258), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_527), .A2(n_188), .B1(n_258), .B2(n_250), .C(n_215), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_491), .A2(n_252), .B1(n_228), .B2(n_204), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_519), .A2(n_215), .B1(n_208), .B2(n_221), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_461), .A2(n_221), .B(n_215), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_484), .A2(n_221), .B(n_214), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_468), .B(n_31), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_508), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_510), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_469), .B(n_214), .Y(n_605) );
INVxp33_ASAP7_75t_L g606 ( .A(n_521), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_470), .A2(n_214), .B1(n_208), .B2(n_204), .C(n_252), .Y(n_607) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_529), .A2(n_32), .B(n_34), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_514), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_571), .A2(n_518), .B(n_460), .C(n_498), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_537), .A2(n_483), .B1(n_476), .B2(n_452), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_538), .B(n_489), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_609), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g614 ( .A1(n_571), .A2(n_459), .B(n_455), .C(n_497), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_570), .B(n_499), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_564), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_574), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_542), .Y(n_618) );
OAI31xp33_ASAP7_75t_L g619 ( .A1(n_544), .A2(n_467), .A3(n_516), .B(n_531), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_552), .Y(n_620) );
INVxp33_ASAP7_75t_L g621 ( .A(n_569), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_533), .B(n_505), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_549), .B(n_516), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_554), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_534), .A2(n_528), .B1(n_487), .B2(n_515), .Y(n_626) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_580), .B(n_517), .Y(n_627) );
AO22x2_ASAP7_75t_L g628 ( .A1(n_574), .A2(n_467), .B1(n_515), .B2(n_509), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_532), .B(n_528), .Y(n_629) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_594), .Y(n_630) );
OA22x2_ASAP7_75t_L g631 ( .A1(n_546), .A2(n_467), .B1(n_507), .B2(n_495), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_556), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_535), .A2(n_509), .B1(n_507), .B2(n_495), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_557), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_559), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_583), .A2(n_492), .B(n_204), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_547), .B(n_492), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_561), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_570), .B(n_584), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g640 ( .A(n_587), .B(n_36), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_584), .B(n_39), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_596), .B(n_208), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_551), .A2(n_252), .B1(n_233), .B2(n_218), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_543), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_562), .Y(n_645) );
NAND2x1_ASAP7_75t_L g646 ( .A(n_586), .B(n_40), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_586), .B(n_41), .Y(n_647) );
NOR2x1_ASAP7_75t_L g648 ( .A(n_596), .B(n_42), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_565), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_545), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_588), .A2(n_224), .B(n_217), .C(n_213), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_539), .B(n_44), .Y(n_653) );
AO22x1_ASAP7_75t_L g654 ( .A1(n_541), .A2(n_46), .B1(n_49), .B2(n_50), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_572), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_578), .Y(n_656) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_536), .A2(n_51), .B(n_54), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_579), .B(n_55), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_582), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_606), .B(n_56), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_618), .B(n_603), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_616), .A2(n_544), .B(n_548), .Y(n_663) );
AOI21xp33_ASAP7_75t_SL g664 ( .A1(n_631), .A2(n_585), .B(n_589), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_629), .B(n_540), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_619), .A2(n_563), .B(n_592), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_620), .B(n_604), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_659), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_614), .A2(n_633), .B1(n_611), .B2(n_624), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_621), .A2(n_577), .B(n_555), .C(n_593), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_614), .A2(n_595), .B1(n_568), .B2(n_550), .Y(n_671) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_626), .A2(n_576), .B1(n_573), .B2(n_560), .C1(n_602), .C2(n_601), .Y(n_672) );
OAI21xp33_ASAP7_75t_L g673 ( .A1(n_631), .A2(n_599), .B(n_576), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_630), .A2(n_573), .B1(n_600), .B2(n_598), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_648), .A2(n_590), .B1(n_607), .B2(n_581), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_610), .A2(n_558), .B(n_575), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_619), .B(n_605), .Y(n_677) );
XNOR2x1_ASAP7_75t_L g678 ( .A(n_627), .B(n_590), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_628), .A2(n_597), .B1(n_608), .B2(n_567), .C(n_591), .Y(n_679) );
XOR2x2_ASAP7_75t_L g680 ( .A(n_640), .B(n_57), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_646), .A2(n_62), .B(n_63), .C(n_64), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_622), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_617), .A2(n_642), .B1(n_612), .B2(n_657), .C(n_613), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_623), .B(n_69), .Y(n_684) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_617), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_639), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_660), .A2(n_71), .B1(n_72), .B2(n_74), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_643), .A2(n_75), .B1(n_77), .B2(n_80), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_664), .A2(n_628), .B1(n_656), .B2(n_655), .C(n_625), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_663), .A2(n_632), .B1(n_634), .B2(n_635), .C(n_650), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_662), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_669), .A2(n_645), .B1(n_638), .B2(n_649), .Y(n_692) );
AOI221x1_ASAP7_75t_L g693 ( .A1(n_673), .A2(n_658), .B1(n_636), .B2(n_647), .C(n_641), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_668), .Y(n_694) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_672), .A2(n_652), .B(n_653), .C(n_658), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_677), .A2(n_637), .B1(n_651), .B2(n_644), .C(n_615), .Y(n_696) );
AOI211x1_ASAP7_75t_SL g697 ( .A1(n_676), .A2(n_654), .B(n_83), .C(n_86), .Y(n_697) );
NOR4xp25_ASAP7_75t_L g698 ( .A(n_670), .B(n_685), .C(n_666), .D(n_683), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_671), .A2(n_81), .B1(n_88), .B2(n_90), .C(n_91), .Y(n_699) );
AOI21xp33_ASAP7_75t_SL g700 ( .A1(n_678), .A2(n_92), .B(n_94), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g701 ( .A(n_679), .B(n_99), .C(n_100), .D(n_101), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_661), .A2(n_103), .B1(n_104), .B2(n_107), .C(n_213), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_691), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_694), .Y(n_704) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_701), .B(n_681), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_689), .A2(n_680), .B1(n_661), .B2(n_667), .C1(n_686), .C2(n_684), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_692), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_696), .B(n_665), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_698), .A2(n_667), .B1(n_674), .B2(n_675), .C(n_688), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_704), .B(n_700), .Y(n_710) );
AOI32xp33_ASAP7_75t_L g711 ( .A1(n_709), .A2(n_695), .A3(n_690), .B1(n_699), .B2(n_693), .Y(n_711) );
INVx2_ASAP7_75t_SL g712 ( .A(n_703), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_707), .B(n_702), .C(n_682), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_713), .B(n_708), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_710), .Y(n_716) );
OAI22x1_ASAP7_75t_L g717 ( .A1(n_714), .A2(n_705), .B1(n_711), .B2(n_706), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_716), .Y(n_718) );
XOR2x2_ASAP7_75t_L g719 ( .A(n_718), .B(n_715), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_717), .Y(n_720) );
OA21x2_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_706), .B(n_687), .Y(n_721) );
AOI22xp33_ASAP7_75t_R g722 ( .A1(n_719), .A2(n_697), .B1(n_217), .B2(n_224), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_721), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_721), .B(n_722), .Y(n_724) );
endmodule