module fake_jpeg_29365_n_12 (n_3, n_2, n_1, n_0, n_4, n_12);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_12;

wire n_11;
wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

CKINVDCx14_ASAP7_75t_R g5 ( 
.A(n_4),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_SL g6 ( 
.A(n_2),
.B(n_3),
.Y(n_6)
);

INVx13_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_0),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_L g10 ( 
.A1(n_6),
.A2(n_1),
.B1(n_3),
.B2(n_8),
.Y(n_10)
);

FAx1_ASAP7_75t_R g12 ( 
.A(n_10),
.B(n_11),
.CI(n_7),
.CON(n_12),
.SN(n_12)
);

AOI321xp33_ASAP7_75t_L g11 ( 
.A1(n_6),
.A2(n_9),
.A3(n_5),
.B1(n_7),
.B2(n_3),
.C(n_0),
.Y(n_11)
);


endmodule