module fake_jpeg_19903_n_356 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_36),
.B(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_0),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_54),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_61),
.A2(n_64),
.B1(n_83),
.B2(n_0),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_36),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_68),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_75),
.B1(n_82),
.B2(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_19),
.B(n_18),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_19),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_26),
.B1(n_34),
.B2(n_20),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_34),
.B1(n_21),
.B2(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_108),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_92),
.B(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_40),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_38),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_104),
.B(n_97),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_104),
.B(n_48),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_37),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_107),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_46),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_17),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_54),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_121),
.C(n_19),
.Y(n_144)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_35),
.B(n_21),
.Y(n_104)
);

OR2x4_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_35),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_37),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_52),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_52),
.B1(n_23),
.B2(n_27),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_120),
.B1(n_127),
.B2(n_59),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_113),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_64),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_19),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_57),
.A2(n_48),
.B1(n_16),
.B2(n_17),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_18),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_107),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_63),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_59),
.B1(n_76),
.B2(n_27),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_78),
.B1(n_79),
.B2(n_71),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_19),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_131),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_60),
.B1(n_70),
.B2(n_72),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_133),
.A2(n_146),
.B1(n_156),
.B2(n_157),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_139),
.B1(n_155),
.B2(n_94),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_85),
.B1(n_59),
.B2(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_141),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_11),
.B(n_10),
.C(n_12),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_153),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_159),
.B(n_1),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

OR2x4_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_120),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_103),
.A2(n_76),
.B1(n_27),
.B2(n_23),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_23),
.B1(n_17),
.B2(n_63),
.Y(n_157)
);

NAND2x1_ASAP7_75t_SL g159 ( 
.A(n_100),
.B(n_0),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_93),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_168),
.B1(n_192),
.B2(n_131),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_100),
.C(n_89),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_175),
.C(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_167),
.B(n_181),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_90),
.B1(n_98),
.B2(n_126),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_129),
.B(n_148),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_178),
.B(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_99),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_186),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_99),
.C(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_141),
.CON(n_208),
.SN(n_208)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_101),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_117),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_119),
.Y(n_212)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_189),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_129),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_134),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_191),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_145),
.A2(n_122),
.B1(n_109),
.B2(n_95),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_138),
.B1(n_155),
.B2(n_139),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_209),
.B1(n_211),
.B2(n_218),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_11),
.C(n_12),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_166),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_213),
.B(n_4),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_175),
.B1(n_171),
.B2(n_190),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_150),
.B1(n_143),
.B2(n_152),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_164),
.A2(n_153),
.B1(n_130),
.B2(n_105),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_176),
.B1(n_186),
.B2(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_130),
.B1(n_118),
.B2(n_105),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_136),
.B(n_3),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_102),
.B1(n_136),
.B2(n_9),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_192),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_2),
.B(n_3),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_216),
.B(n_227),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_102),
.B(n_119),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_225),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_161),
.B1(n_170),
.B2(n_172),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_166),
.A2(n_2),
.B(n_4),
.Y(n_227)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_240),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_232),
.A2(n_241),
.B(n_198),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_233),
.B(n_235),
.Y(n_269)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_174),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_243),
.Y(n_261)
);

OAI22x1_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_178),
.B1(n_190),
.B2(n_168),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_246),
.B1(n_252),
.B2(n_213),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_165),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_179),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_211),
.B1(n_202),
.B2(n_217),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_176),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_193),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_179),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_226),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_200),
.B(n_205),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_183),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_227),
.C(n_214),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_219),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_224),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_253),
.A2(n_256),
.B(n_5),
.C(n_7),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_199),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_215),
.B1(n_221),
.B2(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_255),
.Y(n_271)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_197),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_262),
.C(n_268),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_218),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_263),
.B(n_231),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_259),
.B(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_210),
.C(n_202),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_216),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_265),
.A2(n_272),
.B1(n_246),
.B2(n_254),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_263),
.B1(n_258),
.B2(n_230),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_224),
.C(n_220),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_230),
.A2(n_220),
.B1(n_217),
.B2(n_206),
.Y(n_272)
);

O2A1O1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_267),
.B(n_253),
.C(n_270),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_277),
.B1(n_236),
.B2(n_240),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_200),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_247),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_296),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_233),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_293),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_287),
.B1(n_292),
.B2(n_265),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_255),
.B(n_231),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_288),
.A2(n_273),
.B(n_249),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_297),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_237),
.B1(n_235),
.B2(n_252),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_234),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_277),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_236),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_299),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_257),
.C(n_279),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_291),
.C(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_291),
.B(n_251),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_271),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_259),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_308),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_232),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_273),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_290),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_315),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_288),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_284),
.B(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_316),
.B(n_318),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_298),
.C(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_299),
.C(n_292),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_321),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_314),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_256),
.C(n_206),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_328),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_309),
.A2(n_198),
.B(n_205),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_306),
.B1(n_273),
.B2(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_287),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_SL g330 ( 
.A(n_318),
.B(n_312),
.Y(n_330)
);

OAI21x1_ASAP7_75t_SL g345 ( 
.A1(n_330),
.A2(n_335),
.B(n_5),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_337),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_305),
.B(n_310),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_310),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_320),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_303),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_5),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_345),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_334),
.A2(n_319),
.B(n_325),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_340),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_330),
.A2(n_315),
.B(n_256),
.C(n_325),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_343),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_331),
.A2(n_229),
.B(n_13),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_329),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_348),
.Y(n_351)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_346),
.A2(n_341),
.B(n_332),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g352 ( 
.A(n_350),
.B(n_349),
.C(n_347),
.Y(n_352)
);

OAI32xp33_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_349),
.A3(n_342),
.B1(n_351),
.B2(n_337),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_336),
.B(n_8),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_8),
.Y(n_356)
);


endmodule