module fake_jpeg_16266_n_52 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_52);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_23),
.B1(n_19),
.B2(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_21),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_41),
.C(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_40),
.B1(n_5),
.B2(n_4),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.C(n_45),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_9),
.C(n_10),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_15),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_49),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_47),
.B1(n_46),
.B2(n_18),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_16),
.B(n_17),
.Y(n_52)
);


endmodule