module real_jpeg_14221_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_0),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_24),
.C(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_0),
.B(n_88),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_0),
.A2(n_8),
.B(n_23),
.C(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_0),
.B(n_37),
.C(n_40),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_0),
.B(n_18),
.Y(n_137)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_26),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_10),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_107),
.CON(n_11),
.SN(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_105),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_93),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_14),
.B(n_93),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_14),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_60),
.CI(n_77),
.CON(n_14),
.SN(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_32),
.C(n_46),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_16),
.A2(n_32),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_16),
.A2(n_71),
.B1(n_76),
.B2(n_98),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B(n_27),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_17),
.A2(n_22),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

O2A1O1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_20),
.B(n_24),
.C(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_21),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_19),
.A2(n_20),
.B(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_21),
.B(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_29),
.B(n_64),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_29),
.B(n_43),
.Y(n_149)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_43),
.B(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_45),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_34),
.A2(n_38),
.B1(n_45),
.B2(n_73),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_39),
.B(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_72),
.B(n_74),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_47),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_56),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_81),
.Y(n_80)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_58),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_64),
.B(n_66),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_68),
.B1(n_70),
.B2(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_66),
.B(n_83),
.Y(n_102)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_98),
.C(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_71),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_71),
.A2(n_76),
.B1(n_133),
.B2(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_82),
.A2(n_100),
.B1(n_136),
.B2(n_139),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_82),
.B(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_126),
.C(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_90),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_102),
.C(n_103),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_101),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_101),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_160),
.B(n_164),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_129),
.B(n_159),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_117),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_117),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_111),
.A2(n_112),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_126),
.C(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_128),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_153),
.B(n_158),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_140),
.B(n_152),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B(n_151),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_148),
.B(n_150),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);


endmodule