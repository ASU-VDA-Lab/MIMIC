module fake_aes_11429_n_652 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_652);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_652;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_68), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_43), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_44), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_13), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_35), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_61), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_47), .Y(n_82) );
CKINVDCx14_ASAP7_75t_R g83 ( .A(n_46), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_13), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_4), .Y(n_85) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_67), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_11), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_50), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_56), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_6), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_54), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
BUFx10_ASAP7_75t_L g97 ( .A(n_40), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_18), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_21), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_29), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_58), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_37), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_63), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_33), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_3), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_28), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_21), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_41), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_19), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_22), .Y(n_115) );
BUFx10_ASAP7_75t_L g116 ( .A(n_23), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_45), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_70), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_42), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_65), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_76), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_75), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_109), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_117), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_113), .B(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_78), .B(n_0), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_117), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_120), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_78), .B(n_1), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_80), .B(n_1), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_86), .B(n_2), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_84), .B(n_2), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_97), .B(n_3), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_94), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_87), .B(n_4), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_85), .B(n_5), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_87), .B(n_5), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_103), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_103), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_105), .Y(n_159) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_105), .B(n_32), .Y(n_160) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_160), .B(n_119), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_131), .A2(n_114), .B1(n_99), .B2(n_92), .Y(n_162) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_160), .Y(n_163) );
INVxp67_ASAP7_75t_SL g164 ( .A(n_151), .Y(n_164) );
INVxp67_ASAP7_75t_SL g165 ( .A(n_151), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_141), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_131), .B(n_92), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_135), .B(n_111), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
AND2x6_ASAP7_75t_L g175 ( .A(n_135), .B(n_119), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_126), .B(n_116), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_126), .B(n_116), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_125), .B(n_104), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_122), .B(n_91), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_123), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_123), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_123), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_149), .B(n_102), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_123), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_122), .B(n_91), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_132), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_132), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_124), .B(n_100), .Y(n_199) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_144), .A2(n_107), .B1(n_99), .B2(n_114), .C(n_111), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_124), .B(n_83), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_127), .B(n_116), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_160), .A2(n_107), .B1(n_115), .B2(n_108), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_153), .A2(n_112), .B1(n_110), .B2(n_118), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_127), .B(n_106), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_153), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_130), .B(n_118), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_121), .Y(n_209) );
AO22x2_ASAP7_75t_L g210 ( .A1(n_136), .A2(n_112), .B1(n_110), .B2(n_82), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_130), .B(n_90), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_121), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_129), .B(n_116), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_121), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_137), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_211), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_213), .B(n_159), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_175), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_213), .B(n_159), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_211), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_175), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_169), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_212), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_164), .B(n_136), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_213), .B(n_150), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_212), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_165), .B(n_155), .Y(n_230) );
INVxp67_ASAP7_75t_SL g231 ( .A(n_169), .Y(n_231) );
BUFx2_ASAP7_75t_SL g232 ( .A(n_175), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_195), .B(n_155), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_213), .B(n_152), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_175), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_166), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_178), .B(n_143), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_215), .B(n_152), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_187), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_166), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_215), .B(n_157), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_163), .A2(n_140), .B1(n_157), .B2(n_145), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_163), .A2(n_142), .B1(n_145), .B2(n_147), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_163), .A2(n_142), .B1(n_147), .B2(n_140), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_193), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_161), .A2(n_150), .B1(n_143), .B2(n_154), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_210), .A2(n_156), .B1(n_154), .B2(n_144), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_161), .A2(n_156), .B1(n_146), .B2(n_148), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
INVx4_ASAP7_75t_L g254 ( .A(n_175), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_195), .B(n_158), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_201), .B(n_158), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_193), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_161), .A2(n_158), .B1(n_148), .B2(n_139), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_175), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_166), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_174), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_193), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_174), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_190), .Y(n_265) );
OR2x2_ASAP7_75t_SL g266 ( .A(n_203), .B(n_98), .Y(n_266) );
INVx5_ASAP7_75t_L g267 ( .A(n_175), .Y(n_267) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_174), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_179), .B(n_148), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_189), .B(n_139), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_202), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_168), .B(n_139), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_169), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_168), .B(n_138), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_180), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_190), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g277 ( .A1(n_210), .A2(n_97), .B1(n_138), .B2(n_101), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_254), .B(n_220), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_254), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_240), .B(n_162), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
AND2x6_ASAP7_75t_L g284 ( .A(n_220), .B(n_176), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_SL g286 ( .A1(n_256), .A2(n_206), .B(n_205), .C(n_170), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_244), .B(n_210), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_222), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_246), .A2(n_176), .B1(n_166), .B2(n_168), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_223), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_263), .A2(n_176), .B1(n_168), .B2(n_171), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_218), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_272), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_225), .B(n_184), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_268), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_248), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_223), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_241), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_259), .Y(n_302) );
BUFx4f_ASAP7_75t_L g303 ( .A(n_272), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_248), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_259), .B(n_171), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_271), .B(n_200), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_226), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_259), .Y(n_308) );
AND2x4_ASAP7_75t_SL g309 ( .A(n_233), .B(n_184), .Y(n_309) );
INVx5_ASAP7_75t_L g310 ( .A(n_236), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_251), .A2(n_171), .B1(n_192), .B2(n_184), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_236), .B(n_171), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_275), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_246), .A2(n_199), .B(n_207), .C(n_184), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_226), .Y(n_316) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_233), .A2(n_192), .B1(n_207), .B2(n_97), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_236), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_229), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_261), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_255), .B(n_192), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_255), .B(n_192), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_236), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_314), .A2(n_250), .B1(n_270), .B2(n_258), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_283), .Y(n_326) );
BUFx4_ASAP7_75t_R g327 ( .A(n_284), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_306), .A2(n_230), .B1(n_227), .B2(n_238), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_315), .A2(n_269), .B(n_258), .C(n_252), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_230), .B1(n_227), .B2(n_277), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_296), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_309), .B(n_250), .Y(n_333) );
CKINVDCx8_ASAP7_75t_R g334 ( .A(n_314), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_284), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_317), .A2(n_252), .B1(n_245), .B2(n_247), .C(n_270), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_309), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_296), .B(n_266), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_281), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_281), .A2(n_264), .B(n_239), .Y(n_340) );
CKINVDCx11_ASAP7_75t_R g341 ( .A(n_313), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_303), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_303), .B(n_272), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_312), .A2(n_274), .B1(n_232), .B2(n_266), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_279), .B(n_236), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_293), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_279), .B(n_236), .Y(n_349) );
INVx4_ASAP7_75t_L g350 ( .A(n_284), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_303), .A2(n_232), .B1(n_207), .B2(n_274), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
AO22x2_ASAP7_75t_L g353 ( .A1(n_287), .A2(n_274), .B1(n_229), .B2(n_239), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_305), .A2(n_274), .B1(n_273), .B2(n_268), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_338), .B(n_322), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_342), .Y(n_356) );
INVx6_ASAP7_75t_L g357 ( .A(n_347), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_346), .A2(n_282), .B1(n_290), .B2(n_294), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_342), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_337), .B(n_305), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_344), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_337), .A2(n_294), .B1(n_293), .B2(n_319), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_335), .Y(n_364) );
AOI221x1_ASAP7_75t_SL g365 ( .A1(n_325), .A2(n_138), .B1(n_207), .B2(n_134), .C(n_128), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_331), .A2(n_323), .B1(n_295), .B2(n_311), .C1(n_228), .C2(n_219), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_328), .A2(n_292), .B1(n_234), .B2(n_221), .C(n_204), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_338), .A2(n_307), .B1(n_319), .B2(n_316), .Y(n_368) );
BUFx5_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_333), .A2(n_307), .B1(n_316), .B2(n_273), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_336), .A2(n_286), .B1(n_235), .B2(n_264), .C(n_134), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_339), .B(n_235), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_134), .B1(n_133), .B2(n_128), .C(n_304), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_330), .A2(n_273), .B1(n_284), .B2(n_268), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_348), .Y(n_375) );
OAI31xp33_ASAP7_75t_L g376 ( .A1(n_329), .A2(n_297), .A3(n_285), .B(n_313), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_326), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_340), .A2(n_268), .B(n_297), .C(n_320), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_332), .Y(n_380) );
AOI31xp33_ASAP7_75t_L g381 ( .A1(n_363), .A2(n_327), .A3(n_351), .B(n_332), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_360), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_360), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_364), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_368), .A2(n_353), .B1(n_343), .B2(n_335), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_362), .B(n_352), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_366), .A2(n_353), .B1(n_345), .B2(n_341), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_359), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_362), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_356), .B(n_345), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_376), .A2(n_334), .B(n_341), .C(n_354), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_378), .A2(n_380), .B(n_377), .Y(n_392) );
OAI31xp33_ASAP7_75t_L g393 ( .A1(n_367), .A2(n_285), .A3(n_349), .B(n_347), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_379), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_355), .A2(n_369), .B1(n_358), .B2(n_374), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_375), .A2(n_334), .B(n_128), .C(n_133), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_365), .A2(n_133), .B1(n_298), .B2(n_321), .C(n_320), .Y(n_398) );
OAI222xp33_ASAP7_75t_SL g399 ( .A1(n_369), .A2(n_350), .B1(n_335), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_399) );
OAI31xp33_ASAP7_75t_L g400 ( .A1(n_355), .A2(n_349), .A3(n_347), .B(n_313), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_357), .A2(n_350), .B1(n_343), .B2(n_299), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_370), .A2(n_350), .B1(n_298), .B2(n_304), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_373), .B(n_193), .C(n_173), .Y(n_403) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_379), .B(n_209), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_372), .B(n_321), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_371), .B(n_193), .C(n_173), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_369), .A2(n_349), .B1(n_284), .B2(n_97), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_372), .B(n_209), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_369), .A2(n_284), .B1(n_231), .B2(n_216), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_361), .B(n_214), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g412 ( .A1(n_364), .A2(n_214), .B(n_216), .C(n_279), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_361), .B(n_302), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_357), .A2(n_299), .B1(n_224), .B2(n_308), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_382), .B(n_369), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_382), .B(n_369), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_383), .B(n_369), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_383), .B(n_369), .Y(n_418) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_385), .A2(n_389), .A3(n_396), .B1(n_386), .B2(n_401), .B3(n_410), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_388), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_394), .B(n_357), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_405), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_391), .B(n_197), .C(n_185), .Y(n_425) );
OAI33xp33_ASAP7_75t_L g426 ( .A1(n_386), .A2(n_185), .A3(n_198), .B1(n_197), .B2(n_191), .B3(n_188), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
AOI33xp33_ASAP7_75t_L g428 ( .A1(n_387), .A2(n_395), .A3(n_390), .B1(n_408), .B2(n_405), .B3(n_407), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_411), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_384), .B(n_411), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_384), .B(n_364), .Y(n_431) );
OAI221xp5_ASAP7_75t_SL g432 ( .A1(n_393), .A2(n_186), .B1(n_198), .B2(n_188), .C(n_191), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_412), .B(n_193), .C(n_173), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_408), .Y(n_434) );
NAND4xp25_ASAP7_75t_L g435 ( .A(n_393), .B(n_186), .C(n_172), .D(n_183), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_390), .A2(n_357), .B1(n_364), .B2(n_299), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_381), .B(n_6), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_381), .A2(n_364), .B(n_280), .Y(n_438) );
OAI33xp33_ASAP7_75t_L g439 ( .A1(n_402), .A2(n_170), .A3(n_183), .B1(n_182), .B2(n_177), .B3(n_172), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_404), .B(n_7), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_384), .B(n_7), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
OAI31xp33_ASAP7_75t_L g445 ( .A1(n_399), .A2(n_224), .A3(n_280), .B(n_206), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_398), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_413), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_392), .B(n_9), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_400), .A2(n_167), .B1(n_177), .B2(n_182), .C(n_173), .Y(n_449) );
OAI221xp5_ASAP7_75t_SL g450 ( .A1(n_400), .A2(n_167), .B1(n_194), .B2(n_196), .C(n_16), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_409), .B(n_12), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_414), .A2(n_12), .A3(n_14), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_403), .B(n_310), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_403), .B(n_409), .Y(n_454) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_406), .B(n_308), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_406), .B(n_14), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_405), .B(n_15), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_382), .B(n_17), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_388), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_391), .B(n_194), .C(n_196), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_382), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_412), .B(n_173), .C(n_208), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_423), .B(n_19), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_420), .B(n_20), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_421), .B(n_20), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_421), .B(n_25), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_420), .B(n_26), .Y(n_467) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_437), .A2(n_308), .B1(n_280), .B2(n_278), .C(n_300), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_461), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_461), .B(n_27), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
OAI211xp5_ASAP7_75t_L g472 ( .A1(n_438), .A2(n_310), .B(n_267), .C(n_300), .Y(n_472) );
AND2x4_ASAP7_75t_SL g473 ( .A(n_434), .B(n_289), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_459), .B(n_30), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_446), .A2(n_300), .B1(n_291), .B2(n_289), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_424), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_447), .B(n_31), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_424), .B(n_36), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_429), .B(n_38), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_443), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_427), .Y(n_482) );
OAI33xp33_ASAP7_75t_L g483 ( .A1(n_457), .A2(n_39), .A3(n_49), .B1(n_51), .B2(n_52), .B3(n_53), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_443), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_415), .B(n_55), .Y(n_486) );
AOI31xp33_ASAP7_75t_L g487 ( .A1(n_419), .A2(n_57), .A3(n_60), .B(n_64), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
AOI221x1_ASAP7_75t_L g489 ( .A1(n_433), .A2(n_66), .B1(n_69), .B2(n_71), .C(n_72), .Y(n_489) );
AOI21xp33_ASAP7_75t_SL g490 ( .A1(n_438), .A2(n_73), .B(n_237), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_415), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_458), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_458), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_422), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_416), .B(n_208), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_422), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_452), .B(n_208), .C(n_237), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_428), .B(n_208), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_441), .B(n_278), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_416), .B(n_278), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_451), .A2(n_291), .B(n_289), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_417), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_417), .B(n_300), .Y(n_503) );
NOR2x1_ASAP7_75t_L g504 ( .A(n_433), .B(n_300), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_418), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_418), .B(n_278), .Y(n_506) );
NAND4xp25_ASAP7_75t_L g507 ( .A(n_450), .B(n_237), .C(n_260), .D(n_243), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_441), .B(n_291), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_462), .B(n_291), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_430), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_430), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_448), .B(n_237), .C(n_260), .D(n_243), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_430), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_456), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_448), .B(n_278), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_440), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_440), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_492), .B(n_442), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_464), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_471), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_469), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_477), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_471), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_477), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_496), .B(n_444), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_475), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_482), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_493), .B(n_456), .Y(n_529) );
INVxp67_ASAP7_75t_SL g530 ( .A(n_481), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_514), .B(n_444), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_482), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_491), .B(n_454), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_491), .B(n_454), .Y(n_534) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_487), .A2(n_435), .B(n_455), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_502), .B(n_455), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_502), .B(n_455), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_512), .A2(n_446), .B1(n_435), .B2(n_436), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_513), .B(n_431), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_464), .B(n_446), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_505), .B(n_431), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_475), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_505), .B(n_436), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_494), .B(n_465), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_516), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_465), .B(n_431), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_484), .B(n_462), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_463), .B(n_453), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_517), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_463), .B(n_445), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_473), .B(n_445), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_473), .B(n_449), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_513), .B(n_460), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_474), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_498), .B(n_432), .C(n_426), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_474), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_507), .A2(n_439), .B1(n_425), .B2(n_289), .Y(n_560) );
AOI211x1_ASAP7_75t_L g561 ( .A1(n_468), .A2(n_478), .B(n_472), .C(n_486), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_488), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_467), .A2(n_310), .B1(n_267), .B2(n_318), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_513), .B(n_257), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_467), .B(n_262), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_561), .B(n_490), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_520), .B(n_483), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_534), .B(n_510), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_535), .B(n_504), .Y(n_569) );
XNOR2x1_ASAP7_75t_L g570 ( .A(n_553), .B(n_486), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_552), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g572 ( .A1(n_558), .A2(n_479), .B(n_470), .C(n_466), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_534), .B(n_511), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_533), .B(n_511), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_530), .B(n_510), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_519), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_522), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_547), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_540), .B(n_506), .Y(n_579) );
NOR2xp33_ASAP7_75t_SL g580 ( .A(n_541), .B(n_479), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_563), .A2(n_509), .B(n_489), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_518), .B(n_495), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_523), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_540), .B(n_506), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_525), .Y(n_586) );
XNOR2xp5_ASAP7_75t_L g587 ( .A(n_546), .B(n_495), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_562), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_540), .B(n_503), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_557), .B(n_515), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_559), .B(n_466), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_543), .B(n_500), .Y(n_592) );
XNOR2xp5_ASAP7_75t_L g593 ( .A(n_548), .B(n_503), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_529), .B(n_470), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_551), .B(n_508), .Y(n_595) );
AOI32xp33_ASAP7_75t_L g596 ( .A1(n_541), .A2(n_480), .A3(n_497), .B1(n_476), .B2(n_499), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g597 ( .A1(n_536), .A2(n_480), .B1(n_489), .B2(n_501), .C1(n_500), .C2(n_243), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_528), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_539), .A2(n_560), .B1(n_554), .B2(n_545), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_532), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_562), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_538), .B(n_243), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_542), .B(n_260), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_560), .A2(n_310), .B(n_260), .C(n_318), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_549), .B(n_257), .C(n_265), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_531), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_555), .A2(n_324), .B(n_318), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_543), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_556), .A2(n_267), .B1(n_310), .B2(n_318), .C(n_324), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_536), .A2(n_267), .B1(n_318), .B2(n_324), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g611 ( .A1(n_537), .A2(n_257), .B1(n_276), .B2(n_253), .C(n_242), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_537), .A2(n_242), .B1(n_276), .B2(n_253), .C(n_265), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_556), .A2(n_267), .B1(n_324), .B2(n_249), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_526), .B(n_249), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_521), .B(n_249), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_524), .Y(n_616) );
OAI211xp5_ASAP7_75t_L g617 ( .A1(n_565), .A2(n_249), .B(n_262), .C(n_524), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_527), .B(n_249), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_527), .B(n_262), .Y(n_619) );
OA22x2_ASAP7_75t_L g620 ( .A1(n_544), .A2(n_262), .B1(n_564), .B2(n_565), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_566), .A2(n_596), .B(n_567), .C(n_572), .Y(n_621) );
NOR5xp2_ASAP7_75t_L g622 ( .A(n_601), .B(n_588), .C(n_572), .D(n_611), .E(n_617), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_567), .B(n_606), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_569), .A2(n_620), .B(n_570), .Y(n_624) );
NAND3x1_ASAP7_75t_L g625 ( .A(n_582), .B(n_605), .C(n_591), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_599), .B(n_597), .C(n_604), .D(n_580), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_582), .B(n_609), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_620), .A2(n_588), .B1(n_592), .B2(n_583), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_595), .A2(n_590), .B1(n_608), .B2(n_591), .Y(n_629) );
OAI21xp33_ASAP7_75t_SL g630 ( .A1(n_614), .A2(n_585), .B(n_589), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_579), .A2(n_607), .B1(n_594), .B2(n_587), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_571), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_575), .Y(n_633) );
OA22x2_ASAP7_75t_L g634 ( .A1(n_621), .A2(n_593), .B1(n_579), .B2(n_573), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_628), .A2(n_609), .B(n_610), .C(n_613), .Y(n_635) );
OAI31xp33_ASAP7_75t_L g636 ( .A1(n_624), .A2(n_584), .A3(n_600), .B(n_598), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_630), .A2(n_581), .B(n_578), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_627), .A2(n_602), .B(n_603), .C(n_574), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_631), .B(n_616), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_632), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g641 ( .A(n_636), .B(n_622), .C(n_625), .Y(n_641) );
AOI32xp33_ASAP7_75t_L g642 ( .A1(n_635), .A2(n_623), .A3(n_633), .B1(n_626), .B2(n_568), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_634), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_SL g644 ( .A1(n_637), .A2(n_632), .B(n_586), .C(n_576), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_643), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_641), .B(n_629), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_645), .Y(n_647) );
XNOR2xp5_ASAP7_75t_L g648 ( .A(n_646), .B(n_642), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_644), .B1(n_577), .B2(n_564), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_649), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_647), .B(n_648), .C(n_612), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_618), .A3(n_619), .B(n_615), .Y(n_652) );
endmodule