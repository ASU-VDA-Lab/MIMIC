module fake_ibex_1231_n_3468 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_667, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_673, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_679, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_672, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_675, n_463, n_624, n_411, n_135, n_520, n_658, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3468);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_673;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_679;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_672;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_658;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3468;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_3255;
wire n_3272;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_1668;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2806;
wire n_2283;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_3427;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_3162;
wire n_2732;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_3085;
wire n_3059;
wire n_2567;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_3163;
wire n_2929;
wire n_3343;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_3067;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_2928;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_3124;
wire n_999;
wire n_2634;
wire n_3286;
wire n_2982;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_3081;
wire n_2492;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2618;
wire n_2303;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_3247;
wire n_1891;
wire n_1026;
wire n_2681;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_866;

BUFx2_ASAP7_75t_L g680 ( 
.A(n_195),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_173),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_290),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_536),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_234),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_537),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_266),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_544),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_539),
.B(n_266),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_31),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_138),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_104),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_653),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_658),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_326),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_369),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_27),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_678),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_0),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_513),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_358),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_608),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_519),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_668),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_501),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_597),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_677),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_500),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_477),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_4),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_667),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_85),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_280),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_384),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_376),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_292),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_650),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_225),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_71),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_212),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_483),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_659),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_423),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_169),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_544),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_130),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_184),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_204),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_343),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_230),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_243),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_22),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_633),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_253),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_647),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_216),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_324),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_92),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_481),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_598),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_69),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_232),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_421),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_90),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_453),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_386),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_661),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_231),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_529),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_83),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_203),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_90),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_406),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_298),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_144),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_583),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_557),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_359),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_135),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_593),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_498),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_663),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_258),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_630),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_306),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_20),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_25),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_660),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_81),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_174),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_254),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_285),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_463),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_594),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_8),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_576),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_85),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_649),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_170),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_313),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_578),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_591),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_398),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_340),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_523),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_365),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_196),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_291),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_622),
.Y(n_790)
);

BUFx5_ASAP7_75t_L g791 ( 
.A(n_264),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_441),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_73),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_51),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_560),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_230),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_262),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_107),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_264),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_600),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_542),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_309),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_26),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_442),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_644),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_193),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_289),
.Y(n_807)
);

BUFx8_ASAP7_75t_SL g808 ( 
.A(n_228),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_379),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_552),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_176),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_584),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_35),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_52),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_173),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_675),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_627),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_61),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_545),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_210),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_318),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_643),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_318),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_303),
.B(n_430),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_188),
.Y(n_825)
);

CKINVDCx16_ASAP7_75t_R g826 ( 
.A(n_43),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_140),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_582),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_121),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_289),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_601),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_327),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_258),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_132),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_590),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_129),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_528),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_39),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_122),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_532),
.Y(n_840)
);

BUFx10_ASAP7_75t_L g841 ( 
.A(n_439),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_118),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_22),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_592),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_539),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_99),
.Y(n_846)
);

CKINVDCx16_ASAP7_75t_R g847 ( 
.A(n_512),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_381),
.Y(n_848)
);

BUFx5_ASAP7_75t_L g849 ( 
.A(n_234),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_376),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_311),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_32),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_220),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_276),
.Y(n_854)
);

CKINVDCx16_ASAP7_75t_R g855 ( 
.A(n_103),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_300),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_548),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_260),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_327),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_586),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_50),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_400),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_380),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_589),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_365),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_379),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_347),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_543),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_180),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_464),
.Y(n_870)
);

BUFx10_ASAP7_75t_L g871 ( 
.A(n_95),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_487),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_88),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_133),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_241),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_398),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_384),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_372),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_112),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_634),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_29),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_554),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_298),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_458),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_561),
.Y(n_885)
);

BUFx8_ASAP7_75t_SL g886 ( 
.A(n_101),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_330),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_387),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_344),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_177),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_65),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_374),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_104),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_607),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_123),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_216),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_259),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_311),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_107),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_30),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_301),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_60),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_80),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_423),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_317),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_615),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_247),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_356),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_390),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_399),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_300),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_147),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_673),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_224),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_520),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_364),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_199),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_11),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_175),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_13),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_414),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_293),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_75),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_180),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_461),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_418),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_161),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_474),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_632),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_519),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_207),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_626),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_638),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_651),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_196),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_538),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_275),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_478),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_657),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_282),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_324),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_357),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_172),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_581),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_155),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_165),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_151),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_273),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_171),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_535),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_329),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_197),
.Y(n_952)
);

BUFx10_ASAP7_75t_L g953 ( 
.A(n_25),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_59),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_609),
.Y(n_955)
);

CKINVDCx16_ASAP7_75t_R g956 ( 
.A(n_269),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_504),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_641),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_121),
.Y(n_959)
);

BUFx8_ASAP7_75t_SL g960 ( 
.A(n_78),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_656),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_611),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_540),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_43),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_290),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_382),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_115),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_67),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_75),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_553),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_363),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_112),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_125),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_69),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_116),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_577),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_197),
.Y(n_977)
);

CKINVDCx16_ASAP7_75t_R g978 ( 
.A(n_666),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_532),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_116),
.Y(n_980)
);

BUFx2_ASAP7_75t_SL g981 ( 
.A(n_165),
.Y(n_981)
);

CKINVDCx14_ASAP7_75t_R g982 ( 
.A(n_564),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_31),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_203),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_364),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_416),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_192),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_351),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_23),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_361),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_21),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_646),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_81),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_308),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_7),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_652),
.Y(n_996)
);

BUFx2_ASAP7_75t_SL g997 ( 
.A(n_552),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_L g998 ( 
.A(n_326),
.B(n_531),
.Y(n_998)
);

BUFx8_ASAP7_75t_SL g999 ( 
.A(n_345),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_454),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_255),
.Y(n_1001)
);

CKINVDCx16_ASAP7_75t_R g1002 ( 
.A(n_63),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_480),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_339),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_238),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_629),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_541),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_48),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_88),
.Y(n_1009)
);

BUFx5_ASAP7_75t_L g1010 ( 
.A(n_500),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_482),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_378),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_132),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_87),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_547),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_239),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_227),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_338),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_521),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_19),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_241),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_310),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_635),
.Y(n_1023)
);

BUFx10_ASAP7_75t_L g1024 ( 
.A(n_596),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_429),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_543),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_479),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_636),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_606),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_194),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_42),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_239),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_163),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_511),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_346),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_263),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_469),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_350),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_147),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_458),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_170),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_73),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_54),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_466),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_99),
.Y(n_1045)
);

BUFx10_ASAP7_75t_L g1046 ( 
.A(n_616),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_SL g1047 ( 
.A1(n_699),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_683),
.B(n_1),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_737),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_683),
.B(n_2),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_791),
.Y(n_1051)
);

BUFx8_ASAP7_75t_L g1052 ( 
.A(n_692),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_791),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_737),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_737),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_810),
.B(n_3),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_709),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_791),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_680),
.B(n_3),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_747),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_737),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_791),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_785),
.B(n_5),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_978),
.Y(n_1064)
);

CKINVDCx6p67_ASAP7_75t_R g1065 ( 
.A(n_709),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_814),
.Y(n_1066)
);

AOI22x1_ASAP7_75t_SL g1067 ( 
.A1(n_719),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_752),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_752),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_705),
.B(n_9),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_709),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_791),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_707),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_791),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_808),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_791),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_761),
.Y(n_1077)
);

BUFx8_ASAP7_75t_SL g1078 ( 
.A(n_808),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_707),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_701),
.A2(n_556),
.B(n_555),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_701),
.A2(n_976),
.B(n_706),
.Y(n_1081)
);

OAI22x1_ASAP7_75t_R g1082 ( 
.A1(n_719),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_849),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_752),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_961),
.B(n_10),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_752),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_707),
.Y(n_1087)
);

AOI22x1_ASAP7_75t_SL g1088 ( 
.A1(n_723),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_849),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_SL g1090 ( 
.A1(n_723),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_849),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_886),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_706),
.A2(n_559),
.B(n_558),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_766),
.Y(n_1094)
);

OA21x2_ASAP7_75t_L g1095 ( 
.A1(n_976),
.A2(n_563),
.B(n_562),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_766),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_766),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_849),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_682),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_682),
.B(n_718),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_714),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_718),
.B(n_16),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_766),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_827),
.Y(n_1104)
);

AOI22x1_ASAP7_75t_SL g1105 ( 
.A1(n_727),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1105)
);

AND2x6_ASAP7_75t_L g1106 ( 
.A(n_748),
.B(n_565),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_787),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_693),
.A2(n_567),
.B(n_566),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_703),
.A2(n_569),
.B(n_568),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_848),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_848),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_884),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_827),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_827),
.Y(n_1114)
);

BUFx8_ASAP7_75t_SL g1115 ( 
.A(n_886),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_983),
.B(n_17),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_983),
.B(n_18),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_711),
.A2(n_571),
.B(n_570),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_846),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_846),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_1024),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_834),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1034),
.B(n_19),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1034),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_850),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_846),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_991),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1010),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_684),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_684),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_796),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_991),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_796),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1010),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_991),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_874),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_991),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_932),
.B(n_20),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_990),
.Y(n_1139)
);

CKINVDCx6p67_ASAP7_75t_R g1140 ( 
.A(n_1024),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1020),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1078),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1078),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1056),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_1060),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1056),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1115),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1115),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1075),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1101),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1092),
.Y(n_1151)
);

CKINVDCx16_ASAP7_75t_R g1152 ( 
.A(n_1057),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1064),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_1065),
.B(n_982),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1140),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1052),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1052),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1117),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1066),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1112),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_1108),
.A2(n_734),
.B(n_725),
.Y(n_1161)
);

NAND2xp33_ASAP7_75t_R g1162 ( 
.A(n_1048),
.B(n_712),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1101),
.B(n_1005),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1122),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1049),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1123),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1057),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1122),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1125),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_R g1170 ( 
.A(n_1050),
.B(n_712),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1125),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1099),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1139),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1139),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1071),
.B(n_713),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1082),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1059),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_1100),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1071),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_1073),
.B(n_982),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1121),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1110),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_R g1183 ( 
.A(n_1073),
.B(n_697),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1121),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1079),
.B(n_874),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1111),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1124),
.Y(n_1187)
);

INVx6_ASAP7_75t_L g1188 ( 
.A(n_1049),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1070),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1070),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1087),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_R g1192 ( 
.A(n_1107),
.B(n_697),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_1063),
.B(n_1008),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1067),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1102),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1088),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1105),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_1047),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1102),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_1077),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1085),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1053),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1085),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1090),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1062),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_1129),
.B(n_939),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1138),
.Y(n_1207)
);

CKINVDCx16_ASAP7_75t_R g1208 ( 
.A(n_1106),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1116),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1138),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1130),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1131),
.B(n_951),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1133),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1136),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1106),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1106),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1106),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1080),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1081),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1072),
.B(n_932),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1074),
.Y(n_1221)
);

NAND2xp33_ASAP7_75t_R g1222 ( 
.A(n_1109),
.B(n_713),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1083),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1080),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1098),
.B(n_702),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1128),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1051),
.Y(n_1227)
);

OR2x6_ASAP7_75t_L g1228 ( 
.A(n_1118),
.B(n_981),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1134),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1080),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1058),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1076),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1089),
.B(n_744),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1091),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1049),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1093),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1049),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1054),
.B(n_1024),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_R g1239 ( 
.A(n_1109),
.B(n_715),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1141),
.B(n_715),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_R g1241 ( 
.A(n_1054),
.B(n_958),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1054),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1054),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_1055),
.B(n_958),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1055),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1055),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1141),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1093),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1141),
.Y(n_1249)
);

AND2x6_ASAP7_75t_L g1250 ( 
.A(n_1061),
.B(n_748),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1061),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1068),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1068),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1068),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1069),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1141),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1069),
.B(n_936),
.Y(n_1257)
);

INVxp33_ASAP7_75t_SL g1258 ( 
.A(n_1093),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1137),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1095),
.B(n_781),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1095),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1095),
.B(n_798),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1069),
.B(n_948),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1069),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1084),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1109),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1084),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1084),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1084),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1086),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1086),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_R g1272 ( 
.A(n_1086),
.B(n_717),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1137),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1137),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1086),
.B(n_951),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1094),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1094),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1094),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1096),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1096),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1096),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1097),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_R g1283 ( 
.A(n_1097),
.B(n_722),
.Y(n_1283)
);

NOR2x1p5_ASAP7_75t_L g1284 ( 
.A(n_1097),
.B(n_716),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1103),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1103),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1103),
.Y(n_1287)
);

INVx4_ASAP7_75t_L g1288 ( 
.A(n_1103),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1104),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1135),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1104),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1104),
.Y(n_1292)
);

INVxp67_ASAP7_75t_R g1293 ( 
.A(n_1113),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1113),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_R g1295 ( 
.A(n_1114),
.B(n_722),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1114),
.B(n_1038),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1195),
.Y(n_1297)
);

NAND2xp33_ASAP7_75t_L g1298 ( 
.A(n_1215),
.B(n_758),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1189),
.A2(n_720),
.B1(n_721),
.B2(n_716),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1189),
.B(n_765),
.Y(n_1300)
);

AND2x2_ASAP7_75t_SL g1301 ( 
.A(n_1152),
.B(n_826),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1199),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1190),
.B(n_1046),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1209),
.B(n_1207),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1150),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1153),
.B(n_1150),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1275),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1167),
.B(n_1178),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1174),
.B(n_847),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1200),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1201),
.B(n_782),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1172),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1216),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1203),
.B(n_783),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1193),
.B(n_790),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1182),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1260),
.B(n_1262),
.C(n_1239),
.Y(n_1317)
);

INVx8_ASAP7_75t_L g1318 ( 
.A(n_1155),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1200),
.B(n_805),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1186),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1213),
.B(n_822),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1185),
.B(n_828),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1185),
.B(n_831),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1187),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1158),
.Y(n_1325)
);

NOR3xp33_ASAP7_75t_L g1326 ( 
.A(n_1204),
.B(n_857),
.C(n_855),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1144),
.B(n_844),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_L g1328 ( 
.A(n_1168),
.B(n_901),
.C(n_892),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1278),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1208),
.B(n_860),
.Y(n_1330)
);

NOR3xp33_ASAP7_75t_L g1331 ( 
.A(n_1169),
.B(n_956),
.C(n_910),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1145),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1217),
.Y(n_1333)
);

XOR2xp5_ASAP7_75t_L g1334 ( 
.A(n_1164),
.B(n_727),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1146),
.B(n_864),
.Y(n_1335)
);

NAND3xp33_ASAP7_75t_L g1336 ( 
.A(n_1222),
.B(n_824),
.C(n_688),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1166),
.B(n_885),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1180),
.B(n_894),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1191),
.B(n_913),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1231),
.B(n_929),
.Y(n_1340)
);

AO221x1_ASAP7_75t_L g1341 ( 
.A1(n_1206),
.A2(n_999),
.B1(n_960),
.B2(n_746),
.C(n_786),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1232),
.B(n_934),
.Y(n_1342)
);

NAND2xp33_ASAP7_75t_L g1343 ( 
.A(n_1154),
.B(n_944),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1212),
.Y(n_1344)
);

NOR3xp33_ASAP7_75t_L g1345 ( 
.A(n_1171),
.B(n_1002),
.C(n_694),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1211),
.B(n_955),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1240),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1173),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1214),
.B(n_1221),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1145),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1220),
.A2(n_987),
.B(n_980),
.C(n_690),
.Y(n_1351)
);

AO221x1_ASAP7_75t_L g1352 ( 
.A1(n_1183),
.A2(n_999),
.B1(n_960),
.B2(n_746),
.C(n_786),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1284),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1257),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1219),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1159),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1263),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1296),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1184),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1225),
.B(n_1175),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1163),
.B(n_970),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1226),
.B(n_992),
.Y(n_1362)
);

NOR3xp33_ASAP7_75t_L g1363 ( 
.A(n_1160),
.B(n_738),
.C(n_681),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1227),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_1218),
.B(n_741),
.C(n_736),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1233),
.B(n_1006),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1223),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1179),
.B(n_1023),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1181),
.B(n_1029),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1241),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1228),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1162),
.A2(n_721),
.B1(n_1025),
.B2(n_720),
.Y(n_1372)
);

NAND2xp33_ASAP7_75t_L g1373 ( 
.A(n_1224),
.B(n_1230),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1238),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1177),
.B(n_757),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1228),
.B(n_998),
.Y(n_1376)
);

INVxp33_ASAP7_75t_L g1377 ( 
.A(n_1192),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_1025),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1289),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1228),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1288),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1202),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1244),
.B(n_763),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1205),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1229),
.B(n_685),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1258),
.B(n_1272),
.Y(n_1386)
);

NAND2xp33_ASAP7_75t_L g1387 ( 
.A(n_1236),
.B(n_769),
.Y(n_1387)
);

AO221x1_ASAP7_75t_L g1388 ( 
.A1(n_1156),
.A2(n_815),
.B1(n_875),
.B2(n_733),
.C(n_730),
.Y(n_1388)
);

NOR3xp33_ASAP7_75t_L g1389 ( 
.A(n_1194),
.B(n_829),
.C(n_797),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1161),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1161),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1157),
.B(n_775),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1283),
.B(n_686),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_L g1394 ( 
.A(n_1248),
.B(n_777),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1295),
.B(n_779),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1261),
.B(n_689),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1170),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1250),
.B(n_691),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_SL g1399 ( 
.A(n_1142),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1250),
.B(n_695),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1149),
.B(n_795),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1151),
.B(n_23),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1250),
.B(n_696),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1250),
.B(n_698),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1279),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1281),
.B(n_787),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1266),
.B(n_700),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1282),
.B(n_800),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1288),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1237),
.A2(n_704),
.B(n_708),
.C(n_687),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1198),
.A2(n_1042),
.B1(n_1043),
.B2(n_1041),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1143),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1242),
.B(n_812),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1147),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1243),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1245),
.B(n_710),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1196),
.B(n_817),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1251),
.B(n_724),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1197),
.B(n_787),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1252),
.B(n_835),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1253),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1255),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1264),
.B(n_880),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1267),
.B(n_726),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1269),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1270),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1271),
.B(n_728),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1148),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1277),
.B(n_816),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1280),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1285),
.B(n_882),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1286),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1287),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1291),
.Y(n_1434)
);

AO221x1_ASAP7_75t_L g1435 ( 
.A1(n_1176),
.A2(n_815),
.B1(n_875),
.B2(n_733),
.C(n_730),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1294),
.B(n_729),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1165),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1188),
.B(n_740),
.Y(n_1438)
);

AO221x1_ASAP7_75t_L g1439 ( 
.A1(n_1165),
.A2(n_924),
.B1(n_937),
.B2(n_922),
.C(n_878),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1188),
.B(n_742),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1188),
.B(n_743),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1165),
.Y(n_1442)
);

NOR3xp33_ASAP7_75t_L g1443 ( 
.A(n_1246),
.B(n_1027),
.C(n_1017),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1247),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1249),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1256),
.B(n_745),
.Y(n_1446)
);

NOR3xp33_ASAP7_75t_L g1447 ( 
.A(n_1259),
.B(n_751),
.C(n_749),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1268),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1273),
.B(n_906),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1274),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1276),
.B(n_933),
.Y(n_1451)
);

INVx3_ASAP7_75t_R g1452 ( 
.A(n_1235),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1293),
.Y(n_1453)
);

NAND2x1_ASAP7_75t_L g1454 ( 
.A(n_1290),
.B(n_962),
.Y(n_1454)
);

NOR2xp67_ASAP7_75t_L g1455 ( 
.A(n_1265),
.B(n_24),
.Y(n_1455)
);

AO221x1_ASAP7_75t_L g1456 ( 
.A1(n_1254),
.A2(n_924),
.B1(n_937),
.B2(n_922),
.C(n_878),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1254),
.B(n_996),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1292),
.B(n_754),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1292),
.B(n_1028),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1292),
.B(n_760),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1189),
.B(n_762),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1279),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1174),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1189),
.B(n_764),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1189),
.B(n_767),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1150),
.B(n_792),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1279),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1279),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1275),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1189),
.B(n_771),
.Y(n_1470)
);

NOR3xp33_ASAP7_75t_L g1471 ( 
.A(n_1150),
.B(n_776),
.C(n_774),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1275),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1195),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1195),
.Y(n_1474)
);

NOR2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1157),
.B(n_778),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_SL g1476 ( 
.A(n_1208),
.B(n_816),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1152),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1195),
.B(n_770),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1195),
.B(n_770),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1195),
.B(n_942),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1195),
.B(n_942),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1195),
.B(n_979),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1189),
.B(n_780),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1210),
.B(n_1020),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1195),
.B(n_995),
.Y(n_1485)
);

INVx3_ASAP7_75t_R g1486 ( 
.A(n_1153),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1195),
.B(n_995),
.Y(n_1487)
);

AO221x1_ASAP7_75t_L g1488 ( 
.A1(n_1150),
.A2(n_974),
.B1(n_1000),
.B2(n_965),
.C(n_963),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1189),
.B(n_784),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1150),
.B(n_792),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1189),
.B(n_788),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1195),
.Y(n_1492)
);

NAND2x1_ASAP7_75t_L g1493 ( 
.A(n_1158),
.B(n_1016),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1195),
.Y(n_1494)
);

AO221x1_ASAP7_75t_L g1495 ( 
.A1(n_1150),
.A2(n_1000),
.B1(n_1044),
.B2(n_974),
.C(n_965),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1150),
.B(n_792),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1174),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1215),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1215),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1189),
.B(n_789),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_L g1501 ( 
.A(n_1150),
.B(n_801),
.C(n_799),
.Y(n_1501)
);

NAND2xp33_ASAP7_75t_L g1502 ( 
.A(n_1215),
.B(n_806),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1150),
.B(n_803),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1189),
.B(n_807),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1189),
.B(n_818),
.Y(n_1505)
);

INVxp33_ASAP7_75t_L g1506 ( 
.A(n_1174),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1189),
.B(n_820),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1275),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1195),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1195),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1174),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1297),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1506),
.B(n_1463),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1304),
.A2(n_1044),
.B1(n_732),
.B2(n_735),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1355),
.A2(n_739),
.B(n_731),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1334),
.B(n_997),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1305),
.A2(n_823),
.B1(n_833),
.B2(n_825),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1304),
.B(n_836),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1306),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1497),
.B(n_837),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1511),
.B(n_840),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1371),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1302),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1477),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1371),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1473),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1350),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1474),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1310),
.B(n_839),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

NOR2x2_ASAP7_75t_L g1531 ( 
.A(n_1306),
.B(n_1035),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1462),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1309),
.B(n_858),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1313),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1494),
.B(n_750),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1510),
.B(n_1509),
.Y(n_1536)
);

NOR2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1477),
.B(n_893),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1348),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1325),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1306),
.B(n_803),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1312),
.Y(n_1541)
);

NOR2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1428),
.B(n_904),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1467),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1466),
.B(n_753),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1316),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1317),
.A2(n_756),
.B1(n_759),
.B2(n_755),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1468),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1320),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1318),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1360),
.B(n_1483),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1324),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1336),
.A2(n_772),
.B1(n_773),
.B2(n_768),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1364),
.Y(n_1553)
);

NOR2x2_ASAP7_75t_L g1554 ( 
.A(n_1486),
.B(n_1035),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1489),
.B(n_863),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1344),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1507),
.B(n_865),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1318),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1387),
.A2(n_869),
.B1(n_872),
.B2(n_866),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1476),
.B(n_879),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_R g1561 ( 
.A(n_1318),
.B(n_883),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1461),
.B(n_887),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1406),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1478),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1332),
.B(n_793),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1453),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1390),
.A2(n_802),
.B(n_794),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1356),
.B(n_803),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1301),
.B(n_841),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1464),
.B(n_888),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1405),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1313),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1399),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1490),
.B(n_804),
.Y(n_1574)
);

AO21x1_ASAP7_75t_L g1575 ( 
.A1(n_1391),
.A2(n_811),
.B(n_809),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1300),
.B(n_891),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1414),
.A2(n_899),
.B1(n_902),
.B2(n_898),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1299),
.B(n_1496),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1465),
.B(n_903),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1470),
.B(n_1500),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1367),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1503),
.B(n_905),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1493),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1434),
.B(n_907),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1396),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1412),
.B(n_813),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1475),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1313),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1379),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1479),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1479),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1434),
.B(n_911),
.Y(n_1592)
);

AND2x6_ASAP7_75t_SL g1593 ( 
.A(n_1419),
.B(n_819),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1394),
.A2(n_915),
.B1(n_916),
.B2(n_914),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1376),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1399),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1434),
.Y(n_1597)
);

NOR2xp67_ASAP7_75t_SL g1598 ( 
.A(n_1333),
.B(n_918),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1491),
.B(n_919),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1504),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1480),
.Y(n_1601)
);

NOR3xp33_ASAP7_75t_SL g1602 ( 
.A(n_1375),
.B(n_928),
.C(n_926),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1505),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1407),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1481),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1482),
.B(n_931),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1307),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1372),
.B(n_935),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1471),
.A2(n_940),
.B1(n_941),
.B2(n_938),
.Y(n_1609)
);

BUFx4f_ASAP7_75t_L g1610 ( 
.A(n_1376),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1469),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1485),
.B(n_945),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1333),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1337),
.A2(n_830),
.B(n_821),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1359),
.B(n_832),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1333),
.B(n_1498),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1485),
.B(n_946),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1402),
.B(n_838),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1397),
.B(n_949),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1336),
.A2(n_842),
.B(n_851),
.C(n_845),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1365),
.A2(n_853),
.B1(n_854),
.B2(n_852),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1349),
.B(n_954),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1487),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1487),
.B(n_957),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1472),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1447),
.B(n_856),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1319),
.B(n_1353),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1365),
.A2(n_861),
.B1(n_862),
.B2(n_859),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1347),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1498),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1370),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_SL g1632 ( 
.A(n_1377),
.B(n_966),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1361),
.B(n_841),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1345),
.B(n_841),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1378),
.B(n_968),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1311),
.B(n_972),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1508),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1501),
.A2(n_867),
.B1(n_870),
.B2(n_868),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1314),
.B(n_977),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1351),
.A2(n_876),
.B(n_877),
.C(n_873),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1382),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1381),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1370),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_L g1644 ( 
.A(n_1326),
.B(n_985),
.C(n_984),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1380),
.B(n_881),
.Y(n_1645)
);

INVx5_ASAP7_75t_L g1646 ( 
.A(n_1498),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1303),
.B(n_889),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1308),
.B(n_986),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1329),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1426),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1321),
.B(n_988),
.Y(n_1651)
);

INVx5_ASAP7_75t_L g1652 ( 
.A(n_1499),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1373),
.A2(n_895),
.B1(n_896),
.B2(n_890),
.Y(n_1653)
);

AND2x6_ASAP7_75t_L g1654 ( 
.A(n_1499),
.B(n_897),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1414),
.A2(n_1003),
.B1(n_1009),
.B2(n_1001),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1386),
.A2(n_908),
.B1(n_909),
.B2(n_900),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1340),
.A2(n_917),
.B1(n_920),
.B2(n_912),
.Y(n_1657)
);

NAND2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1338),
.B(n_921),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1328),
.B(n_843),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1385),
.B(n_1011),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1437),
.Y(n_1661)
);

AND2x6_ASAP7_75t_L g1662 ( 
.A(n_1374),
.B(n_923),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1411),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1384),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1429),
.B(n_1014),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1408),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1409),
.Y(n_1667)
);

AND2x4_ASAP7_75t_SL g1668 ( 
.A(n_1331),
.B(n_843),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1346),
.B(n_1019),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1315),
.B(n_1322),
.Y(n_1670)
);

AND3x1_ASAP7_75t_SL g1671 ( 
.A(n_1435),
.B(n_927),
.C(n_925),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1439),
.A2(n_943),
.B1(n_947),
.B2(n_930),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1363),
.B(n_843),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1327),
.A2(n_952),
.B(n_950),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1342),
.B(n_1021),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1335),
.A2(n_964),
.B(n_959),
.Y(n_1676)
);

AND2x6_ASAP7_75t_SL g1677 ( 
.A(n_1388),
.B(n_967),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1354),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1458),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1454),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1456),
.A2(n_971),
.B1(n_973),
.B2(n_969),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1357),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1358),
.Y(n_1683)
);

NAND2x1p5_ASAP7_75t_L g1684 ( 
.A(n_1339),
.B(n_975),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1410),
.B(n_1022),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1437),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1323),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1484),
.A2(n_993),
.B1(n_994),
.B2(n_989),
.Y(n_1688)
);

INVx5_ASAP7_75t_L g1689 ( 
.A(n_1415),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1422),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1488),
.A2(n_1495),
.B1(n_1392),
.B2(n_1401),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1443),
.A2(n_1502),
.B1(n_1431),
.B2(n_1330),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1341),
.A2(n_1030),
.B1(n_1031),
.B2(n_1026),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1446),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1368),
.B(n_1004),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1432),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1433),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1352),
.A2(n_1033),
.B1(n_1037),
.B2(n_1032),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1416),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1418),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1438),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1421),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1362),
.B(n_1040),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1369),
.B(n_1007),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1425),
.A2(n_1013),
.B1(n_1015),
.B2(n_1012),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1383),
.B(n_1045),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1440),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1441),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1430),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1389),
.B(n_1018),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1424),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1427),
.Y(n_1712)
);

BUFx8_ASAP7_75t_L g1713 ( 
.A(n_1343),
.Y(n_1713)
);

INVx5_ASAP7_75t_L g1714 ( 
.A(n_1437),
.Y(n_1714)
);

NOR2xp67_ASAP7_75t_L g1715 ( 
.A(n_1366),
.B(n_21),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1457),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1436),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1393),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1459),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1413),
.B(n_871),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1449),
.Y(n_1721)
);

NOR2x1p5_ASAP7_75t_L g1722 ( 
.A(n_1398),
.B(n_1400),
.Y(n_1722)
);

BUFx12f_ASAP7_75t_L g1723 ( 
.A(n_1442),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1445),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1429),
.B(n_871),
.Y(n_1725)
);

AND2x6_ASAP7_75t_L g1726 ( 
.A(n_1403),
.B(n_1036),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1448),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1420),
.B(n_1039),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1444),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1298),
.A2(n_1395),
.B1(n_1423),
.B2(n_1460),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1451),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1455),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1404),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1452),
.B(n_953),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1450),
.B(n_953),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1306),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1297),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1306),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1355),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1506),
.B(n_28),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1350),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1297),
.Y(n_1742)
);

BUFx4f_ASAP7_75t_L g1743 ( 
.A(n_1310),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1297),
.Y(n_1744)
);

BUFx12f_ASAP7_75t_L g1745 ( 
.A(n_1477),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1417),
.B(n_30),
.C(n_32),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1304),
.B(n_33),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1477),
.B(n_1119),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1310),
.B(n_33),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1334),
.Y(n_1750)
);

INVx5_ASAP7_75t_L g1751 ( 
.A(n_1310),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1297),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1297),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1336),
.A2(n_1120),
.B1(n_1126),
.B2(n_1119),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1390),
.A2(n_573),
.B(n_572),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1304),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1723),
.Y(n_1757)
);

OR2x6_ASAP7_75t_L g1758 ( 
.A(n_1745),
.B(n_34),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1756),
.B(n_36),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1530),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1580),
.A2(n_575),
.B(n_574),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1590),
.A2(n_1126),
.B1(n_1127),
.B2(n_1120),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1586),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1591),
.A2(n_1126),
.B1(n_1127),
.B2(n_1120),
.Y(n_1764)
);

BUFx5_ASAP7_75t_L g1765 ( 
.A(n_1654),
.Y(n_1765)
);

INVx5_ASAP7_75t_L g1766 ( 
.A(n_1522),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1549),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1563),
.B(n_38),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1561),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1661),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1524),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1751),
.B(n_40),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1512),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1585),
.B(n_41),
.Y(n_1774)
);

AOI21xp33_ASAP7_75t_L g1775 ( 
.A1(n_1520),
.A2(n_41),
.B(n_42),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1601),
.B(n_44),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1604),
.B(n_44),
.Y(n_1777)
);

AO32x1_ASAP7_75t_L g1778 ( 
.A1(n_1546),
.A2(n_1132),
.A3(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1620),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1605),
.B(n_48),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1666),
.B(n_49),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1519),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_R g1783 ( 
.A(n_1573),
.B(n_49),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1623),
.B(n_53),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1553),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1751),
.B(n_54),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1586),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1743),
.B(n_1751),
.Y(n_1788)
);

AND2x6_ASAP7_75t_L g1789 ( 
.A(n_1522),
.B(n_55),
.Y(n_1789)
);

NOR2x1_ASAP7_75t_L g1790 ( 
.A(n_1536),
.B(n_56),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1743),
.B(n_56),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1578),
.B(n_57),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1532),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1661),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1596),
.Y(n_1795)
);

INVx6_ASAP7_75t_L g1796 ( 
.A(n_1524),
.Y(n_1796)
);

AOI33xp33_ASAP7_75t_L g1797 ( 
.A1(n_1638),
.A2(n_61),
.A3(n_63),
.B1(n_58),
.B2(n_59),
.B3(n_62),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1670),
.A2(n_65),
.B(n_62),
.C(n_64),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1721),
.A2(n_67),
.B(n_64),
.C(n_66),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1629),
.B(n_66),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1558),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1686),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1512),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1513),
.B(n_1736),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1538),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1737),
.B(n_68),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1738),
.B(n_1600),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1523),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1603),
.B(n_70),
.Y(n_1809)
);

BUFx4f_ASAP7_75t_L g1810 ( 
.A(n_1565),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1514),
.B(n_72),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1527),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1737),
.B(n_72),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1742),
.B(n_74),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1742),
.B(n_74),
.Y(n_1815)
);

AOI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1755),
.A2(n_580),
.B(n_579),
.Y(n_1816)
);

INVx2_ASAP7_75t_SL g1817 ( 
.A(n_1741),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1543),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1526),
.B(n_76),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_SL g1820 ( 
.A(n_1659),
.B(n_76),
.C(n_77),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1721),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1522),
.B(n_79),
.Y(n_1822)
);

O2A1O1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1640),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1528),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1663),
.B(n_82),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1744),
.A2(n_87),
.B1(n_84),
.B2(n_86),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1547),
.Y(n_1827)
);

CKINVDCx14_ASAP7_75t_R g1828 ( 
.A(n_1565),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1744),
.B(n_86),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1752),
.B(n_89),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1752),
.B(n_89),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1753),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1566),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1525),
.B(n_91),
.Y(n_1834)
);

O2A1O1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1656),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1835)
);

O2A1O1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1657),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1699),
.B(n_94),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1749),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_SL g1839 ( 
.A(n_1672),
.B(n_96),
.C(n_97),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1608),
.B(n_98),
.Y(n_1840)
);

AO21x1_ASAP7_75t_L g1841 ( 
.A1(n_1716),
.A2(n_588),
.B(n_587),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1531),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1739),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1686),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1518),
.B(n_1540),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1747),
.B(n_100),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1541),
.B(n_102),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1589),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1545),
.Y(n_1849)
);

BUFx8_ASAP7_75t_L g1850 ( 
.A(n_1587),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1548),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1551),
.Y(n_1852)
);

A2O1A1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1731),
.A2(n_1694),
.B(n_1674),
.C(n_1676),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1718),
.B(n_1533),
.Y(n_1854)
);

OR2x6_ASAP7_75t_L g1855 ( 
.A(n_1537),
.B(n_105),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1687),
.B(n_105),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1750),
.A2(n_109),
.B1(n_106),
.B2(n_108),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1713),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1641),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1552),
.B(n_106),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_SL g1861 ( 
.A(n_1681),
.B(n_108),
.C(n_110),
.Y(n_1861)
);

OAI22x1_ASAP7_75t_L g1862 ( 
.A1(n_1749),
.A2(n_113),
.B1(n_110),
.B2(n_111),
.Y(n_1862)
);

INVxp67_ASAP7_75t_L g1863 ( 
.A(n_1700),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1521),
.A2(n_114),
.B1(n_111),
.B2(n_113),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1664),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_SL g1866 ( 
.A(n_1713),
.B(n_1610),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1686),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1650),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1684),
.B(n_117),
.Y(n_1869)
);

BUFx8_ASAP7_75t_L g1870 ( 
.A(n_1595),
.Y(n_1870)
);

AO21x1_ASAP7_75t_L g1871 ( 
.A1(n_1716),
.A2(n_599),
.B(n_595),
.Y(n_1871)
);

A2O1A1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1731),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_1872)
);

NAND2x1p5_ASAP7_75t_L g1873 ( 
.A(n_1630),
.B(n_119),
.Y(n_1873)
);

AO31x2_ASAP7_75t_L g1874 ( 
.A1(n_1575),
.A2(n_1719),
.A3(n_1733),
.B(n_1679),
.Y(n_1874)
);

A2O1A1Ixp33_ASAP7_75t_L g1875 ( 
.A1(n_1614),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1724),
.Y(n_1876)
);

O2A1O1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1710),
.A2(n_125),
.B(n_120),
.C(n_124),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1643),
.B(n_124),
.Y(n_1878)
);

OAI22x1_ASAP7_75t_L g1879 ( 
.A1(n_1542),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1535),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1606),
.B(n_131),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1649),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1691),
.A2(n_1693),
.B1(n_1577),
.B2(n_1655),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1582),
.B(n_133),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1727),
.Y(n_1885)
);

BUFx12f_ASAP7_75t_L g1886 ( 
.A(n_1593),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1516),
.B(n_1712),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1556),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1714),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1568),
.B(n_134),
.Y(n_1890)
);

INVx6_ASAP7_75t_L g1891 ( 
.A(n_1689),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1610),
.Y(n_1892)
);

OAI21xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1567),
.A2(n_134),
.B(n_135),
.Y(n_1893)
);

OAI22x1_ASAP7_75t_L g1894 ( 
.A1(n_1740),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1653),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.Y(n_1895)
);

OAI22x1_ASAP7_75t_L g1896 ( 
.A1(n_1554),
.A2(n_142),
.B1(n_139),
.B2(n_141),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_SL g1897 ( 
.A1(n_1616),
.A2(n_1733),
.B(n_1665),
.C(n_1725),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1654),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1714),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1714),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1562),
.A2(n_603),
.B(n_602),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1612),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1597),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1711),
.B(n_145),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1617),
.B(n_145),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1515),
.A2(n_605),
.B(n_604),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1631),
.Y(n_1907)
);

OAI22x1_ASAP7_75t_L g1908 ( 
.A1(n_1559),
.A2(n_149),
.B1(n_146),
.B2(n_148),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1717),
.B(n_146),
.Y(n_1909)
);

A2O1A1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1707),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1569),
.B(n_150),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1667),
.Y(n_1912)
);

AOI221x1_ASAP7_75t_L g1913 ( 
.A1(n_1732),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1646),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1624),
.B(n_1544),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1544),
.B(n_152),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1570),
.A2(n_612),
.B(n_610),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_SL g1918 ( 
.A(n_1644),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1579),
.A2(n_614),
.B(n_613),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1534),
.Y(n_1920)
);

BUFx4f_ASAP7_75t_L g1921 ( 
.A(n_1645),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1646),
.Y(n_1922)
);

OAI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1594),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1637),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1729),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1574),
.B(n_156),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1633),
.B(n_157),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1702),
.B(n_158),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1571),
.B(n_158),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1689),
.Y(n_1930)
);

NOR3xp33_ASAP7_75t_L g1931 ( 
.A(n_1634),
.B(n_159),
.C(n_160),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1534),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1534),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1709),
.Y(n_1934)
);

O2A1O1Ixp33_ASAP7_75t_L g1935 ( 
.A1(n_1685),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1654),
.Y(n_1936)
);

CKINVDCx11_ASAP7_75t_R g1937 ( 
.A(n_1677),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1615),
.B(n_162),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1615),
.B(n_163),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1654),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1607),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1599),
.A2(n_618),
.B(n_617),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1635),
.A2(n_620),
.B(n_619),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1572),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1611),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1588),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1675),
.A2(n_623),
.B(n_621),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1636),
.A2(n_625),
.B(n_624),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1748),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1621),
.A2(n_167),
.B1(n_164),
.B2(n_166),
.Y(n_1950)
);

OR2x6_ASAP7_75t_L g1951 ( 
.A(n_1748),
.B(n_166),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1645),
.Y(n_1952)
);

CKINVDCx8_ASAP7_75t_R g1953 ( 
.A(n_1645),
.Y(n_1953)
);

AO32x1_ASAP7_75t_L g1954 ( 
.A1(n_1688),
.A2(n_169),
.A3(n_167),
.B1(n_168),
.B2(n_171),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1639),
.A2(n_631),
.B(n_628),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1628),
.A2(n_175),
.B1(n_172),
.B2(n_174),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1692),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1728),
.B(n_178),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1645),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1576),
.A2(n_639),
.B(n_637),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1652),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1697),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1660),
.A2(n_642),
.B(n_640),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1588),
.B(n_179),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1626),
.B(n_179),
.Y(n_1965)
);

O2A1O1Ixp33_ASAP7_75t_L g1966 ( 
.A1(n_1555),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1966)
);

A2O1A1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1715),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1651),
.A2(n_648),
.B(n_645),
.Y(n_1968)
);

O2A1O1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1557),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_1969)
);

XNOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1698),
.B(n_185),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1539),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1626),
.B(n_186),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_SL g1973 ( 
.A(n_1588),
.B(n_187),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1673),
.B(n_187),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1746),
.B(n_188),
.C(n_189),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1517),
.B(n_189),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1648),
.B(n_190),
.Y(n_1977)
);

BUFx3_ASAP7_75t_L g1978 ( 
.A(n_1689),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1613),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1622),
.B(n_191),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1613),
.B(n_194),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1705),
.B(n_198),
.Y(n_1982)
);

INVxp67_ASAP7_75t_L g1983 ( 
.A(n_1662),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1662),
.B(n_198),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1662),
.B(n_199),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1730),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1702),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1625),
.Y(n_1988)
);

BUFx12f_ASAP7_75t_L g1989 ( 
.A(n_1627),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1613),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1609),
.B(n_205),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1632),
.B(n_206),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1602),
.B(n_208),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1642),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1627),
.B(n_209),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1690),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_SL g1997 ( 
.A(n_1529),
.B(n_211),
.C(n_212),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1690),
.Y(n_1998)
);

INVxp33_ASAP7_75t_SL g1999 ( 
.A(n_1669),
.Y(n_1999)
);

INVx3_ASAP7_75t_SL g2000 ( 
.A(n_1668),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1696),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1618),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1581),
.A2(n_655),
.B(n_654),
.Y(n_2003)
);

A2O1A1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1735),
.A2(n_1706),
.B(n_1696),
.C(n_1647),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1583),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1678),
.Y(n_2006)
);

NOR2xp67_ASAP7_75t_SL g2007 ( 
.A(n_1560),
.B(n_1701),
.Y(n_2007)
);

A2O1A1Ixp33_ASAP7_75t_L g2008 ( 
.A1(n_1619),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1682),
.Y(n_2009)
);

BUFx2_ASAP7_75t_L g2010 ( 
.A(n_1726),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1695),
.B(n_221),
.Y(n_2011)
);

A2O1A1Ixp33_ASAP7_75t_L g2012 ( 
.A1(n_1754),
.A2(n_1703),
.B(n_1683),
.C(n_1695),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1720),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1708),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1658),
.B(n_222),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1726),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1704),
.B(n_223),
.Y(n_2017)
);

OAI22x1_ASAP7_75t_L g2018 ( 
.A1(n_1671),
.A2(n_1734),
.B1(n_1584),
.B2(n_1592),
.Y(n_2018)
);

INVx5_ASAP7_75t_L g2019 ( 
.A(n_1618),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1726),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1726),
.Y(n_2021)
);

NOR2x1_ASAP7_75t_L g2022 ( 
.A(n_1722),
.B(n_229),
.Y(n_2022)
);

BUFx8_ASAP7_75t_L g2023 ( 
.A(n_1680),
.Y(n_2023)
);

INVx5_ASAP7_75t_L g2024 ( 
.A(n_1723),
.Y(n_2024)
);

O2A1O1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1550),
.A2(n_236),
.B(n_233),
.C(n_235),
.Y(n_2025)
);

NOR2xp67_ASAP7_75t_L g2026 ( 
.A(n_1745),
.B(n_235),
.Y(n_2026)
);

AO32x1_ASAP7_75t_L g2027 ( 
.A1(n_1546),
.A2(n_240),
.A3(n_237),
.B1(n_238),
.B2(n_242),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1756),
.B(n_237),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1530),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1561),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1756),
.B(n_240),
.Y(n_2031)
);

NAND2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1524),
.B(n_242),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1756),
.B(n_243),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1756),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2034)
);

A2O1A1Ixp33_ASAP7_75t_SL g2035 ( 
.A1(n_1598),
.A2(n_664),
.B(n_665),
.C(n_662),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1563),
.B(n_244),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1756),
.B(n_245),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1563),
.B(n_246),
.Y(n_2038)
);

NOR2x1_ASAP7_75t_L g2039 ( 
.A(n_1564),
.B(n_247),
.Y(n_2039)
);

NOR3xp33_ASAP7_75t_L g2040 ( 
.A(n_1691),
.B(n_248),
.C(n_249),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1661),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1756),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1530),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_SL g2044 ( 
.A1(n_1586),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2044)
);

O2A1O1Ixp33_ASAP7_75t_L g2045 ( 
.A1(n_1550),
.A2(n_254),
.B(n_251),
.C(n_253),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1563),
.B(n_255),
.Y(n_2046)
);

INVxp67_ASAP7_75t_SL g2047 ( 
.A(n_1756),
.Y(n_2047)
);

AOI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_1756),
.A2(n_259),
.B1(n_256),
.B2(n_257),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_L g2049 ( 
.A(n_1661),
.B(n_669),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1723),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1580),
.A2(n_671),
.B(n_670),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1563),
.B(n_256),
.Y(n_2052)
);

INVx4_ASAP7_75t_L g2053 ( 
.A(n_1745),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1756),
.A2(n_262),
.B1(n_257),
.B2(n_261),
.Y(n_2054)
);

CKINVDCx20_ASAP7_75t_R g2055 ( 
.A(n_1561),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1756),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1580),
.A2(n_676),
.B(n_674),
.Y(n_2057)
);

NAND2x1p5_ASAP7_75t_L g2058 ( 
.A(n_1524),
.B(n_265),
.Y(n_2058)
);

AOI33xp33_ASAP7_75t_L g2059 ( 
.A1(n_1638),
.A2(n_267),
.A3(n_268),
.B1(n_270),
.B2(n_271),
.B3(n_272),
.Y(n_2059)
);

O2A1O1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_1550),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1580),
.A2(n_679),
.B(n_273),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1756),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1756),
.B(n_274),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_1563),
.B(n_277),
.Y(n_2064)
);

BUFx4f_ASAP7_75t_SL g2065 ( 
.A(n_1745),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_1743),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1756),
.B(n_277),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_SL g2068 ( 
.A(n_1745),
.B(n_278),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1745),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1580),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1756),
.B(n_279),
.Y(n_2071)
);

A2O1A1Ixp33_ASAP7_75t_L g2072 ( 
.A1(n_1580),
.A2(n_283),
.B(n_281),
.C(n_282),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_SL g2073 ( 
.A(n_1745),
.B(n_281),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1756),
.B(n_283),
.Y(n_2074)
);

INVx4_ASAP7_75t_L g2075 ( 
.A(n_1745),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_1561),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1756),
.B(n_284),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_SL g2078 ( 
.A1(n_1586),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2078)
);

OAI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1756),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_1580),
.A2(n_287),
.B(n_291),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1756),
.B(n_292),
.Y(n_2081)
);

INVx5_ASAP7_75t_L g2082 ( 
.A(n_1723),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1563),
.B(n_293),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1580),
.A2(n_294),
.B(n_295),
.Y(n_2084)
);

O2A1O1Ixp5_ASAP7_75t_L g2085 ( 
.A1(n_1725),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1530),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1756),
.B(n_296),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1563),
.B(n_297),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1756),
.B(n_297),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1756),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_R g2091 ( 
.A(n_1573),
.B(n_299),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_R g2092 ( 
.A(n_1573),
.B(n_299),
.Y(n_2092)
);

OAI221xp5_ASAP7_75t_L g2093 ( 
.A1(n_1550),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.C(n_304),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1756),
.B(n_302),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1745),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1756),
.B(n_304),
.Y(n_2096)
);

NOR3xp33_ASAP7_75t_SL g2097 ( 
.A(n_1573),
.B(n_305),
.C(n_306),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1530),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1756),
.B(n_305),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1580),
.A2(n_307),
.B(n_308),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1756),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1563),
.B(n_307),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1745),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_R g2104 ( 
.A(n_1573),
.B(n_309),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1563),
.B(n_310),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1756),
.B(n_312),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1756),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1530),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_1723),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_1745),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1756),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2111)
);

OAI22x1_ASAP7_75t_L g2112 ( 
.A1(n_1749),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_SL g2113 ( 
.A1(n_1586),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_2113)
);

OAI21xp33_ASAP7_75t_L g2114 ( 
.A1(n_1550),
.A2(n_322),
.B(n_323),
.Y(n_2114)
);

O2A1O1Ixp33_ASAP7_75t_L g2115 ( 
.A1(n_1550),
.A2(n_325),
.B(n_322),
.C(n_323),
.Y(n_2115)
);

AOI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_1580),
.A2(n_328),
.B(n_329),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1745),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1756),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_1563),
.B(n_331),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1756),
.B(n_331),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1563),
.B(n_332),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1756),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1756),
.B(n_333),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1756),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_1563),
.B(n_334),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1756),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_1756),
.Y(n_2127)
);

A2O1A1Ixp33_ASAP7_75t_L g2128 ( 
.A1(n_1580),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1580),
.A2(n_337),
.B(n_339),
.Y(n_2129)
);

BUFx5_ASAP7_75t_L g2130 ( 
.A(n_1789),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2047),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2131)
);

HB1xp67_ASAP7_75t_L g2132 ( 
.A(n_2127),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2056),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1854),
.B(n_341),
.Y(n_2134)
);

OAI21x1_ASAP7_75t_SL g2135 ( 
.A1(n_1761),
.A2(n_342),
.B(n_343),
.Y(n_2135)
);

BUFx5_ASAP7_75t_L g2136 ( 
.A(n_1789),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_1863),
.B(n_344),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1773),
.Y(n_2138)
);

BUFx3_ASAP7_75t_L g2139 ( 
.A(n_1757),
.Y(n_2139)
);

INVxp67_ASAP7_75t_SL g2140 ( 
.A(n_2094),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_1757),
.Y(n_2141)
);

AO21x2_ASAP7_75t_L g2142 ( 
.A1(n_1816),
.A2(n_347),
.B(n_348),
.Y(n_2142)
);

INVx4_ASAP7_75t_L g2143 ( 
.A(n_1757),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_1810),
.Y(n_2144)
);

OR2x6_ASAP7_75t_L g2145 ( 
.A(n_1951),
.B(n_349),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_SL g2146 ( 
.A1(n_1828),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_2146)
);

AOI22x1_ASAP7_75t_L g2147 ( 
.A1(n_2018),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_2094),
.Y(n_2148)
);

INVx3_ASAP7_75t_SL g2149 ( 
.A(n_2053),
.Y(n_2149)
);

OAI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_1853),
.A2(n_355),
.B(n_357),
.Y(n_2150)
);

INVxp67_ASAP7_75t_SL g2151 ( 
.A(n_1830),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2090),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_2024),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1953),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_2024),
.Y(n_2155)
);

AO21x2_ASAP7_75t_L g2156 ( 
.A1(n_1841),
.A2(n_360),
.B(n_362),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1832),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_1845),
.B(n_362),
.Y(n_2158)
);

BUFx2_ASAP7_75t_R g2159 ( 
.A(n_2095),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_2024),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_2082),
.Y(n_2161)
);

INVx1_ASAP7_75t_SL g2162 ( 
.A(n_1793),
.Y(n_2162)
);

INVx4_ASAP7_75t_L g2163 ( 
.A(n_2082),
.Y(n_2163)
);

INVx4_ASAP7_75t_L g2164 ( 
.A(n_2082),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2101),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2107),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2118),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1915),
.B(n_366),
.Y(n_2168)
);

BUFx2_ASAP7_75t_L g2169 ( 
.A(n_1810),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_1801),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2122),
.B(n_367),
.Y(n_2171)
);

AO21x2_ASAP7_75t_L g2172 ( 
.A1(n_1871),
.A2(n_367),
.B(n_368),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_1951),
.Y(n_2173)
);

AOI22x1_ASAP7_75t_L g2174 ( 
.A1(n_1943),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2126),
.Y(n_2175)
);

AO21x2_ASAP7_75t_L g2176 ( 
.A1(n_1906),
.A2(n_371),
.B(n_372),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2012),
.A2(n_373),
.B(n_374),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1889),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1785),
.Y(n_2179)
);

AOI22x1_ASAP7_75t_L g2180 ( 
.A1(n_1963),
.A2(n_1968),
.B1(n_1917),
.B2(n_1919),
.Y(n_2180)
);

OA21x2_ASAP7_75t_L g2181 ( 
.A1(n_1913),
.A2(n_373),
.B(n_375),
.Y(n_2181)
);

AO21x1_ASAP7_75t_L g2182 ( 
.A1(n_2025),
.A2(n_375),
.B(n_377),
.Y(n_2182)
);

INVxp67_ASAP7_75t_SL g2183 ( 
.A(n_1830),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_2065),
.Y(n_2184)
);

BUFx12f_ASAP7_75t_L g2185 ( 
.A(n_2053),
.Y(n_2185)
);

NAND2x1p5_ASAP7_75t_L g2186 ( 
.A(n_1921),
.B(n_380),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_1889),
.Y(n_2187)
);

INVxp67_ASAP7_75t_SL g2188 ( 
.A(n_1831),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1848),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_2069),
.Y(n_2190)
);

CKINVDCx11_ASAP7_75t_R g2191 ( 
.A(n_2000),
.Y(n_2191)
);

BUFx4f_ASAP7_75t_L g2192 ( 
.A(n_1758),
.Y(n_2192)
);

INVx1_ASAP7_75t_SL g2193 ( 
.A(n_1903),
.Y(n_2193)
);

AOI22x1_ASAP7_75t_L g2194 ( 
.A1(n_1901),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_2103),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_SL g2196 ( 
.A1(n_1831),
.A2(n_383),
.B1(n_385),
.B2(n_387),
.Y(n_2196)
);

BUFx3_ASAP7_75t_L g2197 ( 
.A(n_2023),
.Y(n_2197)
);

INVxp67_ASAP7_75t_SL g2198 ( 
.A(n_1928),
.Y(n_2198)
);

INVx5_ASAP7_75t_L g2199 ( 
.A(n_1789),
.Y(n_2199)
);

OAI21x1_ASAP7_75t_SL g2200 ( 
.A1(n_2039),
.A2(n_385),
.B(n_388),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_2030),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_2051),
.A2(n_2057),
.B(n_1942),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_L g2203 ( 
.A1(n_1947),
.A2(n_1955),
.B(n_1948),
.Y(n_2203)
);

NAND2x1p5_ASAP7_75t_L g2204 ( 
.A(n_1921),
.B(n_2019),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1852),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1808),
.Y(n_2206)
);

AO21x2_ASAP7_75t_L g2207 ( 
.A1(n_2114),
.A2(n_389),
.B(n_390),
.Y(n_2207)
);

AO21x2_ASAP7_75t_L g2208 ( 
.A1(n_1806),
.A2(n_389),
.B(n_391),
.Y(n_2208)
);

OAI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2004),
.A2(n_391),
.B(n_392),
.Y(n_2209)
);

OAI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_1759),
.A2(n_392),
.B(n_393),
.Y(n_2210)
);

AO21x2_ASAP7_75t_L g2211 ( 
.A1(n_1813),
.A2(n_393),
.B(n_394),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1999),
.B(n_394),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1760),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_1887),
.B(n_395),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_1881),
.A2(n_395),
.B(n_396),
.Y(n_2215)
);

AO21x2_ASAP7_75t_L g2216 ( 
.A1(n_1814),
.A2(n_397),
.B(n_399),
.Y(n_2216)
);

BUFx2_ASAP7_75t_L g2217 ( 
.A(n_1787),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_2003),
.A2(n_397),
.B(n_400),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_2023),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2040),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_2220)
);

AOI21x1_ASAP7_75t_L g2221 ( 
.A1(n_1973),
.A2(n_401),
.B(n_402),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1824),
.Y(n_2222)
);

BUFx5_ASAP7_75t_L g2223 ( 
.A(n_1789),
.Y(n_2223)
);

OAI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2028),
.A2(n_2033),
.B(n_2031),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1849),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1889),
.Y(n_2226)
);

BUFx12f_ASAP7_75t_L g2227 ( 
.A(n_2075),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_2110),
.Y(n_2228)
);

AO21x2_ASAP7_75t_L g2229 ( 
.A1(n_1815),
.A2(n_403),
.B(n_404),
.Y(n_2229)
);

AO21x2_ASAP7_75t_L g2230 ( 
.A1(n_1829),
.A2(n_404),
.B(n_405),
.Y(n_2230)
);

AOI22x1_ASAP7_75t_L g2231 ( 
.A1(n_2061),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_2231)
);

AND2x4_ASAP7_75t_L g2232 ( 
.A(n_2019),
.B(n_407),
.Y(n_2232)
);

BUFx8_ASAP7_75t_L g2233 ( 
.A(n_1805),
.Y(n_2233)
);

OAI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2037),
.A2(n_408),
.B(n_409),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2017),
.B(n_1811),
.Y(n_2235)
);

BUFx2_ASAP7_75t_SL g2236 ( 
.A(n_2117),
.Y(n_2236)
);

BUFx2_ASAP7_75t_R g2237 ( 
.A(n_1858),
.Y(n_2237)
);

NAND2x1p5_ASAP7_75t_L g2238 ( 
.A(n_2019),
.B(n_410),
.Y(n_2238)
);

BUFx3_ASAP7_75t_L g2239 ( 
.A(n_1766),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_1766),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1766),
.Y(n_2241)
);

BUFx2_ASAP7_75t_SL g2242 ( 
.A(n_2075),
.Y(n_2242)
);

AO21x2_ASAP7_75t_L g2243 ( 
.A1(n_2074),
.A2(n_2120),
.B(n_2096),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1771),
.B(n_551),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1899),
.Y(n_2245)
);

BUFx8_ASAP7_75t_L g2246 ( 
.A(n_1886),
.Y(n_2246)
);

AOI22x1_ASAP7_75t_L g2247 ( 
.A1(n_1960),
.A2(n_1894),
.B1(n_1908),
.B2(n_2080),
.Y(n_2247)
);

CKINVDCx20_ASAP7_75t_R g2248 ( 
.A(n_2055),
.Y(n_2248)
);

BUFx10_ASAP7_75t_L g2249 ( 
.A(n_1758),
.Y(n_2249)
);

OA21x2_ASAP7_75t_L g2250 ( 
.A1(n_2085),
.A2(n_410),
.B(n_411),
.Y(n_2250)
);

AOI21x1_ASAP7_75t_L g2251 ( 
.A1(n_1822),
.A2(n_411),
.B(n_412),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_1792),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1851),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2017),
.B(n_413),
.Y(n_2254)
);

NOR2x1_ASAP7_75t_R g2255 ( 
.A(n_1769),
.B(n_415),
.Y(n_2255)
);

BUFx3_ASAP7_75t_L g2256 ( 
.A(n_1899),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1934),
.Y(n_2257)
);

AOI22x1_ASAP7_75t_L g2258 ( 
.A1(n_2129),
.A2(n_416),
.B1(n_417),
.B2(n_419),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1859),
.Y(n_2259)
);

OA21x2_ASAP7_75t_L g2260 ( 
.A1(n_1799),
.A2(n_417),
.B(n_419),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1971),
.Y(n_2261)
);

NAND2x1p5_ASAP7_75t_L g2262 ( 
.A(n_1952),
.B(n_420),
.Y(n_2262)
);

NAND2x1p5_ASAP7_75t_L g2263 ( 
.A(n_1959),
.B(n_422),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1888),
.Y(n_2264)
);

INVx4_ASAP7_75t_L g2265 ( 
.A(n_1771),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_1790),
.A2(n_424),
.B(n_425),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_1899),
.Y(n_2267)
);

OA21x2_ASAP7_75t_L g2268 ( 
.A1(n_1821),
.A2(n_426),
.B(n_427),
.Y(n_2268)
);

BUFx2_ASAP7_75t_L g2269 ( 
.A(n_1898),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_SL g2270 ( 
.A1(n_1790),
.A2(n_427),
.B(n_428),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1876),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1885),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2029),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2043),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2086),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_1900),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2098),
.Y(n_2277)
);

BUFx12f_ASAP7_75t_L g2278 ( 
.A(n_1812),
.Y(n_2278)
);

BUFx2_ASAP7_75t_L g2279 ( 
.A(n_1936),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_1900),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_1900),
.Y(n_2281)
);

AO21x2_ASAP7_75t_L g2282 ( 
.A1(n_2123),
.A2(n_428),
.B(n_429),
.Y(n_2282)
);

AO21x2_ASAP7_75t_L g2283 ( 
.A1(n_2035),
.A2(n_430),
.B(n_431),
.Y(n_2283)
);

BUFx2_ASAP7_75t_R g2284 ( 
.A(n_1795),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_1870),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_1834),
.A2(n_431),
.B(n_432),
.Y(n_2286)
);

BUFx2_ASAP7_75t_SL g2287 ( 
.A(n_2076),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2108),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_1928),
.Y(n_2289)
);

BUFx4f_ASAP7_75t_SL g2290 ( 
.A(n_1850),
.Y(n_2290)
);

BUFx2_ASAP7_75t_R g2291 ( 
.A(n_1818),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_1975),
.A2(n_432),
.B1(n_433),
.B2(n_434),
.Y(n_2292)
);

AOI22x1_ASAP7_75t_L g2293 ( 
.A1(n_2084),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_1922),
.Y(n_2294)
);

OAI21x1_ASAP7_75t_L g2295 ( 
.A1(n_1964),
.A2(n_435),
.B(n_436),
.Y(n_2295)
);

BUFx12f_ASAP7_75t_L g2296 ( 
.A(n_1850),
.Y(n_2296)
);

AO21x2_ASAP7_75t_L g2297 ( 
.A1(n_1839),
.A2(n_437),
.B(n_438),
.Y(n_2297)
);

INVx6_ASAP7_75t_L g2298 ( 
.A(n_1870),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2067),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_1869),
.B(n_438),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2077),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1868),
.B(n_439),
.Y(n_2302)
);

OAI21x1_ASAP7_75t_L g2303 ( 
.A1(n_1981),
.A2(n_1764),
.B(n_1762),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_1907),
.B(n_440),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_1914),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1924),
.Y(n_2306)
);

INVx1_ASAP7_75t_SL g2307 ( 
.A(n_1882),
.Y(n_2307)
);

NAND2x1_ASAP7_75t_L g2308 ( 
.A(n_1920),
.B(n_443),
.Y(n_2308)
);

INVx6_ASAP7_75t_L g2309 ( 
.A(n_1827),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1767),
.Y(n_2310)
);

AO21x2_ASAP7_75t_L g2311 ( 
.A1(n_1861),
.A2(n_443),
.B(n_444),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1800),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1800),
.Y(n_2313)
);

BUFx4f_ASAP7_75t_L g2314 ( 
.A(n_1855),
.Y(n_2314)
);

BUFx3_ASAP7_75t_L g2315 ( 
.A(n_2050),
.Y(n_2315)
);

INVx5_ASAP7_75t_L g2316 ( 
.A(n_1932),
.Y(n_2316)
);

OAI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2063),
.A2(n_445),
.B(n_446),
.Y(n_2317)
);

BUFx2_ASAP7_75t_L g2318 ( 
.A(n_1833),
.Y(n_2318)
);

BUFx2_ASAP7_75t_SL g2319 ( 
.A(n_2050),
.Y(n_2319)
);

BUFx12f_ASAP7_75t_L g2320 ( 
.A(n_1855),
.Y(n_2320)
);

BUFx3_ASAP7_75t_L g2321 ( 
.A(n_2109),
.Y(n_2321)
);

INVxp67_ASAP7_75t_SL g2322 ( 
.A(n_1932),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1880),
.B(n_446),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1783),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_1825),
.B(n_447),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_2109),
.Y(n_2326)
);

CKINVDCx6p67_ASAP7_75t_R g2327 ( 
.A(n_1896),
.Y(n_2327)
);

INVx2_ASAP7_75t_SL g2328 ( 
.A(n_1796),
.Y(n_2328)
);

NAND2x1p5_ASAP7_75t_L g2329 ( 
.A(n_1922),
.B(n_447),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_1961),
.Y(n_2330)
);

OR2x6_ASAP7_75t_L g2331 ( 
.A(n_1819),
.B(n_448),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_1961),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_1865),
.B(n_551),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1819),
.Y(n_2334)
);

OAI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2068),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_2335)
);

INVx5_ASAP7_75t_L g2336 ( 
.A(n_1933),
.Y(n_2336)
);

OAI21x1_ASAP7_75t_L g2337 ( 
.A1(n_1776),
.A2(n_452),
.B(n_453),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1995),
.B(n_452),
.Y(n_2338)
);

OAI21x1_ASAP7_75t_L g2339 ( 
.A1(n_1780),
.A2(n_454),
.B(n_455),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_1933),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_1796),
.Y(n_2341)
);

BUFx2_ASAP7_75t_SL g2342 ( 
.A(n_1765),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1770),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2006),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1840),
.B(n_455),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_2091),
.Y(n_2346)
);

AOI21x1_ASAP7_75t_L g2347 ( 
.A1(n_2021),
.A2(n_456),
.B(n_457),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2009),
.Y(n_2348)
);

CKINVDCx8_ASAP7_75t_R g2349 ( 
.A(n_1842),
.Y(n_2349)
);

BUFx2_ASAP7_75t_R g2350 ( 
.A(n_1970),
.Y(n_2350)
);

CKINVDCx20_ASAP7_75t_R g2351 ( 
.A(n_2092),
.Y(n_2351)
);

NAND2x1p5_ASAP7_75t_L g2352 ( 
.A(n_1940),
.B(n_1944),
.Y(n_2352)
);

OAI21x1_ASAP7_75t_L g2353 ( 
.A1(n_1784),
.A2(n_456),
.B(n_457),
.Y(n_2353)
);

OAI21x1_ASAP7_75t_L g2354 ( 
.A1(n_2100),
.A2(n_459),
.B(n_460),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_1995),
.B(n_459),
.Y(n_2355)
);

INVx8_ASAP7_75t_L g2356 ( 
.A(n_1772),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1797),
.Y(n_2357)
);

BUFx5_ASAP7_75t_L g2358 ( 
.A(n_1978),
.Y(n_2358)
);

AND2x6_ASAP7_75t_L g2359 ( 
.A(n_1946),
.B(n_460),
.Y(n_2359)
);

INVx4_ASAP7_75t_L g2360 ( 
.A(n_1946),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2001),
.B(n_550),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1770),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_1765),
.B(n_461),
.Y(n_2363)
);

INVx6_ASAP7_75t_L g2364 ( 
.A(n_1891),
.Y(n_2364)
);

INVx4_ASAP7_75t_L g2365 ( 
.A(n_1979),
.Y(n_2365)
);

INVx2_ASAP7_75t_SL g2366 ( 
.A(n_1891),
.Y(n_2366)
);

BUFx2_ASAP7_75t_L g2367 ( 
.A(n_2014),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1770),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1794),
.Y(n_2369)
);

INVx6_ASAP7_75t_L g2370 ( 
.A(n_1979),
.Y(n_2370)
);

OR2x6_ASAP7_75t_L g2371 ( 
.A(n_2032),
.B(n_462),
.Y(n_2371)
);

OAI21x1_ASAP7_75t_L g2372 ( 
.A1(n_2116),
.A2(n_464),
.B(n_465),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2059),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1794),
.Y(n_2374)
);

INVx6_ASAP7_75t_L g2375 ( 
.A(n_1990),
.Y(n_2375)
);

AO21x2_ASAP7_75t_L g2376 ( 
.A1(n_1905),
.A2(n_467),
.B(n_468),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1838),
.B(n_467),
.Y(n_2377)
);

AOI21x1_ASAP7_75t_L g2378 ( 
.A1(n_2010),
.A2(n_468),
.B(n_469),
.Y(n_2378)
);

HB1xp67_ASAP7_75t_L g2379 ( 
.A(n_1990),
.Y(n_2379)
);

OAI21x1_ASAP7_75t_SL g2380 ( 
.A1(n_1984),
.A2(n_470),
.B(n_471),
.Y(n_2380)
);

BUFx3_ASAP7_75t_L g2381 ( 
.A(n_1765),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_L g2382 ( 
.A1(n_1847),
.A2(n_472),
.B(n_473),
.Y(n_2382)
);

AOI21x1_ASAP7_75t_L g2383 ( 
.A1(n_2016),
.A2(n_472),
.B(n_473),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_1976),
.B(n_474),
.Y(n_2384)
);

BUFx12f_ASAP7_75t_L g2385 ( 
.A(n_1937),
.Y(n_2385)
);

INVx5_ASAP7_75t_SL g2386 ( 
.A(n_1772),
.Y(n_2386)
);

AND2x6_ASAP7_75t_L g2387 ( 
.A(n_1794),
.B(n_475),
.Y(n_2387)
);

OAI21x1_ASAP7_75t_L g2388 ( 
.A1(n_1935),
.A2(n_476),
.B(n_477),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_1786),
.Y(n_2389)
);

BUFx2_ASAP7_75t_R g2390 ( 
.A(n_1788),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_1962),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_2001),
.B(n_1843),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_1786),
.Y(n_2393)
);

BUFx2_ASAP7_75t_SL g2394 ( 
.A(n_1765),
.Y(n_2394)
);

INVx6_ASAP7_75t_SL g2395 ( 
.A(n_1866),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1802),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_1989),
.B(n_476),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_1949),
.Y(n_2398)
);

BUFx12f_ASAP7_75t_L g2399 ( 
.A(n_1817),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2104),
.Y(n_2400)
);

NAND2x1p5_ASAP7_75t_L g2401 ( 
.A(n_1844),
.B(n_479),
.Y(n_2401)
);

INVx8_ASAP7_75t_L g2402 ( 
.A(n_1996),
.Y(n_2402)
);

AOI22x1_ASAP7_75t_L g2403 ( 
.A1(n_1879),
.A2(n_484),
.B1(n_485),
.B2(n_486),
.Y(n_2403)
);

BUFx2_ASAP7_75t_L g2404 ( 
.A(n_1782),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1918),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_1867),
.B(n_486),
.Y(n_2406)
);

INVx2_ASAP7_75t_SL g2407 ( 
.A(n_2066),
.Y(n_2407)
);

INVx5_ASAP7_75t_L g2408 ( 
.A(n_2041),
.Y(n_2408)
);

BUFx8_ASAP7_75t_SL g2409 ( 
.A(n_1996),
.Y(n_2409)
);

AO21x2_ASAP7_75t_L g2410 ( 
.A1(n_1872),
.A2(n_487),
.B(n_488),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_1804),
.B(n_1781),
.Y(n_2411)
);

INVxp67_ASAP7_75t_SL g2412 ( 
.A(n_1873),
.Y(n_2412)
);

AO21x2_ASAP7_75t_L g2413 ( 
.A1(n_2070),
.A2(n_488),
.B(n_489),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_1998),
.Y(n_2414)
);

AO21x2_ASAP7_75t_L g2415 ( 
.A1(n_2072),
.A2(n_489),
.B(n_490),
.Y(n_2415)
);

AO21x2_ASAP7_75t_L g2416 ( 
.A1(n_2128),
.A2(n_490),
.B(n_491),
.Y(n_2416)
);

AO21x2_ASAP7_75t_L g2417 ( 
.A1(n_1798),
.A2(n_491),
.B(n_492),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2071),
.Y(n_2418)
);

INVxp67_ASAP7_75t_L g2419 ( 
.A(n_1926),
.Y(n_2419)
);

AOI22x1_ASAP7_75t_L g2420 ( 
.A1(n_1862),
.A2(n_2112),
.B1(n_2058),
.B2(n_1846),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1927),
.B(n_492),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1809),
.B(n_493),
.Y(n_2422)
);

BUFx2_ASAP7_75t_SL g2423 ( 
.A(n_2026),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_1925),
.B(n_550),
.Y(n_2424)
);

OA21x2_ASAP7_75t_L g2425 ( 
.A1(n_1910),
.A2(n_494),
.B(n_495),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2081),
.Y(n_2426)
);

CKINVDCx20_ASAP7_75t_R g2427 ( 
.A(n_1763),
.Y(n_2427)
);

OAI21x1_ASAP7_75t_SL g2428 ( 
.A1(n_1985),
.A2(n_495),
.B(n_496),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2087),
.Y(n_2429)
);

BUFx3_ASAP7_75t_L g2430 ( 
.A(n_1930),
.Y(n_2430)
);

OR2x6_ASAP7_75t_L g2431 ( 
.A(n_1892),
.B(n_497),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2089),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_1807),
.B(n_498),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_1883),
.A2(n_499),
.B1(n_501),
.B2(n_502),
.Y(n_2434)
);

BUFx10_ASAP7_75t_L g2435 ( 
.A(n_2015),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2099),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2106),
.A2(n_503),
.B(n_504),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1941),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_1912),
.Y(n_2439)
);

OAI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_1977),
.A2(n_505),
.B(n_506),
.Y(n_2440)
);

OAI21x1_ASAP7_75t_L g2441 ( 
.A1(n_2045),
.A2(n_506),
.B(n_507),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_1945),
.Y(n_2442)
);

AO21x1_ASAP7_75t_L g2443 ( 
.A1(n_2060),
.A2(n_507),
.B(n_508),
.Y(n_2443)
);

OAI21x1_ASAP7_75t_L g2444 ( 
.A1(n_2115),
.A2(n_509),
.B(n_510),
.Y(n_2444)
);

CKINVDCx20_ASAP7_75t_R g2445 ( 
.A(n_2044),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1988),
.Y(n_2446)
);

NAND2x1p5_ASAP7_75t_L g2447 ( 
.A(n_2007),
.B(n_511),
.Y(n_2447)
);

AO21x2_ASAP7_75t_L g2448 ( 
.A1(n_1967),
.A2(n_513),
.B(n_514),
.Y(n_2448)
);

AO21x2_ASAP7_75t_L g2449 ( 
.A1(n_2008),
.A2(n_515),
.B(n_516),
.Y(n_2449)
);

OAI21x1_ASAP7_75t_L g2450 ( 
.A1(n_1966),
.A2(n_515),
.B(n_517),
.Y(n_2450)
);

AO21x2_ASAP7_75t_L g2451 ( 
.A1(n_2049),
.A2(n_517),
.B(n_518),
.Y(n_2451)
);

OAI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_1884),
.A2(n_518),
.B(n_520),
.Y(n_2452)
);

OR2x2_ASAP7_75t_L g2453 ( 
.A(n_1916),
.B(n_521),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_1997),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2097),
.Y(n_2455)
);

OAI21x1_ASAP7_75t_L g2456 ( 
.A1(n_1969),
.A2(n_522),
.B(n_523),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_1837),
.B(n_522),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_1994),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2138),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2133),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2327),
.A2(n_1957),
.B1(n_1931),
.B2(n_2002),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2213),
.Y(n_2462)
);

AOI22xp33_ASAP7_75t_L g2463 ( 
.A1(n_2314),
.A2(n_2078),
.B1(n_2113),
.B2(n_1857),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2152),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2165),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2166),
.Y(n_2466)
);

HB1xp67_ASAP7_75t_L g2467 ( 
.A(n_2198),
.Y(n_2467)
);

HB1xp67_ASAP7_75t_L g2468 ( 
.A(n_2198),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2167),
.Y(n_2469)
);

INVx4_ASAP7_75t_L g2470 ( 
.A(n_2290),
.Y(n_2470)
);

AOI22xp33_ASAP7_75t_SL g2471 ( 
.A1(n_2151),
.A2(n_2073),
.B1(n_1893),
.B2(n_2093),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2316),
.Y(n_2472)
);

AOI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2151),
.A2(n_1911),
.B1(n_1895),
.B2(n_1923),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2175),
.Y(n_2474)
);

INVx4_ASAP7_75t_L g2475 ( 
.A(n_2290),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2179),
.Y(n_2476)
);

AOI21x1_ASAP7_75t_L g2477 ( 
.A1(n_2177),
.A2(n_2022),
.B(n_1878),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_2265),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2206),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2222),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2225),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2183),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2253),
.Y(n_2483)
);

INVx3_ASAP7_75t_SL g2484 ( 
.A(n_2228),
.Y(n_2484)
);

AOI22xp33_ASAP7_75t_L g2485 ( 
.A1(n_2314),
.A2(n_1980),
.B1(n_1991),
.B2(n_1890),
.Y(n_2485)
);

AOI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_2320),
.A2(n_1820),
.B1(n_1974),
.B2(n_1856),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2257),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2264),
.Y(n_2488)
);

HB1xp67_ASAP7_75t_L g2489 ( 
.A(n_2183),
.Y(n_2489)
);

INVxp33_ASAP7_75t_L g2490 ( 
.A(n_2191),
.Y(n_2490)
);

AOI22xp33_ASAP7_75t_L g2491 ( 
.A1(n_2320),
.A2(n_1986),
.B1(n_1775),
.B2(n_2111),
.Y(n_2491)
);

NAND2x1p5_ASAP7_75t_L g2492 ( 
.A(n_2199),
.B(n_1791),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2344),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2188),
.A2(n_1950),
.B1(n_1956),
.B2(n_2013),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2348),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2199),
.B(n_2188),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2132),
.Y(n_2497)
);

AO21x1_ASAP7_75t_L g2498 ( 
.A1(n_2335),
.A2(n_2140),
.B(n_2150),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2235),
.B(n_1774),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_2173),
.B(n_1965),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2306),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2157),
.B(n_2357),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2265),
.Y(n_2503)
);

INVx4_ASAP7_75t_L g2504 ( 
.A(n_2296),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2205),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2140),
.Y(n_2506)
);

NOR2x1_ASAP7_75t_SL g2507 ( 
.A(n_2199),
.B(n_1987),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_2316),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2261),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2132),
.B(n_1972),
.Y(n_2510)
);

OAI22xp5_ASAP7_75t_L g2511 ( 
.A1(n_2331),
.A2(n_2048),
.B1(n_2054),
.B2(n_1864),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2331),
.B(n_1777),
.Y(n_2512)
);

INVx4_ASAP7_75t_L g2513 ( 
.A(n_2296),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2189),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2259),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2204),
.Y(n_2516)
);

BUFx2_ASAP7_75t_SL g2517 ( 
.A(n_2197),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2438),
.Y(n_2518)
);

INVx1_ASAP7_75t_SL g2519 ( 
.A(n_2193),
.Y(n_2519)
);

HB1xp67_ASAP7_75t_L g2520 ( 
.A(n_2289),
.Y(n_2520)
);

OAI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_2177),
.A2(n_1779),
.B(n_1823),
.Y(n_2521)
);

INVx4_ASAP7_75t_L g2522 ( 
.A(n_2191),
.Y(n_2522)
);

BUFx2_ASAP7_75t_SL g2523 ( 
.A(n_2197),
.Y(n_2523)
);

CKINVDCx20_ASAP7_75t_R g2524 ( 
.A(n_2246),
.Y(n_2524)
);

BUFx3_ASAP7_75t_L g2525 ( 
.A(n_2219),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2442),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2446),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2271),
.Y(n_2528)
);

NAND2x1p5_ASAP7_75t_L g2529 ( 
.A(n_2143),
.B(n_1992),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2331),
.B(n_1929),
.Y(n_2530)
);

OAI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_2145),
.A2(n_2034),
.B1(n_2124),
.B2(n_2079),
.Y(n_2531)
);

BUFx12f_ASAP7_75t_L g2532 ( 
.A(n_2246),
.Y(n_2532)
);

AOI22xp33_ASAP7_75t_SL g2533 ( 
.A1(n_2427),
.A2(n_2445),
.B1(n_2420),
.B2(n_2148),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2272),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2273),
.Y(n_2535)
);

INVx8_ASAP7_75t_L g2536 ( 
.A(n_2185),
.Y(n_2536)
);

INVx3_ASAP7_75t_L g2537 ( 
.A(n_2204),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2274),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2275),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2277),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2288),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2244),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2245),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_2219),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2439),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2373),
.B(n_1874),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2244),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2145),
.A2(n_1983),
.B1(n_2020),
.B2(n_2062),
.Y(n_2548)
);

OR2x2_ASAP7_75t_L g2549 ( 
.A(n_2162),
.B(n_2307),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2244),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2254),
.B(n_1768),
.Y(n_2551)
);

OAI21x1_ASAP7_75t_SL g2552 ( 
.A1(n_2209),
.A2(n_1877),
.B(n_1836),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2439),
.Y(n_2553)
);

INVxp67_ASAP7_75t_L g2554 ( 
.A(n_2148),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2412),
.B(n_1874),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2171),
.Y(n_2556)
);

INVx2_ASAP7_75t_SL g2557 ( 
.A(n_2298),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2289),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2333),
.Y(n_2559)
);

BUFx2_ASAP7_75t_L g2560 ( 
.A(n_2139),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2239),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2145),
.A2(n_2042),
.B1(n_1860),
.B2(n_1902),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2333),
.Y(n_2563)
);

OR2x2_ASAP7_75t_L g2564 ( 
.A(n_2391),
.B(n_2011),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2143),
.B(n_1904),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2233),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_L g2567 ( 
.A1(n_2192),
.A2(n_2125),
.B1(n_2121),
.B2(n_2119),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2333),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2233),
.Y(n_2569)
);

INVx3_ASAP7_75t_L g2570 ( 
.A(n_2239),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2329),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2139),
.Y(n_2572)
);

OAI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2224),
.A2(n_1875),
.B(n_1835),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2329),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2240),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2240),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2241),
.Y(n_2577)
);

BUFx10_ASAP7_75t_L g2578 ( 
.A(n_2298),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2424),
.Y(n_2579)
);

INVx1_ASAP7_75t_SL g2580 ( 
.A(n_2245),
.Y(n_2580)
);

BUFx8_ASAP7_75t_L g2581 ( 
.A(n_2185),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2340),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2340),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2238),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2302),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2137),
.Y(n_2586)
);

BUFx10_ASAP7_75t_L g2587 ( 
.A(n_2298),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2246),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2447),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2384),
.B(n_2105),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2447),
.Y(n_2591)
);

OAI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2386),
.A2(n_1958),
.B1(n_1938),
.B2(n_1939),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_L g2593 ( 
.A1(n_2192),
.A2(n_2102),
.B1(n_2088),
.B2(n_2083),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2232),
.Y(n_2594)
);

BUFx2_ASAP7_75t_L g2595 ( 
.A(n_2141),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2227),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2232),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2300),
.B(n_2064),
.Y(n_2598)
);

CKINVDCx20_ASAP7_75t_R g2599 ( 
.A(n_2233),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2316),
.Y(n_2600)
);

AOI21xp33_ASAP7_75t_L g2601 ( 
.A1(n_2247),
.A2(n_1909),
.B(n_1982),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2379),
.Y(n_2602)
);

INVx2_ASAP7_75t_SL g2603 ( 
.A(n_2141),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2418),
.B(n_2005),
.Y(n_2604)
);

BUFx2_ASAP7_75t_L g2605 ( 
.A(n_2153),
.Y(n_2605)
);

INVx1_ASAP7_75t_SL g2606 ( 
.A(n_2256),
.Y(n_2606)
);

BUFx4f_ASAP7_75t_SL g2607 ( 
.A(n_2227),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2232),
.Y(n_2608)
);

CKINVDCx6p67_ASAP7_75t_R g2609 ( 
.A(n_2149),
.Y(n_2609)
);

INVx8_ASAP7_75t_L g2610 ( 
.A(n_2356),
.Y(n_2610)
);

BUFx3_ASAP7_75t_L g2611 ( 
.A(n_2149),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2361),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2241),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_2285),
.Y(n_2614)
);

BUFx2_ASAP7_75t_L g2615 ( 
.A(n_2153),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2361),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2427),
.A2(n_1803),
.B1(n_1826),
.B2(n_1993),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_2236),
.Y(n_2618)
);

INVxp67_ASAP7_75t_SL g2619 ( 
.A(n_2130),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2379),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2158),
.B(n_2052),
.Y(n_2621)
);

NAND2x1p5_ASAP7_75t_L g2622 ( 
.A(n_2163),
.B(n_2005),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2426),
.B(n_2046),
.Y(n_2623)
);

OAI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2388),
.A2(n_2038),
.B(n_2036),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2158),
.B(n_524),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_2173),
.B(n_1897),
.Y(n_2626)
);

OAI21x1_ASAP7_75t_SL g2627 ( 
.A1(n_2200),
.A2(n_2027),
.B(n_1954),
.Y(n_2627)
);

BUFx3_ASAP7_75t_L g2628 ( 
.A(n_2228),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2304),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2445),
.A2(n_2027),
.B1(n_1954),
.B2(n_1778),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2134),
.A2(n_1954),
.B1(n_1778),
.B2(n_526),
.Y(n_2631)
);

OAI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2386),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2386),
.A2(n_525),
.B1(n_527),
.B2(n_528),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_2419),
.B(n_527),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2371),
.A2(n_529),
.B1(n_530),
.B2(n_533),
.Y(n_2635)
);

INVx3_ASAP7_75t_L g2636 ( 
.A(n_2163),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2371),
.Y(n_2637)
);

CKINVDCx6p67_ASAP7_75t_R g2638 ( 
.A(n_2242),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2429),
.B(n_530),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2371),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2134),
.A2(n_533),
.B1(n_534),
.B2(n_535),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2431),
.Y(n_2642)
);

AOI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2220),
.A2(n_534),
.B1(n_536),
.B2(n_537),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2338),
.B(n_540),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_2155),
.Y(n_2645)
);

OAI22xp33_ASAP7_75t_SL g2646 ( 
.A1(n_2403),
.A2(n_541),
.B1(n_542),
.B2(n_545),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2164),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2220),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2164),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2168),
.A2(n_546),
.B1(n_549),
.B2(n_2432),
.Y(n_2650)
);

BUFx8_ASAP7_75t_L g2651 ( 
.A(n_2385),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2431),
.Y(n_2652)
);

CKINVDCx20_ASAP7_75t_R g2653 ( 
.A(n_2201),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2411),
.A2(n_549),
.B1(n_2419),
.B2(n_2212),
.Y(n_2654)
);

BUFx2_ASAP7_75t_L g2655 ( 
.A(n_2155),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2212),
.B(n_2454),
.Y(n_2656)
);

BUFx3_ASAP7_75t_L g2657 ( 
.A(n_2161),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2411),
.A2(n_2435),
.B1(n_2168),
.B2(n_2454),
.Y(n_2658)
);

BUFx2_ASAP7_75t_SL g2659 ( 
.A(n_2184),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2455),
.A2(n_2214),
.B1(n_2196),
.B2(n_2436),
.Y(n_2660)
);

BUFx8_ASAP7_75t_L g2661 ( 
.A(n_2385),
.Y(n_2661)
);

OR2x6_ASAP7_75t_L g2662 ( 
.A(n_2356),
.B(n_2186),
.Y(n_2662)
);

OAI21x1_ASAP7_75t_L g2663 ( 
.A1(n_2202),
.A2(n_2203),
.B(n_2180),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2354),
.Y(n_2664)
);

BUFx3_ASAP7_75t_L g2665 ( 
.A(n_2161),
.Y(n_2665)
);

CKINVDCx6p67_ASAP7_75t_R g2666 ( 
.A(n_2249),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2355),
.B(n_2214),
.Y(n_2667)
);

BUFx2_ASAP7_75t_L g2668 ( 
.A(n_2144),
.Y(n_2668)
);

NOR2x1_ASAP7_75t_R g2669 ( 
.A(n_2324),
.B(n_2346),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2376),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2382),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2372),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_2310),
.Y(n_2673)
);

AND2x4_ASAP7_75t_L g2674 ( 
.A(n_2412),
.B(n_2256),
.Y(n_2674)
);

INVx6_ASAP7_75t_L g2675 ( 
.A(n_2399),
.Y(n_2675)
);

AOI22xp33_ASAP7_75t_SL g2676 ( 
.A1(n_2356),
.A2(n_2147),
.B1(n_2393),
.B2(n_2387),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2435),
.A2(n_2325),
.B1(n_2395),
.B2(n_2345),
.Y(n_2677)
);

BUFx10_ASAP7_75t_L g2678 ( 
.A(n_2160),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2393),
.Y(n_2679)
);

BUFx6f_ASAP7_75t_L g2680 ( 
.A(n_2316),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_2336),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2323),
.Y(n_2682)
);

NAND2x1p5_ASAP7_75t_L g2683 ( 
.A(n_2169),
.B(n_2336),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2146),
.B(n_2305),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2267),
.B(n_2276),
.Y(n_2685)
);

CKINVDCx20_ASAP7_75t_R g2686 ( 
.A(n_2248),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2267),
.B(n_2276),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2146),
.B(n_2305),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2404),
.B(n_2430),
.Y(n_2689)
);

BUFx6f_ASAP7_75t_L g2690 ( 
.A(n_2336),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2312),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2280),
.B(n_2281),
.Y(n_2692)
);

HB1xp67_ASAP7_75t_L g2693 ( 
.A(n_2322),
.Y(n_2693)
);

INVxp67_ASAP7_75t_L g2694 ( 
.A(n_2359),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2313),
.Y(n_2695)
);

AO21x2_ASAP7_75t_L g2696 ( 
.A1(n_2135),
.A2(n_2142),
.B(n_2156),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2322),
.Y(n_2697)
);

AOI22xp33_ASAP7_75t_SL g2698 ( 
.A1(n_2359),
.A2(n_2387),
.B1(n_2136),
.B2(n_2223),
.Y(n_2698)
);

AND2x4_ASAP7_75t_L g2699 ( 
.A(n_2280),
.B(n_2281),
.Y(n_2699)
);

BUFx3_ASAP7_75t_L g2700 ( 
.A(n_2310),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2334),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2395),
.Y(n_2702)
);

BUFx3_ASAP7_75t_L g2703 ( 
.A(n_2170),
.Y(n_2703)
);

AOI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2455),
.A2(n_2196),
.B1(n_2252),
.B2(n_2131),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2433),
.Y(n_2705)
);

AOI21x1_ASAP7_75t_L g2706 ( 
.A1(n_2363),
.A2(n_2181),
.B(n_2378),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2395),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_2433),
.A2(n_2452),
.B1(n_2440),
.B2(n_2421),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2409),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_SL g2710 ( 
.A(n_2249),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2262),
.Y(n_2711)
);

INVx2_ASAP7_75t_SL g2712 ( 
.A(n_2309),
.Y(n_2712)
);

HB1xp67_ASAP7_75t_L g2713 ( 
.A(n_2398),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_R g2714 ( 
.A(n_2607),
.B(n_2351),
.Y(n_2714)
);

NAND2xp33_ASAP7_75t_R g2715 ( 
.A(n_2618),
.B(n_2324),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2499),
.B(n_2430),
.Y(n_2716)
);

OR2x6_ASAP7_75t_L g2717 ( 
.A(n_2536),
.B(n_2319),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2644),
.B(n_2217),
.Y(n_2718)
);

AOI22xp33_ASAP7_75t_SL g2719 ( 
.A1(n_2684),
.A2(n_2387),
.B1(n_2359),
.B2(n_2130),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_SL g2720 ( 
.A1(n_2688),
.A2(n_2387),
.B1(n_2359),
.B2(n_2130),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_R g2721 ( 
.A(n_2607),
.B(n_2351),
.Y(n_2721)
);

CKINVDCx16_ASAP7_75t_R g2722 ( 
.A(n_2532),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2460),
.Y(n_2723)
);

HB1xp67_ASAP7_75t_L g2724 ( 
.A(n_2497),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2705),
.B(n_2398),
.Y(n_2725)
);

INVx3_ASAP7_75t_L g2726 ( 
.A(n_2472),
.Y(n_2726)
);

AO32x2_ASAP7_75t_L g2727 ( 
.A1(n_2635),
.A2(n_2389),
.A3(n_2366),
.B1(n_2341),
.B2(n_2328),
.Y(n_2727)
);

OAI222xp33_ASAP7_75t_L g2728 ( 
.A1(n_2660),
.A2(n_2262),
.B1(n_2263),
.B2(n_2335),
.C1(n_2186),
.C2(n_2434),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2497),
.B(n_2318),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2581),
.Y(n_2730)
);

OAI21xp33_ASAP7_75t_SL g2731 ( 
.A1(n_2660),
.A2(n_2434),
.B(n_2353),
.Y(n_2731)
);

OAI222xp33_ASAP7_75t_L g2732 ( 
.A1(n_2533),
.A2(n_2263),
.B1(n_2401),
.B2(n_2406),
.C1(n_2292),
.C2(n_2383),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_SL g2733 ( 
.A1(n_2463),
.A2(n_2292),
.B(n_2397),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2461),
.A2(n_2359),
.B1(n_2387),
.B2(n_2270),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2694),
.B(n_2178),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2545),
.B(n_2190),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_SL g2737 ( 
.A1(n_2599),
.A2(n_2346),
.B1(n_2400),
.B2(n_2248),
.Y(n_2737)
);

BUFx6f_ASAP7_75t_L g2738 ( 
.A(n_2472),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2536),
.Y(n_2739)
);

OR2x6_ASAP7_75t_L g2740 ( 
.A(n_2536),
.B(n_2287),
.Y(n_2740)
);

BUFx2_ASAP7_75t_L g2741 ( 
.A(n_2478),
.Y(n_2741)
);

O2A1O1Ixp33_ASAP7_75t_L g2742 ( 
.A1(n_2635),
.A2(n_2422),
.B(n_2457),
.C(n_2299),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2464),
.B(n_2301),
.Y(n_2743)
);

NAND2xp33_ASAP7_75t_R g2744 ( 
.A(n_2588),
.B(n_2400),
.Y(n_2744)
);

BUFx2_ASAP7_75t_L g2745 ( 
.A(n_2478),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_2713),
.Y(n_2746)
);

INVx1_ASAP7_75t_SL g2747 ( 
.A(n_2638),
.Y(n_2747)
);

OAI21xp33_ASAP7_75t_L g2748 ( 
.A1(n_2533),
.A2(n_2350),
.B(n_2397),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2465),
.Y(n_2749)
);

OR2x6_ASAP7_75t_L g2750 ( 
.A(n_2610),
.B(n_2278),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2466),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2469),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2713),
.Y(n_2753)
);

OAI21x1_ASAP7_75t_L g2754 ( 
.A1(n_2663),
.A2(n_2303),
.B(n_2218),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2694),
.B(n_2178),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2553),
.B(n_2519),
.Y(n_2756)
);

BUFx2_ASAP7_75t_L g2757 ( 
.A(n_2503),
.Y(n_2757)
);

BUFx12f_ASAP7_75t_L g2758 ( 
.A(n_2581),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2611),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2519),
.B(n_2549),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2474),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2476),
.B(n_2269),
.Y(n_2762)
);

NAND2xp33_ASAP7_75t_R g2763 ( 
.A(n_2709),
.B(n_2405),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2479),
.B(n_2279),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_R g2765 ( 
.A(n_2524),
.B(n_2278),
.Y(n_2765)
);

OR2x6_ASAP7_75t_L g2766 ( 
.A(n_2610),
.B(n_2399),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_R g2767 ( 
.A(n_2596),
.B(n_2405),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2609),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2651),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2480),
.B(n_2208),
.Y(n_2770)
);

INVx2_ASAP7_75t_SL g2771 ( 
.A(n_2566),
.Y(n_2771)
);

NOR3xp33_ASAP7_75t_SL g2772 ( 
.A(n_2656),
.B(n_2215),
.C(n_2377),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2467),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2481),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2667),
.B(n_2367),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2483),
.B(n_2211),
.Y(n_2776)
);

NAND2xp33_ASAP7_75t_SL g2777 ( 
.A(n_2506),
.B(n_2154),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2461),
.A2(n_2293),
.B1(n_2258),
.B2(n_2428),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2534),
.B(n_2315),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2487),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2488),
.B(n_2211),
.Y(n_2781)
);

AOI22xp33_ASAP7_75t_L g2782 ( 
.A1(n_2511),
.A2(n_2380),
.B1(n_2182),
.B2(n_2443),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2689),
.B(n_2315),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2493),
.B(n_2216),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2495),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2501),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2629),
.B(n_2321),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2555),
.B(n_2187),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2625),
.B(n_2321),
.Y(n_2789)
);

AOI22xp33_ASAP7_75t_L g2790 ( 
.A1(n_2511),
.A2(n_2448),
.B1(n_2231),
.B2(n_2417),
.Y(n_2790)
);

NAND3xp33_ASAP7_75t_SL g2791 ( 
.A(n_2463),
.B(n_2349),
.C(n_2234),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2459),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2586),
.B(n_2326),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2585),
.B(n_2326),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2531),
.A2(n_2448),
.B1(n_2417),
.B2(n_2449),
.Y(n_2795)
);

BUFx2_ASAP7_75t_L g2796 ( 
.A(n_2503),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2514),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2515),
.B(n_2229),
.Y(n_2798)
);

OR2x6_ASAP7_75t_L g2799 ( 
.A(n_2610),
.B(n_2195),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2541),
.B(n_2294),
.Y(n_2800)
);

CKINVDCx20_ASAP7_75t_R g2801 ( 
.A(n_2651),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_R g2802 ( 
.A(n_2653),
.B(n_2686),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2462),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2472),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2569),
.Y(n_2805)
);

CKINVDCx20_ASAP7_75t_R g2806 ( 
.A(n_2661),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2467),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2518),
.Y(n_2808)
);

NAND2xp33_ASAP7_75t_R g2809 ( 
.A(n_2709),
.B(n_2154),
.Y(n_2809)
);

CKINVDCx11_ASAP7_75t_R g2810 ( 
.A(n_2504),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2526),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2531),
.A2(n_2449),
.B1(n_2437),
.B2(n_2317),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_R g2813 ( 
.A(n_2470),
.B(n_2130),
.Y(n_2813)
);

A2O1A1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2704),
.A2(n_2210),
.B(n_2215),
.C(n_2456),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2527),
.B(n_2229),
.Y(n_2815)
);

CKINVDCx8_ASAP7_75t_R g2816 ( 
.A(n_2517),
.Y(n_2816)
);

INVx1_ASAP7_75t_SL g2817 ( 
.A(n_2523),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2704),
.A2(n_2406),
.B1(n_2401),
.B2(n_2390),
.Y(n_2818)
);

CKINVDCx16_ASAP7_75t_R g2819 ( 
.A(n_2470),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2650),
.A2(n_2453),
.B1(n_2260),
.B2(n_2268),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2505),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2509),
.Y(n_2822)
);

NAND3xp33_ASAP7_75t_SL g2823 ( 
.A(n_2632),
.B(n_2255),
.C(n_2159),
.Y(n_2823)
);

BUFx4f_ASAP7_75t_SL g2824 ( 
.A(n_2661),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2504),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2560),
.B(n_2187),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2548),
.A2(n_2416),
.B1(n_2415),
.B2(n_2413),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_2484),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2621),
.A2(n_2416),
.B1(n_2415),
.B2(n_2413),
.Y(n_2829)
);

OAI222xp33_ASAP7_75t_L g2830 ( 
.A1(n_2662),
.A2(n_2347),
.B1(n_2194),
.B2(n_2174),
.C1(n_2308),
.C2(n_2221),
.Y(n_2830)
);

NOR2x1_ASAP7_75t_L g2831 ( 
.A(n_2636),
.B(n_2423),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_R g2832 ( 
.A(n_2475),
.B(n_2130),
.Y(n_2832)
);

CKINVDCx20_ASAP7_75t_R g2833 ( 
.A(n_2525),
.Y(n_2833)
);

AOI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2548),
.A2(n_2311),
.B1(n_2297),
.B2(n_2410),
.Y(n_2834)
);

OR2x6_ASAP7_75t_L g2835 ( 
.A(n_2475),
.B(n_2309),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2578),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_SL g2837 ( 
.A(n_2632),
.B(n_2633),
.C(n_2658),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2528),
.B(n_2230),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2555),
.B(n_2226),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2678),
.Y(n_2840)
);

HB1xp67_ASAP7_75t_L g2841 ( 
.A(n_2468),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2471),
.A2(n_2450),
.B(n_2456),
.Y(n_2842)
);

AO21x2_ASAP7_75t_L g2843 ( 
.A1(n_2627),
.A2(n_2207),
.B(n_2142),
.Y(n_2843)
);

OAI222xp33_ASAP7_75t_L g2844 ( 
.A1(n_2662),
.A2(n_2251),
.B1(n_2294),
.B2(n_2330),
.C1(n_2332),
.C2(n_2352),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2572),
.B(n_2226),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2595),
.B(n_2330),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2605),
.B(n_2332),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2615),
.B(n_2358),
.Y(n_2848)
);

NAND3xp33_ASAP7_75t_SL g2849 ( 
.A(n_2633),
.B(n_2284),
.C(n_2237),
.Y(n_2849)
);

AND2x4_ASAP7_75t_L g2850 ( 
.A(n_2674),
.B(n_2336),
.Y(n_2850)
);

NAND2xp33_ASAP7_75t_R g2851 ( 
.A(n_2662),
.B(n_2181),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2535),
.Y(n_2852)
);

O2A1O1Ixp33_ASAP7_75t_SL g2853 ( 
.A1(n_2589),
.A2(n_2407),
.B(n_2136),
.C(n_2130),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2513),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2538),
.Y(n_2855)
);

NAND2xp33_ASAP7_75t_R g2856 ( 
.A(n_2636),
.B(n_2181),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2539),
.B(n_2230),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2540),
.Y(n_2858)
);

CKINVDCx16_ASAP7_75t_R g2859 ( 
.A(n_2513),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2691),
.Y(n_2860)
);

BUFx10_ASAP7_75t_L g2861 ( 
.A(n_2675),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2695),
.Y(n_2862)
);

CKINVDCx16_ASAP7_75t_R g2863 ( 
.A(n_2522),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_2710),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2701),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2502),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2502),
.Y(n_2867)
);

NOR2xp33_ASAP7_75t_R g2868 ( 
.A(n_2675),
.B(n_2136),
.Y(n_2868)
);

OAI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2650),
.A2(n_2260),
.B1(n_2268),
.B2(n_2425),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2655),
.B(n_2358),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2657),
.B(n_2358),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2665),
.B(n_2358),
.Y(n_2872)
);

CKINVDCx16_ASAP7_75t_R g2873 ( 
.A(n_2522),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2551),
.B(n_2392),
.Y(n_2874)
);

AND2x4_ASAP7_75t_L g2875 ( 
.A(n_2674),
.B(n_2408),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2556),
.B(n_2500),
.Y(n_2876)
);

NAND2xp33_ASAP7_75t_R g2877 ( 
.A(n_2647),
.B(n_2260),
.Y(n_2877)
);

NAND3xp33_ASAP7_75t_SL g2878 ( 
.A(n_2677),
.B(n_2291),
.C(n_2352),
.Y(n_2878)
);

BUFx3_ASAP7_75t_L g2879 ( 
.A(n_2544),
.Y(n_2879)
);

NAND2xp33_ASAP7_75t_R g2880 ( 
.A(n_2647),
.B(n_2268),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2639),
.Y(n_2881)
);

OR2x6_ASAP7_75t_L g2882 ( 
.A(n_2659),
.B(n_2309),
.Y(n_2882)
);

OR2x6_ASAP7_75t_L g2883 ( 
.A(n_2683),
.B(n_2402),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2710),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2637),
.B(n_2364),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2590),
.B(n_2392),
.Y(n_2886)
);

NOR3xp33_ASAP7_75t_SL g2887 ( 
.A(n_2640),
.B(n_2592),
.C(n_2634),
.Y(n_2887)
);

INVx4_ASAP7_75t_L g2888 ( 
.A(n_2508),
.Y(n_2888)
);

OAI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2471),
.A2(n_2425),
.B1(n_2392),
.B2(n_2394),
.Y(n_2889)
);

NAND2xp33_ASAP7_75t_R g2890 ( 
.A(n_2649),
.B(n_2702),
.Y(n_2890)
);

CKINVDCx5p33_ASAP7_75t_R g2891 ( 
.A(n_2666),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2673),
.B(n_2364),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_2614),
.Y(n_2893)
);

A2O1A1Ixp33_ASAP7_75t_L g2894 ( 
.A1(n_2676),
.A2(n_2266),
.B(n_2444),
.C(n_2441),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2639),
.Y(n_2895)
);

NAND3xp33_ASAP7_75t_SL g2896 ( 
.A(n_2591),
.B(n_2458),
.C(n_2360),
.Y(n_2896)
);

CKINVDCx5p33_ASAP7_75t_R g2897 ( 
.A(n_2578),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2587),
.Y(n_2898)
);

AOI221xp5_ASAP7_75t_L g2899 ( 
.A1(n_2654),
.A2(n_2282),
.B1(n_2176),
.B2(n_2207),
.C(n_2172),
.Y(n_2899)
);

CKINVDCx20_ASAP7_75t_R g2900 ( 
.A(n_2587),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2700),
.B(n_2364),
.Y(n_2901)
);

INVxp67_ASAP7_75t_SL g2902 ( 
.A(n_2468),
.Y(n_2902)
);

AO31x2_ASAP7_75t_L g2903 ( 
.A1(n_2498),
.A2(n_2374),
.A3(n_2343),
.B(n_2368),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_R g2904 ( 
.A(n_2516),
.B(n_2136),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2642),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2598),
.B(n_2337),
.Y(n_2906)
);

OR2x2_ASAP7_75t_L g2907 ( 
.A(n_2520),
.B(n_2458),
.Y(n_2907)
);

AOI22xp33_ASAP7_75t_L g2908 ( 
.A1(n_2491),
.A2(n_2136),
.B1(n_2223),
.B2(n_2243),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2652),
.Y(n_2909)
);

INVxp67_ASAP7_75t_SL g2910 ( 
.A(n_2506),
.Y(n_2910)
);

INVx4_ASAP7_75t_L g2911 ( 
.A(n_2508),
.Y(n_2911)
);

NAND2xp33_ASAP7_75t_R g2912 ( 
.A(n_2649),
.B(n_2250),
.Y(n_2912)
);

BUFx2_ASAP7_75t_L g2913 ( 
.A(n_2561),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_2558),
.B(n_2362),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2604),
.Y(n_2915)
);

OAI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2708),
.A2(n_2295),
.B(n_2286),
.Y(n_2916)
);

OR2x2_ASAP7_75t_L g2917 ( 
.A(n_2558),
.B(n_2368),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2604),
.Y(n_2918)
);

CKINVDCx8_ASAP7_75t_R g2919 ( 
.A(n_2668),
.Y(n_2919)
);

AND4x1_ASAP7_75t_L g2920 ( 
.A(n_2643),
.B(n_2409),
.C(n_2136),
.D(n_2223),
.Y(n_2920)
);

AND2x4_ASAP7_75t_SL g2921 ( 
.A(n_2678),
.B(n_2360),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2682),
.B(n_2623),
.Y(n_2922)
);

CKINVDCx5p33_ASAP7_75t_R g2923 ( 
.A(n_2628),
.Y(n_2923)
);

INVx3_ASAP7_75t_L g2924 ( 
.A(n_2600),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2603),
.B(n_2339),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2623),
.B(n_2414),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_2703),
.Y(n_2927)
);

OR2x6_ASAP7_75t_L g2928 ( 
.A(n_2683),
.B(n_2402),
.Y(n_2928)
);

CKINVDCx5p33_ASAP7_75t_R g2929 ( 
.A(n_2557),
.Y(n_2929)
);

NOR3xp33_ASAP7_75t_SL g2930 ( 
.A(n_2592),
.B(n_2223),
.C(n_2156),
.Y(n_2930)
);

HB1xp67_ASAP7_75t_L g2931 ( 
.A(n_2482),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2645),
.B(n_2286),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2582),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_2707),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2564),
.B(n_2561),
.Y(n_2935)
);

NAND3xp33_ASAP7_75t_SL g2936 ( 
.A(n_2490),
.B(n_2365),
.C(n_2369),
.Y(n_2936)
);

NAND2x1_ASAP7_75t_L g2937 ( 
.A(n_2496),
.B(n_2365),
.Y(n_2937)
);

BUFx3_ASAP7_75t_L g2938 ( 
.A(n_2712),
.Y(n_2938)
);

INVx4_ASAP7_75t_L g2939 ( 
.A(n_2600),
.Y(n_2939)
);

OR2x2_ASAP7_75t_L g2940 ( 
.A(n_2679),
.B(n_2396),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2679),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2489),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_2537),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2510),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2491),
.A2(n_2223),
.B1(n_2243),
.B2(n_2451),
.Y(n_2945)
);

NAND2xp33_ASAP7_75t_R g2946 ( 
.A(n_2537),
.B(n_2250),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2562),
.A2(n_2342),
.B1(n_2408),
.B2(n_2381),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_R g2948 ( 
.A(n_2570),
.B(n_2408),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2554),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2693),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2792),
.Y(n_2951)
);

NAND2xp33_ASAP7_75t_R g2952 ( 
.A(n_2948),
.B(n_2496),
.Y(n_2952)
);

HB1xp67_ASAP7_75t_L g2953 ( 
.A(n_2773),
.Y(n_2953)
);

INVx5_ASAP7_75t_L g2954 ( 
.A(n_2717),
.Y(n_2954)
);

INVx3_ASAP7_75t_L g2955 ( 
.A(n_2741),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2935),
.B(n_2582),
.Y(n_2956)
);

BUFx3_ASAP7_75t_L g2957 ( 
.A(n_2921),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2874),
.B(n_2583),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_2791),
.A2(n_2552),
.B1(n_2573),
.B2(n_2617),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2723),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2866),
.B(n_2546),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2775),
.B(n_2583),
.Y(n_2962)
);

OAI31xp33_ASAP7_75t_SL g2963 ( 
.A1(n_2837),
.A2(n_2676),
.A3(n_2698),
.B(n_2711),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2749),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2716),
.B(n_2602),
.Y(n_2965)
);

OA21x2_ASAP7_75t_L g2966 ( 
.A1(n_2754),
.A2(n_2842),
.B(n_2916),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2751),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2729),
.B(n_2602),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2752),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2783),
.B(n_2620),
.Y(n_2970)
);

HB1xp67_ASAP7_75t_L g2971 ( 
.A(n_2807),
.Y(n_2971)
);

INVxp67_ASAP7_75t_L g2972 ( 
.A(n_2841),
.Y(n_2972)
);

OR2x2_ASAP7_75t_L g2973 ( 
.A(n_2756),
.B(n_2760),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2944),
.B(n_2620),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2867),
.B(n_2546),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2718),
.B(n_2693),
.Y(n_2976)
);

AOI22xp33_ASAP7_75t_L g2977 ( 
.A1(n_2849),
.A2(n_2573),
.B1(n_2617),
.B2(n_2512),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2793),
.B(n_2697),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2803),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2902),
.B(n_2697),
.Y(n_2980)
);

BUFx2_ASAP7_75t_L g2981 ( 
.A(n_2717),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2886),
.B(n_2554),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2761),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2789),
.B(n_2542),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2736),
.B(n_2547),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2787),
.B(n_2550),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2724),
.B(n_2543),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2794),
.B(n_2543),
.Y(n_2988)
);

AND2x4_ASAP7_75t_L g2989 ( 
.A(n_2910),
.B(n_2619),
.Y(n_2989)
);

OAI221xp5_ASAP7_75t_L g2990 ( 
.A1(n_2733),
.A2(n_2486),
.B1(n_2562),
.B2(n_2485),
.C(n_2648),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2906),
.B(n_2580),
.Y(n_2991)
);

AOI22xp33_ASAP7_75t_SL g2992 ( 
.A1(n_2731),
.A2(n_2646),
.B1(n_2574),
.B2(n_2571),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2774),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2780),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2745),
.B(n_2580),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2942),
.B(n_2670),
.Y(n_2996)
);

INVxp67_ASAP7_75t_L g2997 ( 
.A(n_2931),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2785),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2786),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2748),
.B(n_2530),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_2757),
.B(n_2606),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2797),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2746),
.B(n_2606),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2796),
.B(n_2612),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2834),
.A2(n_2601),
.B(n_2671),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2808),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2788),
.B(n_2619),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2848),
.B(n_2616),
.Y(n_3008)
);

AND2x2_ASAP7_75t_SL g3009 ( 
.A(n_2920),
.B(n_2698),
.Y(n_3009)
);

INVxp67_ASAP7_75t_L g3010 ( 
.A(n_2753),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2915),
.B(n_2630),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2811),
.Y(n_3012)
);

BUFx2_ASAP7_75t_L g3013 ( 
.A(n_2888),
.Y(n_3013)
);

BUFx2_ASAP7_75t_L g3014 ( 
.A(n_2888),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2918),
.B(n_2630),
.Y(n_3015)
);

INVxp67_ASAP7_75t_L g3016 ( 
.A(n_2950),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2821),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2941),
.B(n_2559),
.Y(n_3018)
);

HB1xp67_ASAP7_75t_L g3019 ( 
.A(n_2933),
.Y(n_3019)
);

BUFx3_ASAP7_75t_L g3020 ( 
.A(n_2816),
.Y(n_3020)
);

AND2x4_ASAP7_75t_L g3021 ( 
.A(n_2788),
.B(n_2570),
.Y(n_3021)
);

INVx3_ASAP7_75t_L g3022 ( 
.A(n_2911),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2823),
.B(n_2584),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2870),
.B(n_2905),
.Y(n_3024)
);

OAI21x1_ASAP7_75t_SL g3025 ( 
.A1(n_2831),
.A2(n_2507),
.B(n_2706),
.Y(n_3025)
);

BUFx3_ASAP7_75t_L g3026 ( 
.A(n_2850),
.Y(n_3026)
);

AND2x2_ASAP7_75t_L g3027 ( 
.A(n_2909),
.B(n_2846),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2881),
.B(n_2563),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2822),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2847),
.B(n_2575),
.Y(n_3030)
);

OR2x2_ASAP7_75t_L g3031 ( 
.A(n_2725),
.B(n_2575),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2852),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2855),
.Y(n_3033)
);

HB1xp67_ASAP7_75t_L g3034 ( 
.A(n_2914),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2858),
.B(n_2826),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2860),
.Y(n_3036)
);

INVx3_ASAP7_75t_L g3037 ( 
.A(n_2911),
.Y(n_3037)
);

HB1xp67_ASAP7_75t_L g3038 ( 
.A(n_2917),
.Y(n_3038)
);

HB1xp67_ASAP7_75t_L g3039 ( 
.A(n_2940),
.Y(n_3039)
);

OR2x2_ASAP7_75t_L g3040 ( 
.A(n_2876),
.B(n_2576),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2862),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2865),
.Y(n_3042)
);

INVx5_ASAP7_75t_SL g3043 ( 
.A(n_2766),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2845),
.B(n_2871),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2895),
.B(n_2568),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2949),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2800),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2779),
.Y(n_3048)
);

OR2x2_ASAP7_75t_L g3049 ( 
.A(n_2922),
.B(n_2907),
.Y(n_3049)
);

INVx3_ASAP7_75t_L g3050 ( 
.A(n_2939),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2762),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2872),
.B(n_2576),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2926),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2764),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2743),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2913),
.B(n_2850),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_2875),
.B(n_2577),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2875),
.B(n_2577),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2892),
.B(n_2613),
.Y(n_3059)
);

AND2x4_ASAP7_75t_L g3060 ( 
.A(n_2839),
.B(n_2613),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2901),
.B(n_2594),
.Y(n_3061)
);

INVx4_ASAP7_75t_L g3062 ( 
.A(n_2766),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_2885),
.B(n_2597),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2838),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2817),
.B(n_2579),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2879),
.B(n_2608),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2857),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2770),
.Y(n_3068)
);

INVx2_ASAP7_75t_SL g3069 ( 
.A(n_2739),
.Y(n_3069)
);

BUFx2_ASAP7_75t_L g3070 ( 
.A(n_2939),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2776),
.Y(n_3071)
);

AND2x4_ASAP7_75t_L g3072 ( 
.A(n_2839),
.B(n_2685),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2781),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2784),
.B(n_2626),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2727),
.B(n_2685),
.Y(n_3075)
);

OR2x2_ASAP7_75t_L g3076 ( 
.A(n_2798),
.B(n_2687),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_2727),
.B(n_2687),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2727),
.B(n_2692),
.Y(n_3078)
);

AND2x2_ASAP7_75t_L g3079 ( 
.A(n_2938),
.B(n_2692),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2759),
.B(n_2699),
.Y(n_3080)
);

BUFx3_ASAP7_75t_L g3081 ( 
.A(n_2882),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2815),
.B(n_2696),
.Y(n_3082)
);

INVx3_ASAP7_75t_L g3083 ( 
.A(n_2937),
.Y(n_3083)
);

INVx4_ASAP7_75t_L g3084 ( 
.A(n_2740),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2840),
.B(n_2699),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2919),
.B(n_2600),
.Y(n_3086)
);

OR2x2_ASAP7_75t_L g3087 ( 
.A(n_2882),
.B(n_2622),
.Y(n_3087)
);

INVx5_ASAP7_75t_SL g3088 ( 
.A(n_2750),
.Y(n_3088)
);

OAI22xp5_ASAP7_75t_L g3089 ( 
.A1(n_2812),
.A2(n_2473),
.B1(n_2643),
.B2(n_2648),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2843),
.Y(n_3090)
);

BUFx3_ASAP7_75t_L g3091 ( 
.A(n_2738),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2925),
.B(n_2680),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2960),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2964),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2951),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2991),
.B(n_2903),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2967),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_3051),
.B(n_2829),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3044),
.B(n_2968),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2976),
.B(n_2932),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2951),
.Y(n_3101)
);

OR2x2_ASAP7_75t_L g3102 ( 
.A(n_2973),
.B(n_2863),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2969),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2983),
.Y(n_3104)
);

BUFx2_ASAP7_75t_L g3105 ( 
.A(n_3013),
.Y(n_3105)
);

INVx2_ASAP7_75t_SL g3106 ( 
.A(n_3083),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2979),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_3064),
.B(n_3067),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2993),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2994),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2979),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_3068),
.B(n_2903),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_3071),
.B(n_2903),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2998),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_R g3115 ( 
.A(n_2952),
.B(n_2859),
.Y(n_3115)
);

OR2x2_ASAP7_75t_L g3116 ( 
.A(n_3034),
.B(n_2873),
.Y(n_3116)
);

AND2x2_ASAP7_75t_SL g3117 ( 
.A(n_3009),
.B(n_2819),
.Y(n_3117)
);

INVx5_ASAP7_75t_SL g3118 ( 
.A(n_3009),
.Y(n_3118)
);

AND2x4_ASAP7_75t_SL g3119 ( 
.A(n_3062),
.B(n_2740),
.Y(n_3119)
);

HB1xp67_ASAP7_75t_L g3120 ( 
.A(n_2953),
.Y(n_3120)
);

OR2x2_ASAP7_75t_L g3121 ( 
.A(n_3034),
.B(n_3038),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3073),
.B(n_2664),
.Y(n_3122)
);

OR2x2_ASAP7_75t_L g3123 ( 
.A(n_3038),
.B(n_2771),
.Y(n_3123)
);

AND2x4_ASAP7_75t_SL g3124 ( 
.A(n_3062),
.B(n_2750),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_3024),
.B(n_2672),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_3054),
.B(n_2795),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2999),
.Y(n_3127)
);

NOR3xp33_ASAP7_75t_L g3128 ( 
.A(n_2990),
.B(n_2728),
.C(n_2818),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_3055),
.B(n_2827),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3002),
.Y(n_3130)
);

INVx1_ASAP7_75t_SL g3131 ( 
.A(n_2957),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3006),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2956),
.B(n_2719),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3012),
.Y(n_3134)
);

AOI221xp5_ASAP7_75t_L g3135 ( 
.A1(n_2990),
.A2(n_2742),
.B1(n_2814),
.B2(n_2772),
.C(n_2820),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3017),
.Y(n_3136)
);

OR2x2_ASAP7_75t_L g3137 ( 
.A(n_3039),
.B(n_2805),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_3039),
.B(n_2887),
.Y(n_3138)
);

AND2x4_ASAP7_75t_L g3139 ( 
.A(n_3075),
.B(n_2930),
.Y(n_3139)
);

INVx2_ASAP7_75t_SL g3140 ( 
.A(n_3083),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3032),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3033),
.Y(n_3142)
);

OAI21xp33_ASAP7_75t_L g3143 ( 
.A1(n_2963),
.A2(n_2778),
.B(n_2790),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_2987),
.B(n_2720),
.Y(n_3144)
);

OR2x2_ASAP7_75t_L g3145 ( 
.A(n_3049),
.B(n_2828),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_3035),
.B(n_2735),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2978),
.B(n_2735),
.Y(n_3147)
);

BUFx2_ASAP7_75t_L g3148 ( 
.A(n_3014),
.Y(n_3148)
);

HB1xp67_ASAP7_75t_L g3149 ( 
.A(n_2953),
.Y(n_3149)
);

HB1xp67_ASAP7_75t_L g3150 ( 
.A(n_2971),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_3053),
.B(n_2782),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3036),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3041),
.Y(n_3153)
);

NOR2x1_ASAP7_75t_L g3154 ( 
.A(n_3084),
.B(n_2801),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_3077),
.B(n_2755),
.Y(n_3155)
);

INVx2_ASAP7_75t_SL g3156 ( 
.A(n_3026),
.Y(n_3156)
);

OR2x2_ASAP7_75t_L g3157 ( 
.A(n_2971),
.B(n_2836),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_3042),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2962),
.B(n_2755),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3029),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3019),
.Y(n_3161)
);

AND2x4_ASAP7_75t_L g3162 ( 
.A(n_3078),
.B(n_2738),
.Y(n_3162)
);

INVx3_ASAP7_75t_L g3163 ( 
.A(n_3119),
.Y(n_3163)
);

OR2x2_ASAP7_75t_L g3164 ( 
.A(n_3121),
.B(n_2972),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_3120),
.Y(n_3165)
);

OR2x2_ASAP7_75t_L g3166 ( 
.A(n_3120),
.B(n_2972),
.Y(n_3166)
);

AND2x4_ASAP7_75t_L g3167 ( 
.A(n_3106),
.B(n_3140),
.Y(n_3167)
);

HB1xp67_ASAP7_75t_L g3168 ( 
.A(n_3149),
.Y(n_3168)
);

NOR3xp33_ASAP7_75t_SL g3169 ( 
.A(n_3143),
.B(n_2722),
.C(n_2952),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_3099),
.B(n_3092),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3100),
.B(n_3056),
.Y(n_3171)
);

BUFx2_ASAP7_75t_L g3172 ( 
.A(n_3115),
.Y(n_3172)
);

OR2x2_ASAP7_75t_L g3173 ( 
.A(n_3149),
.B(n_2997),
.Y(n_3173)
);

OR2x2_ASAP7_75t_L g3174 ( 
.A(n_3150),
.B(n_2997),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_3108),
.B(n_3046),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3095),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_3155),
.B(n_3146),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3155),
.B(n_3027),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3155),
.B(n_3019),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_3138),
.B(n_3023),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_3108),
.B(n_3010),
.Y(n_3181)
);

AOI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_3128),
.A2(n_2959),
.B1(n_2977),
.B2(n_3023),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3150),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_3112),
.B(n_3010),
.Y(n_3184)
);

NOR2xp67_ASAP7_75t_L g3185 ( 
.A(n_3116),
.B(n_3084),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_3147),
.B(n_2970),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_SL g3187 ( 
.A(n_3115),
.B(n_2963),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_3159),
.B(n_2965),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3093),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_3112),
.B(n_3082),
.Y(n_3190)
);

OR2x2_ASAP7_75t_L g3191 ( 
.A(n_3161),
.B(n_3016),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_3105),
.B(n_2988),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3113),
.B(n_3082),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_3148),
.B(n_3030),
.Y(n_3194)
);

AND2x4_ASAP7_75t_L g3195 ( 
.A(n_3106),
.B(n_2980),
.Y(n_3195)
);

NOR2xp67_ASAP7_75t_SL g3196 ( 
.A(n_3156),
.B(n_2758),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3094),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3097),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_3140),
.B(n_3156),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_3095),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3113),
.B(n_3011),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3103),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3160),
.B(n_3011),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3104),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3109),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_3101),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3098),
.B(n_3015),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3110),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3114),
.B(n_3015),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3127),
.Y(n_3210)
);

OAI21xp33_ASAP7_75t_L g3211 ( 
.A1(n_3128),
.A2(n_2959),
.B(n_2992),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3101),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3144),
.B(n_3133),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_3130),
.B(n_3074),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_3162),
.B(n_3052),
.Y(n_3215)
);

NOR2x1_ASAP7_75t_L g3216 ( 
.A(n_3154),
.B(n_2957),
.Y(n_3216)
);

NOR2x1_ASAP7_75t_SL g3217 ( 
.A(n_3102),
.B(n_2954),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3123),
.B(n_3016),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3162),
.B(n_2958),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3162),
.B(n_3048),
.Y(n_3220)
);

OR2x2_ASAP7_75t_L g3221 ( 
.A(n_3137),
.B(n_2980),
.Y(n_3221)
);

NOR4xp25_ASAP7_75t_SL g3222 ( 
.A(n_3135),
.B(n_2981),
.C(n_2890),
.D(n_2851),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_3125),
.B(n_2995),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_3125),
.B(n_3001),
.Y(n_3224)
);

AOI31xp33_ASAP7_75t_L g3225 ( 
.A1(n_3131),
.A2(n_2992),
.A3(n_2747),
.B(n_3086),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3132),
.Y(n_3226)
);

OR2x2_ASAP7_75t_L g3227 ( 
.A(n_3190),
.B(n_3129),
.Y(n_3227)
);

A2O1A1Ixp33_ASAP7_75t_L g3228 ( 
.A1(n_3216),
.A2(n_3124),
.B(n_3119),
.C(n_3117),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3207),
.B(n_3096),
.Y(n_3229)
);

AND2x2_ASAP7_75t_L g3230 ( 
.A(n_3179),
.B(n_3096),
.Y(n_3230)
);

OR2x2_ASAP7_75t_L g3231 ( 
.A(n_3190),
.B(n_3126),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3166),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3207),
.B(n_3151),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3173),
.Y(n_3234)
);

HB1xp67_ASAP7_75t_L g3235 ( 
.A(n_3168),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_3177),
.B(n_3139),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3215),
.B(n_3139),
.Y(n_3237)
);

OAI33xp33_ASAP7_75t_L g3238 ( 
.A1(n_3187),
.A2(n_3145),
.A3(n_3157),
.B1(n_3089),
.B2(n_3074),
.B3(n_3142),
.Y(n_3238)
);

AOI22xp5_ASAP7_75t_L g3239 ( 
.A1(n_3211),
.A2(n_3187),
.B1(n_3117),
.B2(n_3182),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3174),
.Y(n_3240)
);

NOR2x1p5_ASAP7_75t_SL g3241 ( 
.A(n_3169),
.B(n_3090),
.Y(n_3241)
);

INVx1_ASAP7_75t_SL g3242 ( 
.A(n_3172),
.Y(n_3242)
);

NAND4xp75_ASAP7_75t_L g3243 ( 
.A(n_3169),
.B(n_3000),
.C(n_3069),
.D(n_3080),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3184),
.Y(n_3244)
);

XOR2x2_ASAP7_75t_L g3245 ( 
.A(n_3185),
.B(n_2824),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3201),
.B(n_3134),
.Y(n_3246)
);

OR2x2_ASAP7_75t_L g3247 ( 
.A(n_3193),
.B(n_3107),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3201),
.B(n_3136),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3184),
.Y(n_3249)
);

O2A1O1Ixp33_ASAP7_75t_L g3250 ( 
.A1(n_3225),
.A2(n_2977),
.B(n_3089),
.C(n_3020),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_3163),
.B(n_2810),
.Y(n_3251)
);

INVx2_ASAP7_75t_SL g3252 ( 
.A(n_3163),
.Y(n_3252)
);

INVx3_ASAP7_75t_L g3253 ( 
.A(n_3167),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3203),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3203),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3165),
.Y(n_3256)
);

HB1xp67_ASAP7_75t_L g3257 ( 
.A(n_3168),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3183),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3189),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3197),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3198),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3202),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3209),
.B(n_3141),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_3178),
.B(n_3139),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3204),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3209),
.B(n_3152),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3205),
.Y(n_3267)
);

INVx6_ASAP7_75t_L g3268 ( 
.A(n_3199),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_3180),
.B(n_3124),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_3199),
.B(n_2955),
.Y(n_3270)
);

INVxp67_ASAP7_75t_SL g3271 ( 
.A(n_3217),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3176),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3208),
.Y(n_3273)
);

NAND2x2_ASAP7_75t_L g3274 ( 
.A(n_3196),
.B(n_3020),
.Y(n_3274)
);

AOI32xp33_ASAP7_75t_L g3275 ( 
.A1(n_3180),
.A2(n_3000),
.A3(n_2777),
.B1(n_3081),
.B2(n_2734),
.Y(n_3275)
);

OAI322xp33_ASAP7_75t_L g3276 ( 
.A1(n_3214),
.A2(n_3158),
.A3(n_3153),
.B1(n_3040),
.B2(n_3031),
.C1(n_3065),
.C2(n_3047),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_3225),
.B(n_3167),
.Y(n_3277)
);

OA222x2_ASAP7_75t_L g3278 ( 
.A1(n_3221),
.A2(n_2955),
.B1(n_3081),
.B2(n_3026),
.C1(n_3022),
.C2(n_3050),
.Y(n_3278)
);

OR2x2_ASAP7_75t_L g3279 ( 
.A(n_3193),
.B(n_3111),
.Y(n_3279)
);

INVxp33_ASAP7_75t_L g3280 ( 
.A(n_3195),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3214),
.B(n_3122),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3213),
.B(n_3122),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3247),
.Y(n_3283)
);

INVx1_ASAP7_75t_SL g3284 ( 
.A(n_3242),
.Y(n_3284)
);

INVx1_ASAP7_75t_SL g3285 ( 
.A(n_3245),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3279),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3254),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3255),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3244),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3249),
.Y(n_3290)
);

NAND3xp33_ASAP7_75t_L g3291 ( 
.A(n_3239),
.B(n_3250),
.C(n_3275),
.Y(n_3291)
);

AOI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3239),
.A2(n_3118),
.B1(n_3088),
.B2(n_3043),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3256),
.Y(n_3293)
);

XNOR2x1_ASAP7_75t_L g3294 ( 
.A(n_3243),
.B(n_2769),
.Y(n_3294)
);

INVxp67_ASAP7_75t_SL g3295 ( 
.A(n_3235),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3258),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3233),
.B(n_3181),
.Y(n_3297)
);

OR2x2_ASAP7_75t_L g3298 ( 
.A(n_3227),
.B(n_3181),
.Y(n_3298)
);

INVxp67_ASAP7_75t_L g3299 ( 
.A(n_3251),
.Y(n_3299)
);

NAND2x1_ASAP7_75t_SL g3300 ( 
.A(n_3253),
.B(n_3195),
.Y(n_3300)
);

AND2x4_ASAP7_75t_L g3301 ( 
.A(n_3271),
.B(n_3194),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3259),
.Y(n_3302)
);

AOI211xp5_ASAP7_75t_L g3303 ( 
.A1(n_3228),
.A2(n_2878),
.B(n_2737),
.C(n_2721),
.Y(n_3303)
);

OAI21xp33_ASAP7_75t_SL g3304 ( 
.A1(n_3277),
.A2(n_3192),
.B(n_3170),
.Y(n_3304)
);

OAI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_3280),
.A2(n_3118),
.B1(n_3088),
.B2(n_3043),
.Y(n_3305)
);

XOR2x2_ASAP7_75t_L g3306 ( 
.A(n_3269),
.B(n_2806),
.Y(n_3306)
);

O2A1O1Ixp33_ASAP7_75t_L g3307 ( 
.A1(n_3238),
.A2(n_2732),
.B(n_2646),
.C(n_2894),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3231),
.B(n_3175),
.Y(n_3308)
);

OAI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3252),
.A2(n_2954),
.B(n_2833),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_3257),
.A2(n_3253),
.B(n_3278),
.Y(n_3310)
);

NOR2x1p5_ASAP7_75t_L g3311 ( 
.A(n_3278),
.B(n_2730),
.Y(n_3311)
);

AOI22xp5_ASAP7_75t_SL g3312 ( 
.A1(n_3270),
.A2(n_2768),
.B1(n_2900),
.B2(n_2854),
.Y(n_3312)
);

XOR2x2_ASAP7_75t_L g3313 ( 
.A(n_3274),
.B(n_2765),
.Y(n_3313)
);

NOR3xp33_ASAP7_75t_L g3314 ( 
.A(n_3276),
.B(n_2936),
.C(n_2844),
.Y(n_3314)
);

AOI211xp5_ASAP7_75t_SL g3315 ( 
.A1(n_3276),
.A2(n_3022),
.B(n_3050),
.C(n_3037),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3260),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3261),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3262),
.Y(n_3318)
);

NAND4xp25_ASAP7_75t_SL g3319 ( 
.A(n_3304),
.B(n_3291),
.C(n_3292),
.D(n_3310),
.Y(n_3319)
);

AOI22x1_ASAP7_75t_L g3320 ( 
.A1(n_3311),
.A2(n_2891),
.B1(n_2825),
.B2(n_2893),
.Y(n_3320)
);

OAI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3304),
.A2(n_2927),
.B(n_2954),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3292),
.A2(n_3268),
.B1(n_3118),
.B2(n_3270),
.Y(n_3322)
);

OAI21xp33_ASAP7_75t_SL g3323 ( 
.A1(n_3300),
.A2(n_3236),
.B(n_3264),
.Y(n_3323)
);

OAI221xp5_ASAP7_75t_L g3324 ( 
.A1(n_3315),
.A2(n_3268),
.B1(n_3234),
.B2(n_3240),
.C(n_3232),
.Y(n_3324)
);

AOI21xp33_ASAP7_75t_L g3325 ( 
.A1(n_3285),
.A2(n_2809),
.B(n_2763),
.Y(n_3325)
);

INVx1_ASAP7_75t_SL g3326 ( 
.A(n_3284),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3289),
.B(n_3263),
.Y(n_3327)
);

NOR2x1_ASAP7_75t_L g3328 ( 
.A(n_3294),
.B(n_2799),
.Y(n_3328)
);

OAI322xp33_ASAP7_75t_L g3329 ( 
.A1(n_3312),
.A2(n_3164),
.A3(n_3218),
.B1(n_3248),
.B2(n_3246),
.C1(n_3229),
.C2(n_3266),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_3301),
.A2(n_3237),
.B1(n_3088),
.B2(n_3281),
.Y(n_3330)
);

NOR3xp33_ASAP7_75t_SL g3331 ( 
.A(n_3305),
.B(n_2884),
.C(n_2864),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3298),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3301),
.B(n_3230),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3295),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3302),
.Y(n_3335)
);

O2A1O1Ixp33_ASAP7_75t_L g3336 ( 
.A1(n_3299),
.A2(n_3267),
.B(n_3273),
.C(n_3265),
.Y(n_3336)
);

INVxp67_ASAP7_75t_SL g3337 ( 
.A(n_3314),
.Y(n_3337)
);

OAI322xp33_ASAP7_75t_L g3338 ( 
.A1(n_3297),
.A2(n_3175),
.A3(n_3191),
.B1(n_3226),
.B2(n_3210),
.C1(n_3282),
.C2(n_3272),
.Y(n_3338)
);

OR2x2_ASAP7_75t_L g3339 ( 
.A(n_3308),
.B(n_3223),
.Y(n_3339)
);

OAI221xp5_ASAP7_75t_L g3340 ( 
.A1(n_3303),
.A2(n_2908),
.B1(n_2945),
.B2(n_2954),
.C(n_3070),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3316),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3290),
.B(n_3224),
.Y(n_3342)
);

OAI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3307),
.A2(n_2889),
.B(n_2869),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3317),
.Y(n_3344)
);

OAI22xp33_ASAP7_75t_SL g3345 ( 
.A1(n_3318),
.A2(n_3241),
.B1(n_3037),
.B2(n_2923),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3287),
.B(n_3171),
.Y(n_3346)
);

AO21x1_ASAP7_75t_L g3347 ( 
.A1(n_3293),
.A2(n_3079),
.B(n_3087),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3313),
.B(n_3043),
.Y(n_3348)
);

OAI221xp5_ASAP7_75t_L g3349 ( 
.A1(n_3309),
.A2(n_3288),
.B1(n_3306),
.B2(n_3283),
.C(n_3286),
.Y(n_3349)
);

INVxp67_ASAP7_75t_SL g3350 ( 
.A(n_3296),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3298),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3301),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3298),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_3297),
.B(n_3176),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_3285),
.B(n_3186),
.Y(n_3355)
);

OAI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_3315),
.A2(n_2877),
.B1(n_2880),
.B2(n_3219),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_L g3357 ( 
.A(n_3326),
.B(n_2861),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3321),
.B(n_3222),
.Y(n_3358)
);

OAI211xp5_ASAP7_75t_L g3359 ( 
.A1(n_3337),
.A2(n_2714),
.B(n_2802),
.C(n_2767),
.Y(n_3359)
);

INVx3_ASAP7_75t_SL g3360 ( 
.A(n_3326),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3332),
.B(n_3188),
.Y(n_3361)
);

AOI211xp5_ASAP7_75t_L g3362 ( 
.A1(n_3319),
.A2(n_2669),
.B(n_2898),
.C(n_2897),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3351),
.B(n_3353),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3334),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3350),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3342),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_3348),
.B(n_2861),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3321),
.B(n_3220),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3355),
.B(n_2929),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3327),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3354),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_3352),
.B(n_3085),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3328),
.A2(n_2799),
.B(n_2835),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3335),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3341),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_3323),
.B(n_2813),
.Y(n_3376)
);

NAND3xp33_ASAP7_75t_L g3377 ( 
.A(n_3343),
.B(n_2934),
.C(n_2641),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3349),
.B(n_2943),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_3345),
.B(n_2832),
.Y(n_3379)
);

AND2x4_ASAP7_75t_L g3380 ( 
.A(n_3331),
.B(n_3059),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3344),
.B(n_3212),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3346),
.Y(n_3382)
);

OR2x2_ASAP7_75t_L g3383 ( 
.A(n_3347),
.B(n_3212),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3360),
.B(n_3336),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3365),
.B(n_3339),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3370),
.B(n_3333),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3382),
.B(n_3366),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3371),
.Y(n_3388)
);

OAI211xp5_ASAP7_75t_SL g3389 ( 
.A1(n_3362),
.A2(n_3359),
.B(n_3364),
.C(n_3373),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3363),
.B(n_3330),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3376),
.A2(n_3320),
.B(n_3329),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3367),
.A2(n_3325),
.B(n_3322),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3363),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3374),
.B(n_3356),
.Y(n_3394)
);

INVxp67_ASAP7_75t_L g3395 ( 
.A(n_3357),
.Y(n_3395)
);

NOR2x1_ASAP7_75t_L g3396 ( 
.A(n_3379),
.B(n_3324),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3361),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3361),
.Y(n_3398)
);

AOI211x1_ASAP7_75t_L g3399 ( 
.A1(n_3358),
.A2(n_3340),
.B(n_3338),
.C(n_3066),
.Y(n_3399)
);

AOI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3378),
.A2(n_2974),
.B1(n_3058),
.B2(n_3057),
.Y(n_3400)
);

AOI211xp5_ASAP7_75t_L g3401 ( 
.A1(n_3377),
.A2(n_2947),
.B(n_2853),
.C(n_2868),
.Y(n_3401)
);

OAI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3375),
.A2(n_2835),
.B(n_2593),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3369),
.A2(n_2896),
.B(n_3025),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3380),
.A2(n_2928),
.B(n_2883),
.Y(n_3404)
);

INVx1_ASAP7_75t_SL g3405 ( 
.A(n_3384),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_SL g3406 ( 
.A(n_3388),
.B(n_3383),
.Y(n_3406)
);

NAND5xp2_ASAP7_75t_L g3407 ( 
.A(n_3391),
.B(n_3392),
.C(n_3402),
.D(n_3404),
.E(n_3403),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3395),
.A2(n_3381),
.B(n_3368),
.Y(n_3408)
);

OAI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_3399),
.A2(n_3380),
.B1(n_3381),
.B2(n_3372),
.Y(n_3409)
);

O2A1O1Ixp33_ASAP7_75t_L g3410 ( 
.A1(n_3389),
.A2(n_2565),
.B(n_2830),
.C(n_2567),
.Y(n_3410)
);

NAND3xp33_ASAP7_75t_SL g3411 ( 
.A(n_3402),
.B(n_2565),
.C(n_2744),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_3390),
.B(n_3072),
.Y(n_3412)
);

AOI322xp5_ASAP7_75t_L g3413 ( 
.A1(n_3396),
.A2(n_2982),
.A3(n_2984),
.B1(n_2985),
.B2(n_2986),
.C1(n_3061),
.C2(n_2473),
.Y(n_3413)
);

OAI211xp5_ASAP7_75t_L g3414 ( 
.A1(n_3394),
.A2(n_2715),
.B(n_2494),
.C(n_2624),
.Y(n_3414)
);

AOI22xp5_ASAP7_75t_L g3415 ( 
.A1(n_3397),
.A2(n_3060),
.B1(n_3021),
.B2(n_3005),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3398),
.A2(n_3060),
.B1(n_3021),
.B2(n_3005),
.Y(n_3416)
);

AOI221xp5_ASAP7_75t_L g3417 ( 
.A1(n_3393),
.A2(n_3028),
.B1(n_3045),
.B2(n_2899),
.C(n_3090),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3385),
.Y(n_3418)
);

AOI211xp5_ASAP7_75t_L g3419 ( 
.A1(n_3387),
.A2(n_2624),
.B(n_2521),
.C(n_3003),
.Y(n_3419)
);

AO21x1_ASAP7_75t_L g3420 ( 
.A1(n_3386),
.A2(n_2529),
.B(n_2492),
.Y(n_3420)
);

AOI221xp5_ASAP7_75t_L g3421 ( 
.A1(n_3401),
.A2(n_3028),
.B1(n_3045),
.B2(n_3018),
.C(n_3063),
.Y(n_3421)
);

AOI221xp5_ASAP7_75t_L g3422 ( 
.A1(n_3400),
.A2(n_3018),
.B1(n_2961),
.B2(n_2975),
.C(n_2996),
.Y(n_3422)
);

AOI32xp33_ASAP7_75t_L g3423 ( 
.A1(n_3389),
.A2(n_3072),
.A3(n_3007),
.B1(n_2989),
.B2(n_3004),
.Y(n_3423)
);

OAI211xp5_ASAP7_75t_SL g3424 ( 
.A1(n_3405),
.A2(n_2494),
.B(n_2521),
.C(n_2631),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3418),
.Y(n_3425)
);

O2A1O1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_3407),
.A2(n_2529),
.B(n_2492),
.C(n_2451),
.Y(n_3426)
);

NOR2x1_ASAP7_75t_L g3427 ( 
.A(n_3411),
.B(n_2883),
.Y(n_3427)
);

NOR3x1_ASAP7_75t_L g3428 ( 
.A(n_3414),
.B(n_3409),
.C(n_3423),
.Y(n_3428)
);

INVx2_ASAP7_75t_SL g3429 ( 
.A(n_3412),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3408),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3415),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3419),
.Y(n_3432)
);

AOI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3406),
.A2(n_2856),
.B1(n_2966),
.B2(n_3007),
.Y(n_3433)
);

AOI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3420),
.A2(n_2966),
.B1(n_2946),
.B2(n_2912),
.Y(n_3434)
);

OAI22xp5_ASAP7_75t_L g3435 ( 
.A1(n_3416),
.A2(n_3076),
.B1(n_3206),
.B2(n_3200),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3410),
.Y(n_3436)
);

OAI211xp5_ASAP7_75t_L g3437 ( 
.A1(n_3430),
.A2(n_3413),
.B(n_3417),
.C(n_3421),
.Y(n_3437)
);

AND2x4_ASAP7_75t_L g3438 ( 
.A(n_3429),
.B(n_3008),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_SL g3439 ( 
.A(n_3427),
.B(n_2680),
.Y(n_3439)
);

NOR2x1_ASAP7_75t_L g3440 ( 
.A(n_3425),
.B(n_3436),
.Y(n_3440)
);

NAND3xp33_ASAP7_75t_L g3441 ( 
.A(n_3426),
.B(n_3432),
.C(n_3427),
.Y(n_3441)
);

OA22x2_ASAP7_75t_L g3442 ( 
.A1(n_3431),
.A2(n_3422),
.B1(n_2928),
.B2(n_2924),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3428),
.Y(n_3443)
);

NOR2x1_ASAP7_75t_L g3444 ( 
.A(n_3424),
.B(n_2283),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3433),
.Y(n_3445)
);

OAI211xp5_ASAP7_75t_L g3446 ( 
.A1(n_3434),
.A2(n_2477),
.B(n_2402),
.C(n_2904),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3440),
.Y(n_3447)
);

CKINVDCx20_ASAP7_75t_R g3448 ( 
.A(n_3443),
.Y(n_3448)
);

CKINVDCx5p33_ASAP7_75t_R g3449 ( 
.A(n_3445),
.Y(n_3449)
);

CKINVDCx5p33_ASAP7_75t_R g3450 ( 
.A(n_3441),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3438),
.Y(n_3451)
);

INVxp67_ASAP7_75t_L g3452 ( 
.A(n_3447),
.Y(n_3452)
);

INVx1_ASAP7_75t_SL g3453 ( 
.A(n_3449),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3448),
.A2(n_3442),
.B1(n_3437),
.B2(n_3435),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3451),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3450),
.Y(n_3456)
);

OAI31xp33_ASAP7_75t_L g3457 ( 
.A1(n_3453),
.A2(n_3446),
.A3(n_3439),
.B(n_3444),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3455),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3454),
.A2(n_2680),
.B1(n_2681),
.B2(n_2690),
.Y(n_3459)
);

AOI211xp5_ASAP7_75t_L g3460 ( 
.A1(n_3452),
.A2(n_2690),
.B(n_2681),
.C(n_2295),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3458),
.Y(n_3461)
);

INVxp67_ASAP7_75t_L g3462 ( 
.A(n_3459),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3461),
.Y(n_3463)
);

AOI21x1_ASAP7_75t_L g3464 ( 
.A1(n_3463),
.A2(n_3456),
.B(n_3457),
.Y(n_3464)
);

NAND3xp33_ASAP7_75t_L g3465 ( 
.A(n_3463),
.B(n_3462),
.C(n_3460),
.Y(n_3465)
);

AOI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3465),
.A2(n_3464),
.B1(n_3091),
.B2(n_2726),
.Y(n_3466)
);

AOI221xp5_ASAP7_75t_L g3467 ( 
.A1(n_3466),
.A2(n_2690),
.B1(n_2681),
.B2(n_2726),
.C(n_2924),
.Y(n_3467)
);

AOI22xp5_ASAP7_75t_L g3468 ( 
.A1(n_3467),
.A2(n_2370),
.B1(n_2375),
.B2(n_2804),
.Y(n_3468)
);


endmodule