module real_aes_1418_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_0), .B(n_197), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_1), .A2(n_180), .B(n_230), .Y(n_229) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_2), .A2(n_55), .B1(n_89), .B2(n_102), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_3), .B(n_187), .Y(n_243) );
INVx1_ASAP7_75t_L g163 ( .A(n_4), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_5), .B(n_187), .Y(n_207) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_6), .A2(n_21), .B1(n_89), .B2(n_99), .Y(n_98) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_7), .B(n_191), .Y(n_224) );
INVx2_ASAP7_75t_L g177 ( .A(n_8), .Y(n_177) );
AOI221x1_ASAP7_75t_L g266 ( .A1(n_9), .A2(n_17), .B1(n_180), .B2(n_197), .C(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_10), .B(n_197), .Y(n_220) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_11), .A2(n_218), .B(n_219), .Y(n_217) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_12), .A2(n_65), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_12), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_13), .B(n_210), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_14), .B(n_187), .Y(n_186) );
AO21x1_ASAP7_75t_L g238 ( .A1(n_15), .A2(n_197), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g492 ( .A(n_16), .Y(n_492) );
NAND2x1_ASAP7_75t_L g252 ( .A(n_18), .B(n_187), .Y(n_252) );
NAND2x1_ASAP7_75t_L g206 ( .A(n_19), .B(n_191), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_20), .A2(n_48), .B1(n_118), .B2(n_120), .Y(n_117) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_21), .A2(n_55), .B1(n_59), .B2(n_503), .C(n_505), .Y(n_502) );
OR2x2_ASAP7_75t_L g176 ( .A(n_22), .B(n_67), .Y(n_176) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_22), .A2(n_67), .B(n_177), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_23), .A2(n_39), .B1(n_124), .B2(n_128), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_24), .A2(n_71), .B1(n_133), .B2(n_135), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_25), .B(n_191), .Y(n_232) );
INVx3_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_27), .B(n_187), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_28), .B(n_191), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_29), .A2(n_180), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g527 ( .A(n_29), .Y(n_527) );
INVx1_ASAP7_75t_SL g94 ( .A(n_30), .Y(n_94) );
INVx1_ASAP7_75t_L g165 ( .A(n_31), .Y(n_165) );
AND2x2_ASAP7_75t_L g181 ( .A(n_31), .B(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g195 ( .A(n_31), .B(n_163), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_32), .B(n_197), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_33), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_34), .B(n_191), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_34), .A2(n_487), .B1(n_501), .B2(n_509), .Y(n_486) );
INVx1_ASAP7_75t_L g517 ( .A(n_34), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_35), .A2(n_63), .B1(n_140), .B2(n_142), .Y(n_139) );
AOI22xp33_ASAP7_75t_SL g147 ( .A1(n_36), .A2(n_62), .B1(n_148), .B2(n_150), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_37), .A2(n_180), .B(n_205), .Y(n_204) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_38), .A2(n_59), .B1(n_89), .B2(n_90), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_40), .B(n_191), .Y(n_253) );
INVx1_ASAP7_75t_L g184 ( .A(n_41), .Y(n_184) );
INVx1_ASAP7_75t_L g193 ( .A(n_41), .Y(n_193) );
INVx1_ASAP7_75t_L g95 ( .A(n_42), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_43), .B(n_155), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_44), .A2(n_80), .B1(n_158), .B2(n_159), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_44), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_45), .B(n_187), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_46), .A2(n_180), .B(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_47), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_47), .Y(n_493) );
AO21x1_ASAP7_75t_L g240 ( .A1(n_49), .A2(n_180), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_50), .B(n_197), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g83 ( .A1(n_51), .A2(n_53), .B1(n_84), .B2(n_103), .Y(n_83) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_52), .A2(n_66), .B1(n_111), .B2(n_114), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_54), .B(n_197), .Y(n_208) );
INVxp33_ASAP7_75t_L g507 ( .A(n_55), .Y(n_507) );
AND2x2_ASAP7_75t_L g289 ( .A(n_56), .B(n_211), .Y(n_289) );
INVx1_ASAP7_75t_L g182 ( .A(n_57), .Y(n_182) );
INVx1_ASAP7_75t_L g189 ( .A(n_57), .Y(n_189) );
AND2x2_ASAP7_75t_L g212 ( .A(n_58), .B(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g506 ( .A(n_59), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_60), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g226 ( .A(n_61), .B(n_213), .Y(n_226) );
AND2x2_ASAP7_75t_L g239 ( .A(n_64), .B(n_175), .Y(n_239) );
INVx1_ASAP7_75t_L g498 ( .A(n_65), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_68), .B(n_191), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_68), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_68), .Y(n_495) );
AND2x2_ASAP7_75t_L g256 ( .A(n_69), .B(n_213), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_70), .B(n_187), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_72), .A2(n_180), .B(n_185), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_73), .B(n_191), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_74), .B(n_187), .Y(n_231) );
BUFx2_ASAP7_75t_SL g504 ( .A(n_75), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_76), .A2(n_180), .B(n_222), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_160), .B1(n_166), .B2(n_483), .C(n_485), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
INVx1_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
OAI222xp33_ASAP7_75t_R g485 ( .A1(n_80), .A2(n_159), .B1(n_486), .B2(n_514), .C1(n_519), .C2(n_527), .Y(n_485) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_131), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_110), .C(n_117), .D(n_123), .Y(n_82) );
INVx2_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
INVx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_96), .Y(n_86) );
AND2x2_ASAP7_75t_L g119 ( .A(n_87), .B(n_108), .Y(n_119) );
AND2x4_ASAP7_75t_L g141 ( .A(n_87), .B(n_116), .Y(n_141) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
INVx2_ASAP7_75t_L g107 ( .A(n_88), .Y(n_107) );
BUFx2_ASAP7_75t_L g121 ( .A(n_88), .Y(n_121) );
AND2x2_ASAP7_75t_L g146 ( .A(n_88), .B(n_92), .Y(n_146) );
INVx1_ASAP7_75t_L g90 ( .A(n_89), .Y(n_90) );
OAI22x1_ASAP7_75t_L g92 ( .A1(n_89), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx2_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
INVx1_ASAP7_75t_L g102 ( .A(n_89), .Y(n_102) );
AND2x4_ASAP7_75t_L g106 ( .A(n_91), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g127 ( .A(n_92), .B(n_107), .Y(n_127) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
AND2x4_ASAP7_75t_L g113 ( .A(n_96), .B(n_106), .Y(n_113) );
AND2x4_ASAP7_75t_L g126 ( .A(n_96), .B(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g157 ( .A(n_96), .B(n_146), .Y(n_157) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_100), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx1_ASAP7_75t_L g109 ( .A(n_98), .Y(n_109) );
AND2x4_ASAP7_75t_L g116 ( .A(n_98), .B(n_100), .Y(n_116) );
AND2x2_ASAP7_75t_L g122 ( .A(n_98), .B(n_101), .Y(n_122) );
INVxp67_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g108 ( .A(n_101), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx8_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x4_ASAP7_75t_L g115 ( .A(n_106), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g130 ( .A(n_106), .B(n_122), .Y(n_130) );
AND2x2_ASAP7_75t_L g149 ( .A(n_108), .B(n_127), .Y(n_149) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx8_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g134 ( .A(n_116), .B(n_127), .Y(n_134) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x2_ASAP7_75t_L g137 ( .A(n_122), .B(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx6_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_139), .C(n_147), .D(n_154), .Y(n_131) );
BUFx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
INVx6_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g151 ( .A(n_146), .B(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx4f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx6_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g508 ( .A(n_162), .Y(n_508) );
AND2x2_ASAP7_75t_L g525 ( .A(n_162), .B(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g183 ( .A(n_163), .B(n_184), .Y(n_183) );
AND3x1_ASAP7_75t_SL g501 ( .A(n_164), .B(n_502), .C(n_508), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_164), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_381), .Y(n_167) );
NAND3xp33_ASAP7_75t_SL g168 ( .A(n_169), .B(n_293), .C(n_348), .Y(n_168) );
AOI221xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_233), .B1(n_257), .B2(n_261), .C(n_271), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_216), .Y(n_170) );
AND2x2_ASAP7_75t_SL g259 ( .A(n_171), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g292 ( .A(n_171), .Y(n_292) );
AND2x2_ASAP7_75t_L g337 ( .A(n_171), .B(n_274), .Y(n_337) );
AND2x4_ASAP7_75t_L g171 ( .A(n_172), .B(n_201), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g325 ( .A(n_173), .Y(n_325) );
INVx1_ASAP7_75t_L g335 ( .A(n_173), .Y(n_335) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_178), .B(n_199), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_174), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_174), .A2(n_178), .B(n_199), .Y(n_299) );
INVx1_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_175), .A2(n_220), .B(n_221), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_175), .B(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_176), .B(n_177), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_196), .Y(n_178) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_180), .Y(n_484) );
AND2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_183), .Y(n_180) );
BUFx3_ASAP7_75t_L g523 ( .A(n_181), .Y(n_523) );
AND2x6_ASAP7_75t_L g191 ( .A(n_182), .B(n_192), .Y(n_191) );
AND2x4_ASAP7_75t_L g187 ( .A(n_184), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g526 ( .A(n_184), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_190), .B(n_194), .Y(n_185) );
AND2x4_ASAP7_75t_L g198 ( .A(n_188), .B(n_192), .Y(n_198) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_194), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_194), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_194), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_194), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_194), .A2(n_252), .B(n_253), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_194), .A2(n_268), .B(n_269), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_194), .A2(n_286), .B(n_287), .Y(n_285) );
INVx5_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x4_ASAP7_75t_L g197 ( .A(n_195), .B(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g314 ( .A(n_201), .B(n_217), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_201), .B(n_260), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_201), .B(n_225), .Y(n_358) );
INVx2_ASAP7_75t_L g367 ( .A(n_201), .Y(n_367) );
AND2x2_ASAP7_75t_L g388 ( .A(n_201), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g472 ( .A(n_201), .B(n_291), .Y(n_472) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g300 ( .A(n_202), .B(n_225), .Y(n_300) );
AND2x2_ASAP7_75t_L g433 ( .A(n_202), .B(n_260), .Y(n_433) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_202), .Y(n_459) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_209), .B(n_212), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_208), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_210), .A2(n_228), .B(n_229), .Y(n_227) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_210), .A2(n_266), .B(n_270), .Y(n_265) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_210), .A2(n_266), .B(n_270), .Y(n_277) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
INVx4_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_215), .Y(n_218) );
AND2x4_ASAP7_75t_L g387 ( .A(n_216), .B(n_388), .Y(n_387) );
AOI321xp33_ASAP7_75t_L g401 ( .A1(n_216), .A2(n_330), .A3(n_331), .B1(n_363), .B2(n_402), .C(n_405), .Y(n_401) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_225), .Y(n_216) );
BUFx3_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
INVx2_ASAP7_75t_L g291 ( .A(n_217), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_217), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g324 ( .A(n_217), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g357 ( .A(n_217), .Y(n_357) );
INVx5_ASAP7_75t_L g260 ( .A(n_225), .Y(n_260) );
NOR2x1_ASAP7_75t_SL g309 ( .A(n_225), .B(n_299), .Y(n_309) );
BUFx2_ASAP7_75t_L g404 ( .A(n_225), .Y(n_404) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVxp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_246), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_235), .B(n_303), .Y(n_302) );
NOR4xp25_ASAP7_75t_L g405 ( .A(n_235), .B(n_399), .C(n_403), .D(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g443 ( .A(n_235), .Y(n_443) );
AND2x2_ASAP7_75t_L g477 ( .A(n_235), .B(n_417), .Y(n_477) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g332 ( .A(n_237), .Y(n_332) );
OAI21x1_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_240), .B(n_244), .Y(n_237) );
INVx1_ASAP7_75t_L g245 ( .A(n_239), .Y(n_245) );
AOI33xp33_ASAP7_75t_L g473 ( .A1(n_246), .A2(n_275), .A3(n_306), .B1(n_322), .B2(n_428), .B3(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g263 ( .A(n_247), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g273 ( .A(n_247), .B(n_274), .Y(n_273) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
INVxp67_ASAP7_75t_L g361 ( .A(n_248), .Y(n_361) );
AND2x2_ASAP7_75t_L g417 ( .A(n_248), .B(n_282), .Y(n_417) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_255), .B(n_256), .Y(n_248) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_249), .A2(n_255), .B(n_256), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_255), .A2(n_283), .B(n_289), .Y(n_282) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_255), .A2(n_283), .B(n_289), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_257), .A2(n_439), .B(n_440), .Y(n_438) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g426 ( .A(n_258), .B(n_300), .Y(n_426) );
AND3x2_ASAP7_75t_L g428 ( .A(n_258), .B(n_312), .C(n_367), .Y(n_428) );
INVx3_ASAP7_75t_SL g380 ( .A(n_259), .Y(n_380) );
INVx4_ASAP7_75t_L g274 ( .A(n_260), .Y(n_274) );
AND2x2_ASAP7_75t_L g312 ( .A(n_260), .B(n_299), .Y(n_312) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g306 ( .A(n_264), .Y(n_306) );
AND2x4_ASAP7_75t_L g331 ( .A(n_264), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g394 ( .A(n_264), .B(n_282), .Y(n_394) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g364 ( .A(n_265), .Y(n_364) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_265), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_R g271 ( .A1(n_272), .A2(n_275), .B(n_279), .C(n_290), .Y(n_271) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g323 ( .A(n_274), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_274), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_274), .B(n_291), .Y(n_452) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g434 ( .A(n_276), .B(n_424), .Y(n_434) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_277), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g303 ( .A(n_277), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g319 ( .A(n_277), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g352 ( .A(n_277), .B(n_332), .Y(n_352) );
AND2x4_ASAP7_75t_L g317 ( .A(n_278), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g341 ( .A(n_278), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g379 ( .A(n_278), .B(n_304), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g307 ( .A(n_280), .B(n_304), .Y(n_307) );
AND2x2_ASAP7_75t_L g322 ( .A(n_280), .B(n_282), .Y(n_322) );
BUFx2_ASAP7_75t_L g378 ( .A(n_280), .Y(n_378) );
AND2x2_ASAP7_75t_L g392 ( .A(n_280), .B(n_303), .Y(n_392) );
INVx2_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_288), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_290), .A2(n_341), .B1(n_343), .B2(n_347), .Y(n_340) );
INVx2_ASAP7_75t_SL g371 ( .A(n_290), .Y(n_371) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g346 ( .A(n_291), .B(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g453 ( .A(n_292), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_326), .C(n_340), .Y(n_293) );
OAI221xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_301), .B1(n_305), .B2(n_308), .C(n_310), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVxp67_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g354 ( .A(n_298), .Y(n_354) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_298), .Y(n_482) );
INVx1_ASAP7_75t_L g445 ( .A(n_300), .Y(n_445) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_300), .B(n_324), .Y(n_455) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_304), .B(n_332), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OR2x2_ASAP7_75t_L g338 ( .A(n_306), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g416 ( .A(n_306), .Y(n_416) );
AND2x2_ASAP7_75t_L g351 ( .A(n_307), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g397 ( .A(n_309), .B(n_357), .Y(n_397) );
AND2x2_ASAP7_75t_L g474 ( .A(n_309), .B(n_472), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .B1(n_322), .B2(n_323), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx2_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
AND2x4_ASAP7_75t_L g363 ( .A(n_317), .B(n_364), .Y(n_363) );
OAI21xp33_ASAP7_75t_SL g393 ( .A1(n_317), .A2(n_394), .B(n_395), .Y(n_393) );
AND2x2_ASAP7_75t_L g420 ( .A(n_317), .B(n_378), .Y(n_420) );
INVx2_ASAP7_75t_L g342 ( .A(n_318), .Y(n_342) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_318), .Y(n_375) );
INVx1_ASAP7_75t_SL g399 ( .A(n_319), .Y(n_399) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g330 ( .A(n_321), .Y(n_330) );
AND2x4_ASAP7_75t_SL g424 ( .A(n_321), .B(n_342), .Y(n_424) );
AND2x2_ASAP7_75t_L g421 ( .A(n_324), .B(n_367), .Y(n_421) );
AND2x2_ASAP7_75t_L g447 ( .A(n_324), .B(n_433), .Y(n_447) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_325), .Y(n_369) );
INVx1_ASAP7_75t_L g389 ( .A(n_325), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_333), .B1(n_336), .B2(n_338), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_331), .B(n_342), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_331), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g470 ( .A(n_331), .Y(n_470) );
INVx2_ASAP7_75t_SL g395 ( .A(n_333), .Y(n_395) );
AND2x2_ASAP7_75t_L g407 ( .A(n_335), .B(n_367), .Y(n_407) );
INVx2_ASAP7_75t_L g413 ( .A(n_335), .Y(n_413) );
INVxp33_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_341), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g463 ( .A(n_341), .Y(n_463) );
INVx1_ASAP7_75t_L g391 ( .A(n_343), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_344), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g402 ( .A(n_346), .B(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_346), .A2(n_476), .B1(n_477), .B2(n_478), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_370), .C(n_373), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B1(n_355), .B2(n_359), .C(n_362), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g468 ( .A(n_353), .Y(n_468) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g437 ( .A(n_354), .B(n_403), .Y(n_437) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g368 ( .A(n_357), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g439 ( .A(n_359), .Y(n_439) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g436 ( .A(n_360), .Y(n_436) );
INVx1_ASAP7_75t_L g442 ( .A(n_361), .Y(n_442) );
OR2x2_ASAP7_75t_L g465 ( .A(n_361), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_SL g374 ( .A(n_364), .Y(n_374) );
AND2x2_ASAP7_75t_L g444 ( .A(n_364), .B(n_424), .Y(n_444) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_364), .B(n_377), .Y(n_476) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g481 ( .A(n_367), .Y(n_481) );
INVx1_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_376), .C(n_380), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_374), .B(n_424), .Y(n_448) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_377), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g385 ( .A(n_379), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g466 ( .A(n_379), .Y(n_466) );
NAND4xp75_ASAP7_75t_L g381 ( .A(n_382), .B(n_438), .C(n_454), .D(n_475), .Y(n_381) );
NOR3x1_ASAP7_75t_L g382 ( .A(n_383), .B(n_400), .C(n_422), .Y(n_382) );
NAND4xp75_ASAP7_75t_L g383 ( .A(n_384), .B(n_390), .C(n_393), .D(n_396), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_387), .Y(n_384) );
AND2x2_ASAP7_75t_L g435 ( .A(n_386), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g460 ( .A(n_387), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g449 ( .A(n_392), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_408), .Y(n_400) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_404), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_414), .B(n_418), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI322xp33_ASAP7_75t_L g440 ( .A1(n_412), .A2(n_441), .A3(n_445), .B1(n_446), .B2(n_448), .C1(n_449), .C2(n_450), .Y(n_440) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_413), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_416), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_417), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B(n_427), .C(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_434), .B1(n_435), .B2(n_437), .Y(n_429) );
NOR2xp33_ASAP7_75t_SL g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B(n_444), .Y(n_441) );
INVxp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_447), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_453), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g457 ( .A(n_452), .B(n_458), .Y(n_457) );
O2A1O1Ixp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_461), .C(n_464), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI221xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_467), .B1(n_469), .B2(n_471), .C(n_473), .Y(n_464) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_488), .A2(n_515), .B1(n_517), .B2(n_518), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_494), .B2(n_500), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_494), .Y(n_500) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_501), .Y(n_516) );
INVxp67_ASAP7_75t_L g513 ( .A(n_502), .Y(n_513) );
CKINVDCx8_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_508), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_508), .A2(n_521), .B(n_524), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_510), .Y(n_518) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
INVxp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
endmodule