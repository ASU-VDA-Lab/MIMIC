module fake_jpeg_2099_n_203 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_35),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_17),
.A2(n_10),
.B(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_2),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_51),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_50),
.B1(n_59),
.B2(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_80),
.B1(n_54),
.B2(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_62),
.B1(n_59),
.B2(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_86),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_57),
.B1(n_48),
.B2(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_89),
.B1(n_46),
.B2(n_58),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_67),
.B1(n_49),
.B2(n_53),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_58),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_48),
.B1(n_57),
.B2(n_65),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_67),
.B1(n_49),
.B2(n_63),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_52),
.C(n_47),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_69),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_94),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_3),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_102),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_101),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_44),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_74),
.A3(n_66),
.B1(n_61),
.B2(n_54),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_83),
.B1(n_82),
.B2(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_2),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_54),
.B1(n_61),
.B2(n_74),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_90),
.B(n_74),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_109),
.B(n_34),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_127),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_12),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_12),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_42),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_6),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_100),
.B1(n_109),
.B2(n_98),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_145),
.B1(n_28),
.B2(n_18),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_142),
.B(n_135),
.C(n_150),
.D(n_140),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_142),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_54),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_139),
.C(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_40),
.C(n_37),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_148),
.C(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_30),
.B(n_11),
.Y(n_146)
);

NOR4xp25_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_19),
.C(n_20),
.D(n_21),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_7),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_15),
.C(n_16),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_156),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_158),
.C(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_14),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_14),
.B(n_15),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_24),
.B(n_28),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_22),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_16),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_18),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_20),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_22),
.C(n_23),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_149),
.C(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_174),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_23),
.A3(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_178),
.Y(n_189)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_164),
.C(n_157),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_162),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_187),
.C(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_180),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_170),
.Y(n_187)
);

OAI322xp33_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_155),
.A3(n_159),
.B1(n_160),
.B2(n_163),
.C1(n_168),
.C2(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_190),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_182),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_178),
.B(n_179),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_174),
.A3(n_183),
.B1(n_184),
.B2(n_185),
.C1(n_187),
.C2(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

OA21x2_ASAP7_75t_SL g202 ( 
.A1(n_201),
.A2(n_199),
.B(n_198),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_202),
.Y(n_203)
);


endmodule