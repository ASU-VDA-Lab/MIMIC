module fake_jpeg_23153_n_230 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_36),
.B1(n_21),
.B2(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_31),
.B1(n_21),
.B2(n_18),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_40),
.B1(n_46),
.B2(n_50),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_31),
.B1(n_21),
.B2(n_14),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_34),
.B(n_32),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_14),
.B1(n_21),
.B2(n_16),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_18),
.B1(n_16),
.B2(n_23),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_49),
.B(n_13),
.C(n_29),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_18),
.B1(n_16),
.B2(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_14),
.B1(n_25),
.B2(n_24),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_25),
.C(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_29),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_66),
.Y(n_72)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_54),
.B(n_55),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_20),
.B1(n_25),
.B2(n_19),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_13),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_20),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_37),
.B1(n_51),
.B2(n_38),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_55),
.B1(n_63),
.B2(n_57),
.Y(n_93)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_81),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_38),
.B1(n_40),
.B2(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_82),
.B1(n_65),
.B2(n_69),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_51),
.C(n_43),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_42),
.C(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_88),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_19),
.B(n_15),
.Y(n_95)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_55),
.B(n_62),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_74),
.B(n_80),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_104),
.B1(n_107),
.B2(n_73),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_87),
.B1(n_76),
.B2(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_89),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_42),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_100),
.C(n_102),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_74),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_35),
.C(n_25),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_13),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_72),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_75),
.B1(n_80),
.B2(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_68),
.B1(n_64),
.B2(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_129),
.B(n_95),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_125),
.B1(n_93),
.B2(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_79),
.C(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

OAI211xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_112),
.B(n_114),
.C(n_28),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_90),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_90),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_72),
.B1(n_82),
.B2(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_67),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_120),
.C(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_106),
.B1(n_92),
.B2(n_107),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_103),
.B1(n_100),
.B2(n_79),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_67),
.B1(n_28),
.B2(n_15),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_149),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_86),
.B(n_19),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_114),
.B(n_128),
.C(n_116),
.D(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_148),
.C(n_139),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_15),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_28),
.B1(n_13),
.B2(n_17),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_162),
.B1(n_156),
.B2(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_166),
.C(n_132),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_24),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_130),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_140),
.B(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_17),
.B(n_1),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_17),
.C(n_26),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_176),
.B1(n_26),
.B2(n_17),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_158),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_161),
.B(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_163),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_142),
.B1(n_131),
.B2(n_143),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_177),
.B(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_141),
.C(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_173),
.C(n_176),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_186),
.C(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_7),
.B(n_9),
.Y(n_201)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_185),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_135),
.C(n_164),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_172),
.C(n_170),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_17),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_170),
.C(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.C(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_168),
.C(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_174),
.C(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_209),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_185),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_6),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_183),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_197),
.C(n_202),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_204),
.B(n_210),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_26),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_208),
.A2(n_7),
.B(n_12),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_5),
.C(n_11),
.Y(n_218)
);

OAI21x1_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_10),
.B(n_11),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_216),
.B(n_5),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_220),
.A2(n_216),
.B(n_215),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_223),
.B(n_224),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_221),
.B(n_10),
.C(n_11),
.D(n_4),
.Y(n_225)
);

NOR4xp25_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_10),
.C(n_1),
.D(n_3),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_226),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_0),
.B(n_3),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_4),
.B(n_26),
.Y(n_230)
);


endmodule