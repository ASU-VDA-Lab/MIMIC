module fake_jpeg_27570_n_133 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_0),
.B(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_4),
.A2(n_1),
.B(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_36),
.B1(n_28),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_49),
.B1(n_30),
.B2(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.C(n_17),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_27),
.C(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_18),
.B1(n_24),
.B2(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_63),
.B1(n_49),
.B2(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_42),
.B1(n_44),
.B2(n_37),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_2),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_46),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_30),
.B1(n_33),
.B2(n_13),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_40),
.B1(n_14),
.B2(n_13),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_40),
.B1(n_53),
.B2(n_62),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_42),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_41),
.C(n_45),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_55),
.C(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_61),
.B1(n_59),
.B2(n_63),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_83),
.B(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_72),
.C(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_91),
.B1(n_65),
.B2(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_98),
.B1(n_101),
.B2(n_71),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_70),
.B(n_76),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_84),
.B1(n_89),
.B2(n_19),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_81),
.B1(n_66),
.B2(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_33),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_71),
.B1(n_74),
.B2(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_91),
.B1(n_76),
.B2(n_85),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_100),
.A3(n_76),
.B1(n_93),
.B2(n_69),
.C1(n_99),
.C2(n_95),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

OA21x2_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_94),
.B(n_16),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_33),
.C(n_14),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_117),
.C(n_105),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_19),
.B1(n_33),
.B2(n_6),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_110),
.C(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_119),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_112),
.B1(n_103),
.B2(n_115),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_120),
.B1(n_5),
.B2(n_6),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_4),
.B(n_5),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_7),
.B(n_9),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_125),
.B(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_122),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_9),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_118),
.B1(n_9),
.B2(n_10),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_129),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_131),
.Y(n_133)
);


endmodule