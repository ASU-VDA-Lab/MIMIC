module fake_jpeg_30963_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_54),
.Y(n_103)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_53),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_55),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_18),
.B1(n_47),
.B2(n_21),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_58),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_62),
.Y(n_109)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_81),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_31),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_77),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_22),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_88),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_99),
.Y(n_145)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_36),
.B(n_15),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_44),
.Y(n_154)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_24),
.B(n_23),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_102),
.B(n_60),
.C(n_66),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_42),
.B1(n_37),
.B2(n_36),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_104),
.A2(n_116),
.B1(n_118),
.B2(n_120),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_51),
.A2(n_18),
.B1(n_47),
.B2(n_21),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_48),
.B1(n_39),
.B2(n_45),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_42),
.B1(n_37),
.B2(n_26),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_124),
.B(n_135),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_22),
.B1(n_45),
.B2(n_43),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_137),
.B1(n_67),
.B2(n_55),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_72),
.A2(n_26),
.B1(n_49),
.B2(n_34),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_84),
.A2(n_43),
.B1(n_39),
.B2(n_29),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_62),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_15),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_80),
.A2(n_44),
.B1(n_29),
.B2(n_25),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_147),
.A2(n_44),
.B1(n_83),
.B2(n_92),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_56),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_33),
.Y(n_203)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_33),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_102),
.A2(n_128),
.B(n_136),
.C(n_109),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_206),
.B(n_125),
.C(n_115),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_68),
.B1(n_64),
.B2(n_61),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_166),
.A2(n_182),
.B1(n_190),
.B2(n_95),
.Y(n_243)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_171),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_169),
.B(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_105),
.B(n_98),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_11),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_175),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_119),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_178),
.Y(n_225)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_120),
.A2(n_79),
.B1(n_63),
.B2(n_78),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_90),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_198),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_130),
.B(n_12),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_185),
.B(n_32),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_101),
.B1(n_94),
.B2(n_75),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_65),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_203),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_12),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_140),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_194),
.B(n_196),
.Y(n_235)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_140),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_210),
.B1(n_125),
.B2(n_107),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_111),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_134),
.B(n_11),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_200),
.B(n_205),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_134),
.A2(n_157),
.B(n_147),
.C(n_133),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_201),
.A2(n_146),
.B(n_127),
.C(n_150),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_123),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_122),
.B(n_44),
.Y(n_205)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_91),
.B1(n_44),
.B2(n_85),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_117),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_106),
.B(n_33),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_212),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_33),
.B1(n_32),
.B2(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_216),
.B(n_252),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_163),
.A2(n_141),
.B1(n_150),
.B2(n_121),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_226),
.A2(n_132),
.B1(n_112),
.B2(n_194),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_242),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_233),
.B(n_241),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_146),
.C(n_155),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_191),
.C(n_188),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_164),
.Y(n_241)
);

AOI22x1_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_157),
.B1(n_107),
.B2(n_141),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_162),
.B1(n_127),
.B2(n_174),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_113),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_248),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_183),
.A2(n_32),
.B(n_3),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_108),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_185),
.B(n_113),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_209),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_203),
.B(n_163),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_161),
.B(n_213),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_192),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_212),
.B(n_196),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_161),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_112),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_257),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_274),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_190),
.B1(n_182),
.B2(n_168),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_261),
.A2(n_272),
.B1(n_283),
.B2(n_284),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_165),
.B1(n_178),
.B2(n_206),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_262),
.A2(n_279),
.B1(n_280),
.B2(n_247),
.Y(n_310)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_266),
.A2(n_239),
.B(n_235),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_273),
.B(n_215),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_173),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_268),
.B(n_278),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_269),
.B(n_285),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_281),
.C(n_253),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_233),
.B(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_296),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_242),
.A2(n_228),
.B1(n_232),
.B2(n_254),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_229),
.A2(n_181),
.B1(n_208),
.B2(n_132),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_229),
.A2(n_180),
.B1(n_160),
.B2(n_177),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_204),
.C(n_189),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_195),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_282),
.B(n_293),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_214),
.A2(n_187),
.B1(n_186),
.B2(n_167),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_214),
.A2(n_238),
.B(n_244),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_215),
.B(n_239),
.Y(n_306)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_228),
.A2(n_179),
.B1(n_161),
.B2(n_32),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_223),
.B1(n_234),
.B2(n_252),
.Y(n_304)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_216),
.A2(n_179),
.B1(n_5),
.B2(n_6),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_292),
.B1(n_7),
.B2(n_8),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_243),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_294),
.B(n_295),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_257),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_304),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_300),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_330),
.Y(n_344)
);

A2O1A1O1Ixp25_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_255),
.B(n_224),
.C(n_239),
.D(n_258),
.Y(n_308)
);

OA21x2_ASAP7_75t_SL g357 ( 
.A1(n_308),
.A2(n_290),
.B(n_289),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_309),
.A2(n_240),
.B(n_230),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_317),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_298),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_258),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_329),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_273),
.A2(n_247),
.B(n_223),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_297),
.B(n_271),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_263),
.A2(n_259),
.B(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_324),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_261),
.A2(n_237),
.B1(n_234),
.B2(n_231),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_280),
.B1(n_279),
.B2(n_271),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_321),
.C(n_325),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_231),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_241),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_270),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_259),
.B(n_217),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_328),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_217),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_298),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_218),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_269),
.B(n_218),
.CI(n_219),
.CON(n_331),
.SN(n_331)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_333),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_265),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_230),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_263),
.B(n_278),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_337),
.A2(n_343),
.B(n_350),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_362),
.B1(n_310),
.B2(n_321),
.Y(n_379)
);

OAI22x1_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_263),
.B1(n_295),
.B2(n_267),
.Y(n_342)
);

OA22x2_ASAP7_75t_L g382 ( 
.A1(n_342),
.A2(n_348),
.B1(n_312),
.B2(n_331),
.Y(n_382)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

AO21x2_ASAP7_75t_L g348 ( 
.A1(n_315),
.A2(n_292),
.B(n_272),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_311),
.A2(n_262),
.B(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_296),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_320),
.C(n_332),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_294),
.B(n_293),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_365),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_306),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_322),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_359),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_302),
.A2(n_287),
.B1(n_264),
.B2(n_237),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_309),
.B(n_240),
.Y(n_363)
);

AND2x4_ASAP7_75t_SL g374 ( 
.A(n_363),
.B(n_331),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_364),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_302),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_366),
.A2(n_367),
.B1(n_307),
.B2(n_316),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_323),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_375),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_355),
.C(n_335),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_375),
.C(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_347),
.B(n_300),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_367),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_372),
.B(n_396),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_374),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_330),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_346),
.A2(n_312),
.B1(n_327),
.B2(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_332),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_395),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_379),
.A2(n_388),
.B1(n_389),
.B2(n_392),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_382),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_317),
.B1(n_307),
.B2(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_346),
.A2(n_316),
.B1(n_313),
.B2(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_350),
.A2(n_313),
.B1(n_305),
.B2(n_303),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_336),
.A2(n_303),
.B1(n_250),
.B2(n_222),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_336),
.A2(n_352),
.B1(n_349),
.B2(n_340),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_336),
.A2(n_250),
.B1(n_222),
.B2(n_9),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_393),
.A2(n_394),
.B1(n_362),
.B2(n_338),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_345),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_337),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_7),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_404),
.C(n_418),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_399),
.A2(n_413),
.B1(n_393),
.B2(n_348),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_387),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_401),
.B(n_411),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_360),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_419),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_377),
.C(n_339),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_339),
.C(n_358),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_420),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_380),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_351),
.B1(n_338),
.B2(n_348),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_414),
.Y(n_426)
);

INVx11_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_416),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_343),
.C(n_356),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_357),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_378),
.B(n_361),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g421 ( 
.A(n_374),
.B(n_391),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_421),
.A2(n_391),
.B(n_363),
.Y(n_431)
);

AO22x1_ASAP7_75t_L g422 ( 
.A1(n_421),
.A2(n_374),
.B1(n_413),
.B2(n_382),
.Y(n_422)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_359),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_439),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_342),
.C(n_381),
.Y(n_425)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_361),
.Y(n_429)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_434),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_388),
.B(n_389),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_432),
.A2(n_348),
.B(n_397),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_382),
.C(n_396),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_436),
.C(n_418),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_365),
.Y(n_434)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_435),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_382),
.C(n_390),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_407),
.B(n_394),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_419),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_386),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_428),
.B(n_415),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_448),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_427),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_441),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_454),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_456),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_409),
.C(n_406),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_452),
.B(n_433),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_420),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_424),
.B(n_400),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_441),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_406),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_453),
.A2(n_429),
.B1(n_436),
.B2(n_440),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_461),
.A2(n_465),
.B1(n_468),
.B2(n_430),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_462),
.B(n_466),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_447),
.A2(n_442),
.B1(n_422),
.B2(n_457),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_430),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_435),
.B1(n_432),
.B2(n_422),
.Y(n_464)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_442),
.A2(n_400),
.B1(n_431),
.B2(n_348),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_457),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_467),
.B(n_469),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_451),
.A2(n_348),
.B1(n_438),
.B2(n_410),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_446),
.B(n_449),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_456),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_353),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_471),
.A2(n_354),
.B(n_417),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_458),
.A2(n_452),
.B(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_463),
.A2(n_445),
.B(n_443),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_SL g474 ( 
.A(n_470),
.B(n_443),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_474),
.B(n_479),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_465),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_476),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_481),
.Y(n_489)
);

AOI21xp33_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_460),
.B(n_459),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_483),
.A2(n_475),
.B(n_417),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_471),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_477),
.A2(n_459),
.B(n_464),
.Y(n_490)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_490),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_484),
.B(n_476),
.Y(n_492)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_493),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_485),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_495),
.A2(n_488),
.B(n_489),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_494),
.B(n_487),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_499),
.B(n_500),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_496),
.A2(n_491),
.B(n_486),
.Y(n_500)
);

MAJx2_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_498),
.C(n_8),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_9),
.Y(n_503)
);


endmodule