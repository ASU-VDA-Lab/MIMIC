module fake_jpeg_31985_n_405 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_405);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_68),
.Y(n_120)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_22),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_36),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_85),
.Y(n_124)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_1),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_28),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_84),
.Y(n_104)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_88),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_1),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_32),
.B1(n_38),
.B2(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_92),
.A2(n_96),
.B1(n_105),
.B2(n_111),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_32),
.B1(n_20),
.B2(n_43),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_32),
.B1(n_20),
.B2(n_43),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_110),
.B(n_100),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_20),
.B1(n_43),
.B2(n_26),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_47),
.A2(n_20),
.B1(n_29),
.B2(n_34),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_137),
.B1(n_39),
.B2(n_28),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_34),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_116),
.B(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_46),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_123),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_55),
.B(n_42),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_58),
.B(n_44),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_44),
.C(n_42),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_53),
.B(n_41),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_67),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_60),
.A2(n_39),
.B1(n_26),
.B2(n_19),
.Y(n_137)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_61),
.B1(n_81),
.B2(n_77),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_145),
.A2(n_177),
.B1(n_122),
.B2(n_98),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_19),
.B1(n_26),
.B2(n_56),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_151),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_152),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_149),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_35),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_33),
.B1(n_25),
.B2(n_23),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_33),
.B1(n_25),
.B2(n_23),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_52),
.B1(n_35),
.B2(n_86),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_179),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_84),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_175),
.C(n_108),
.Y(n_187)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_28),
.B(n_37),
.C(n_67),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_170),
.Y(n_185)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_37),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_174),
.Y(n_210)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_99),
.B(n_64),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_66),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_52),
.B1(n_5),
.B2(n_6),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_112),
.B1(n_115),
.B2(n_129),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_121),
.A2(n_130),
.B1(n_119),
.B2(n_93),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_156),
.B1(n_106),
.B2(n_122),
.Y(n_193)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_103),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_186),
.B(n_159),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_211),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_177),
.B1(n_175),
.B2(n_157),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_197),
.B1(n_208),
.B2(n_221),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_127),
.B1(n_90),
.B2(n_126),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_128),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_158),
.C(n_166),
.Y(n_228)
);

XOR2x1_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_119),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_R g232 ( 
.A1(n_206),
.A2(n_207),
.B1(n_215),
.B2(n_146),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_101),
.B1(n_102),
.B2(n_93),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_148),
.A2(n_126),
.B1(n_139),
.B2(n_106),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_102),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_173),
.B1(n_155),
.B2(n_129),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_139),
.B1(n_130),
.B2(n_112),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_161),
.A2(n_138),
.B1(n_97),
.B2(n_115),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_234),
.B1(n_236),
.B2(n_248),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_184),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_227),
.Y(n_259)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_238),
.C(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_149),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_244),
.Y(n_266)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_216),
.B1(n_202),
.B2(n_141),
.Y(n_280)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_157),
.B1(n_175),
.B2(n_169),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_144),
.B1(n_163),
.B2(n_181),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_235),
.A2(n_200),
.B(n_195),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_201),
.B1(n_211),
.B2(n_190),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_179),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_142),
.C(n_143),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_209),
.A2(n_147),
.B1(n_178),
.B2(n_179),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_242),
.B1(n_246),
.B2(n_192),
.Y(n_264)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_209),
.A2(n_160),
.B1(n_152),
.B2(n_151),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_165),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_185),
.B(n_176),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_133),
.B1(n_183),
.B2(n_153),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_186),
.B(n_182),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_168),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_206),
.B(n_154),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_192),
.B(n_207),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_257),
.A2(n_261),
.B(n_263),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_192),
.B(n_212),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_258),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_211),
.C(n_192),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_243),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_192),
.B(n_200),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_275),
.B1(n_277),
.B2(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_198),
.C(n_213),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_247),
.C(n_242),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_236),
.A2(n_215),
.B(n_217),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_271),
.A2(n_229),
.B(n_237),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_213),
.B1(n_198),
.B2(n_189),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_278),
.B1(n_226),
.B2(n_245),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_222),
.A2(n_189),
.B1(n_219),
.B2(n_217),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_219),
.B1(n_172),
.B2(n_214),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_214),
.B1(n_202),
.B2(n_216),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_218),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_239),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_253),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_269),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_250),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_284),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_259),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_238),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_290),
.C(n_291),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_286),
.A2(n_300),
.B(n_305),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_296),
.B1(n_275),
.B2(n_256),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_252),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_292),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_244),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_301),
.C(n_263),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_303),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_276),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_297),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_227),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_227),
.B(n_233),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_248),
.C(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_262),
.A2(n_224),
.B(n_241),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_262),
.A2(n_224),
.B(n_249),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_258),
.B(n_257),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_318),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_264),
.B1(n_273),
.B2(n_258),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_312),
.A2(n_315),
.B1(n_321),
.B2(n_304),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_289),
.A2(n_258),
.B1(n_256),
.B2(n_255),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_285),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_278),
.B1(n_280),
.B2(n_300),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_280),
.B1(n_281),
.B2(n_276),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_282),
.C(n_306),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_294),
.C(n_301),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_325),
.Y(n_339)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_328),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_280),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_290),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_331),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_335),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_291),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_334),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_320),
.A2(n_280),
.B1(n_265),
.B2(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_261),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_342),
.C(n_309),
.Y(n_350)
);

OAI31xp33_ASAP7_75t_L g338 ( 
.A1(n_325),
.A2(n_272),
.A3(n_270),
.B(n_302),
.Y(n_338)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_270),
.B1(n_299),
.B2(n_274),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_340),
.B(n_341),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_323),
.B(n_267),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_315),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_312),
.A2(n_267),
.B1(n_196),
.B2(n_138),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_346),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_196),
.B1(n_97),
.B2(n_8),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_307),
.B(n_4),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_308),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_350),
.B(n_331),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_322),
.Y(n_364)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_356),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_326),
.C(n_311),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_360),
.C(n_335),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_326),
.C(n_328),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_333),
.A2(n_319),
.B(n_322),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_345),
.B(n_346),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_361),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_351),
.A2(n_343),
.B(n_342),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_348),
.B(n_357),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_367),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_334),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_370),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_358),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_341),
.C(n_337),
.Y(n_370)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_371),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_316),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_373),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_313),
.C(n_316),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_376),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_371),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_384),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_349),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_378),
.B(n_382),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_348),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_350),
.Y(n_384)
);

AOI322xp5_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_365),
.A3(n_354),
.B1(n_358),
.B2(n_313),
.C1(n_310),
.C2(n_367),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_385),
.A2(n_386),
.B1(n_379),
.B2(n_383),
.Y(n_393)
);

AOI322xp5_ASAP7_75t_L g386 ( 
.A1(n_383),
.A2(n_310),
.A3(n_370),
.B1(n_366),
.B2(n_352),
.C1(n_7),
.C2(n_9),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_381),
.A2(n_352),
.B(n_8),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_388),
.A2(n_9),
.B(n_387),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_376),
.A2(n_4),
.B(n_8),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_392),
.Y(n_396)
);

NOR2x1_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_8),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_394),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_374),
.C(n_375),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_397),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_385),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_386),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_399),
.B(n_396),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_402),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_399),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_403),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_398),
.Y(n_405)
);


endmodule