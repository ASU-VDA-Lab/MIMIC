module real_jpeg_16702_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_378),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_0),
.B(n_379),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_1),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_2),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_3),
.Y(n_321)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_4),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_5),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_5),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_5),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_5),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_5),
.B(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_5),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_6),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_6),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

AND2x4_ASAP7_75t_SL g196 ( 
.A(n_6),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_8),
.Y(n_379)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

AND2x4_ASAP7_75t_SL g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

NAND2x1p5_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_10),
.B(n_76),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_59),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_11),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_12),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_12),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_12),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_12),
.B(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_160),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_159),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_19),
.B(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.C(n_114),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_20),
.B(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.C(n_78),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_21),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_46),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_22),
.B(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_23),
.A2(n_36),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_31),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_28),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_24),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_98),
.C(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_24),
.A2(n_80),
.B1(n_98),
.B2(n_99),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_24),
.A2(n_80),
.B1(n_180),
.B2(n_181),
.Y(n_251)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_40),
.B(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_32),
.C(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_28),
.A2(n_177),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_28),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_28),
.A2(n_40),
.B1(n_186),
.B2(n_213),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_29),
.Y(n_271)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_31),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_31),
.B(n_32),
.C(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_32),
.A2(n_37),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_32),
.A2(n_37),
.B1(n_236),
.B2(n_240),
.Y(n_235)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_36),
.A2(n_191),
.B(n_196),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_67),
.C(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_38),
.B(n_46),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_40),
.A2(n_192),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_40),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_40),
.A2(n_63),
.B1(n_213),
.B2(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_40),
.B(n_63),
.C(n_249),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_43),
.B(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_43),
.B(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_48),
.A2(n_49),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_48),
.A2(n_49),
.B1(n_98),
.B2(n_99),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_49),
.B(n_52),
.C(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_49),
.B(n_82),
.C(n_119),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_49),
.A2(n_99),
.B(n_170),
.C(n_215),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_56),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_56),
.A2(n_69),
.B1(n_130),
.B2(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_56),
.B(n_153),
.C(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_56),
.A2(n_130),
.B1(n_236),
.B2(n_240),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_101),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_57),
.B(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_60),
.B(n_78),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.C(n_74),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_61),
.A2(n_62),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.C(n_69),
.Y(n_62)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_63),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_63),
.A2(n_69),
.B1(n_153),
.B2(n_264),
.Y(n_338)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_89),
.B1(n_90),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_67),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_67),
.A2(n_134),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_67),
.B(n_75),
.C(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_69),
.A2(n_106),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_69),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_69),
.B(n_113),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_69),
.A2(n_155),
.B(n_156),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_71),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_71),
.B(n_75),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_72),
.B(n_181),
.C(n_295),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_74),
.A2(n_75),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_79),
.C(n_82),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_75),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_75),
.B(n_316),
.C(n_318),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_80),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_84),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_82),
.A2(n_84),
.B1(n_105),
.B2(n_112),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_82),
.B(n_99),
.C(n_106),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_85),
.B(n_114),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_104),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_96),
.B2(n_97),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_87),
.B(n_97),
.C(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_98),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_98),
.B(n_222),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_126),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_100),
.A2(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_100),
.B(n_270),
.Y(n_272)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_106),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_108),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_106),
.A2(n_196),
.B(n_212),
.C(n_215),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_106),
.B(n_196),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_106),
.A2(n_152),
.B1(n_196),
.B2(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_106),
.A2(n_152),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_108),
.Y(n_113)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_152),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_123),
.C(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_131),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_125),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_129),
.B(n_131),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_130),
.B(n_240),
.C(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_134),
.B(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_158),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_148),
.B1(n_149),
.B2(n_157),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_372),
.B(n_376),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_304),
.A3(n_359),
.B1(n_365),
.B2(n_370),
.C(n_371),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_275),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_253),
.B(n_274),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_230),
.B(n_252),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_209),
.B(n_229),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_188),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_188),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.C(n_184),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_170),
.A2(n_174),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_184),
.B1(n_185),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_176),
.A2(n_177),
.B(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_180),
.A2(n_181),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_199),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_200),
.C(n_208),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_221),
.B(n_223),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_196),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_207),
.B2(n_208),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_204),
.A2(n_249),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_219),
.B(n_228),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_216),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_225),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_224),
.B(n_227),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_232),
.Y(n_252)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_241),
.C(n_242),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

OR2x6_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_247),
.C(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_255),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_266),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_258),
.C(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_262),
.C(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_273),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_269),
.C(n_273),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_276),
.B(n_277),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_290),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_278),
.B(n_291),
.C(n_303),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_285),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_284),
.C(n_288),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_303),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_301),
.C(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_346),
.Y(n_304)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_339),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_306),
.B(n_339),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.C(n_323),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_324),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_312),
.A2(n_314),
.B1(n_315),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_331),
.C(n_332),
.Y(n_340)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.C(n_337),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_333),
.A2(n_334),
.B1(n_336),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_342),
.C(n_344),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

AOI31xp67_ASAP7_75t_L g365 ( 
.A1(n_346),
.A2(n_360),
.A3(n_366),
.B(n_369),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_349),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.C(n_355),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_350),
.A2(n_351),
.B1(n_355),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_355),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_361),
.B(n_364),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

AND2x4_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);


endmodule