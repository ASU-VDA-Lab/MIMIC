module fake_jpeg_1021_n_193 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_29),
.B1(n_23),
.B2(n_19),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_70),
.B1(n_26),
.B2(n_2),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_23),
.B1(n_51),
.B2(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_20),
.B1(n_26),
.B2(n_21),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_32),
.B1(n_25),
.B2(n_22),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_22),
.B1(n_28),
.B2(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_15),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_17),
.B(n_2),
.C(n_4),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_19),
.B1(n_33),
.B2(n_28),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_22),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_26),
.C(n_4),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_88),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_20),
.B1(n_15),
.B2(n_17),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_71),
.B1(n_60),
.B2(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_96),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_1),
.Y(n_93)
);

NAND2x1_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_68),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_117),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_71),
.C(n_52),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_84),
.C(n_92),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_98),
.B1(n_99),
.B2(n_78),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_72),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_102),
.A3(n_101),
.B1(n_86),
.B2(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_135),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_89),
.B(n_79),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_130),
.B(n_108),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_131),
.C(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_87),
.C(n_52),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_65),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_139),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_65),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_111),
.B1(n_123),
.B2(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_143),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_90),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_123),
.C(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_149),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_141),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_125),
.B1(n_112),
.B2(n_107),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_151),
.B(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_126),
.B1(n_138),
.B2(n_134),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_108),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_143),
.B(n_120),
.C(n_105),
.D(n_124),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_131),
.C(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_148),
.C(n_154),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_107),
.B1(n_142),
.B2(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_164),
.B1(n_153),
.B2(n_155),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_165),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_116),
.B(n_106),
.C(n_117),
.D(n_11),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_106),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_171),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_144),
.B(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_170),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_148),
.C(n_149),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_179),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_172),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_159),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_167),
.B(n_175),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_175),
.C(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_185),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_181),
.B(n_178),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_145),
.C(n_116),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_181),
.B1(n_9),
.B2(n_12),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_186),
.B(n_90),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_189),
.C(n_7),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_7),
.Y(n_193)
);


endmodule