module real_jpeg_30349_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_605;
wire n_216;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_667;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_636;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_0),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_0),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_1),
.A2(n_60),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_1),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_1),
.A2(n_360),
.B1(n_435),
.B2(n_440),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_1),
.A2(n_118),
.B1(n_360),
.B2(n_584),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_1),
.A2(n_360),
.B1(n_637),
.B2(n_638),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_2),
.A2(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_2),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_2),
.A2(n_384),
.B1(n_478),
.B2(n_481),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_2),
.A2(n_384),
.B1(n_584),
.B2(n_618),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_2),
.A2(n_384),
.B1(n_626),
.B2(n_627),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_4),
.A2(n_309),
.B1(n_313),
.B2(n_314),
.Y(n_308)
);

INVx2_ASAP7_75t_R g313 ( 
.A(n_4),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_4),
.A2(n_313),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_4),
.A2(n_313),
.B1(n_536),
.B2(n_539),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_4),
.A2(n_313),
.B1(n_601),
.B2(n_605),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_138),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_5),
.A2(n_214),
.B1(n_321),
.B2(n_325),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_5),
.A2(n_365),
.B(n_369),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_5),
.A2(n_214),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_6),
.A2(n_355),
.B(n_357),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_6),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_6),
.B(n_453),
.Y(n_452)
);

OAI32xp33_ASAP7_75t_L g544 ( 
.A1(n_6),
.A2(n_147),
.A3(n_545),
.B1(n_548),
.B2(n_554),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_6),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_6),
.B(n_177),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_6),
.A2(n_290),
.B1(n_636),
.B2(n_644),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_6),
.A2(n_555),
.B1(n_662),
.B2(n_667),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_7),
.A2(n_125),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx2_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_7),
.A2(n_267),
.B1(n_372),
.B2(n_375),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_7),
.A2(n_267),
.B1(n_276),
.B2(n_470),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_7),
.A2(n_267),
.B1(n_562),
.B2(n_566),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_10),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_11),
.Y(n_569)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_13),
.A2(n_74),
.B1(n_77),
.B2(n_84),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_13),
.A2(n_84),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_13),
.A2(n_84),
.B1(n_180),
.B2(n_184),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_13),
.A2(n_84),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_14),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_14),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_14),
.A2(n_127),
.B1(n_182),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_14),
.A2(n_127),
.B1(n_301),
.B2(n_305),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_14),
.A2(n_127),
.B1(n_415),
.B2(n_418),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_15),
.B(n_23),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_16),
.A2(n_58),
.B1(n_65),
.B2(n_70),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_16),
.A2(n_70),
.B1(n_167),
.B2(n_173),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_16),
.A2(n_70),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_16),
.A2(n_70),
.B1(n_245),
.B2(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_17),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_17),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_18),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_18),
.Y(n_159)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_18),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_19),
.A2(n_134),
.B1(n_137),
.B2(n_143),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_19),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_19),
.A2(n_143),
.B1(n_182),
.B2(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_19),
.A2(n_143),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_19),
.A2(n_143),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_693),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_196),
.B(n_692),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_29),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_23),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_SL g693 ( 
.A(n_29),
.B(n_197),
.C(n_694),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_195),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_85),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_32),
.B(n_85),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_57),
.B1(n_71),
.B2(n_73),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_33),
.A2(n_123),
.B1(n_131),
.B2(n_133),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_33),
.A2(n_131),
.B1(n_308),
.B2(n_316),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_33),
.A2(n_71),
.B1(n_354),
.B2(n_359),
.Y(n_353)
);

OAI22x1_ASAP7_75t_L g500 ( 
.A1(n_33),
.A2(n_71),
.B1(n_308),
.B2(n_477),
.Y(n_500)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_34),
.B(n_213),
.Y(n_212)
);

NAND2x1p5_ASAP7_75t_L g265 ( 
.A(n_34),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_34),
.A2(n_210),
.B1(n_476),
.B2(n_483),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_37),
.Y(n_327)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_38),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_38),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_38),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_38),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_41),
.Y(n_399)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_41),
.Y(n_408)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_43),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_43),
.Y(n_388)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_48),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_49),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_49),
.Y(n_480)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_57),
.A2(n_71),
.B1(n_133),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_62),
.Y(n_269)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_63),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_71),
.Y(n_453)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g430 ( 
.A1(n_78),
.A2(n_395),
.A3(n_400),
.B1(n_404),
.B2(n_412),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_82),
.Y(n_356)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_188),
.C(n_190),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_86),
.A2(n_87),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_122),
.C(n_144),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_88),
.A2(n_145),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_88),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_88),
.A2(n_207),
.B1(n_218),
.B2(n_336),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_100),
.B(n_113),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_89),
.A2(n_100),
.B1(n_250),
.B2(n_256),
.Y(n_249)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_89),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_89),
.A2(n_100),
.B1(n_250),
.B2(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_89),
.A2(n_100),
.B1(n_364),
.B2(n_371),
.Y(n_363)
);

OAI22x1_ASAP7_75t_SL g462 ( 
.A1(n_89),
.A2(n_100),
.B1(n_300),
.B2(n_364),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_89),
.A2(n_100),
.B1(n_371),
.B2(n_534),
.Y(n_533)
);

OAI22x1_ASAP7_75t_L g615 ( 
.A1(n_89),
.A2(n_100),
.B1(n_616),
.B2(n_617),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_89),
.B(n_555),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO21x2_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_101),
.B(n_108),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_91),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_91)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_92),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_93),
.Y(n_241)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_93),
.Y(n_248)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_93),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_93),
.Y(n_604)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_93),
.Y(n_608)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_96),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_97),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_101),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_107),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_107),
.Y(n_541)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_107),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_108),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_113),
.Y(n_284)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_120),
.Y(n_258)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_120),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_121),
.Y(n_255)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_121),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_121),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_122),
.B(n_205),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_123),
.A2(n_209),
.B(n_212),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g394 ( 
.A1(n_138),
.A2(n_395),
.A3(n_400),
.B1(n_404),
.B2(n_412),
.Y(n_394)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_142),
.Y(n_312)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_142),
.Y(n_315)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_142),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_166),
.B1(n_176),
.B2(n_179),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_146),
.A2(n_166),
.B1(n_176),
.B2(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_146),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_146),
.A2(n_176),
.B1(n_385),
.B2(n_469),
.Y(n_468)
);

OAI22x1_ASAP7_75t_L g498 ( 
.A1(n_146),
.A2(n_176),
.B1(n_320),
.B2(n_469),
.Y(n_498)
);

AO21x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_153),
.B(n_160),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_148),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_149),
.Y(n_411)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_159),
.Y(n_383)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_160)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_162),
.Y(n_368)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_162),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_172),
.Y(n_392)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_176),
.A2(n_379),
.B1(n_380),
.B2(n_385),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_176),
.A2(n_192),
.B1(n_380),
.B2(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_191),
.B(n_194),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_177),
.A2(n_193),
.B1(n_220),
.B2(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_177),
.A2(n_275),
.B1(n_319),
.B2(n_328),
.Y(n_318)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_178),
.A2(n_379),
.B1(n_434),
.B2(n_661),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_183),
.Y(n_440)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_190),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_224),
.B(n_687),
.Y(n_197)
);

OA21x2_ASAP7_75t_SL g687 ( 
.A1(n_198),
.A2(n_688),
.B(n_691),
.Y(n_687)
);

NOR2x1_ASAP7_75t_R g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_199),
.B(n_202),
.Y(n_691)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.C(n_217),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_204),
.B(n_208),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_208),
.C(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_208),
.A2(n_286),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_208),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_208),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_209),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_214),
.B(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_217),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_218),
.Y(n_336)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_223),
.Y(n_403)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_223),
.Y(n_474)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_223),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_347),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_341),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_329),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_227),
.B(n_329),
.Y(n_689)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_271),
.C(n_287),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_229),
.B(n_504),
.Y(n_503)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_262),
.Y(n_229)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_230),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_249),
.Y(n_230)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_231),
.A2(n_339),
.B(n_340),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_231),
.B(n_249),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_235),
.B(n_242),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g461 ( 
.A(n_234),
.Y(n_461)
);

INVx4_ASAP7_75t_SL g644 ( 
.A(n_234),
.Y(n_644)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_235),
.A2(n_414),
.B1(n_421),
.B2(n_423),
.Y(n_413)
);

AO22x1_ASAP7_75t_L g560 ( 
.A1(n_235),
.A2(n_421),
.B1(n_447),
.B2(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_236),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_236),
.A2(n_291),
.B1(n_424),
.B2(n_459),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_236),
.A2(n_625),
.B1(n_636),
.B2(n_639),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_241),
.Y(n_417)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_241),
.Y(n_448)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_290),
.B1(n_291),
.B2(n_295),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_248),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_255),
.Y(n_370)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_255),
.Y(n_618)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_272),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_286),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_278),
.Y(n_286)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_279),
.A2(n_577),
.B1(n_582),
.B2(n_583),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_279),
.A2(n_285),
.B1(n_535),
.B2(n_671),
.Y(n_670)
);

OA21x2_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B(n_282),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g586 ( 
.A1(n_281),
.A2(n_587),
.B(n_590),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_282),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_286),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_287),
.B(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_306),
.C(n_317),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_288),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_299),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_289),
.B(n_299),
.Y(n_515)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_293),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_293),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx6_ASAP7_75t_L g589 ( 
.A(n_294),
.Y(n_589)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_294),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_294),
.Y(n_651)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx4f_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_304),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g491 ( 
.A1(n_307),
.A2(n_317),
.B1(n_318),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_307),
.Y(n_492)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_338),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_334),
.B1(n_335),
.B2(n_337),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_338),
.C(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_342),
.A2(n_689),
.B(n_690),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_343),
.B(n_345),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_525),
.B(n_682),
.Y(n_347)
);

NAND4xp25_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_487),
.C(n_505),
.D(n_518),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_454),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_350),
.B(n_454),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_393),
.C(n_432),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_351),
.B(n_528),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_362),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_353),
.B(n_363),
.C(n_378),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_359),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_378),
.Y(n_362)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_392),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_393),
.B(n_432),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_413),
.B1(n_429),
.B2(n_431),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_431),
.Y(n_486)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_409),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

AO22x1_ASAP7_75t_SL g441 ( 
.A1(n_414),
.A2(n_442),
.B1(n_446),
.B2(n_447),
.Y(n_441)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_441),
.C(n_451),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_433),
.B(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_441),
.B(n_452),
.Y(n_531)
);

INVx3_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

INVx8_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_445),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_445),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_445),
.Y(n_648)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_446),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_446),
.A2(n_460),
.B1(n_624),
.B2(n_631),
.Y(n_623)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_465),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_457),
.B1(n_463),
.B2(n_464),
.Y(n_455)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_456),
.Y(n_463)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_462),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_462),
.Y(n_501)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_464),
.B(n_466),
.C(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_486),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_475),
.B1(n_484),
.B2(n_485),
.Y(n_467)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_475),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_475),
.Y(n_513)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_484),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g512 ( 
.A(n_486),
.Y(n_512)
);

A2O1A1O1Ixp25_ASAP7_75t_L g682 ( 
.A1(n_487),
.A2(n_505),
.B(n_683),
.C(n_685),
.D(n_686),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_502),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_488),
.B(n_502),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_493),
.C(n_495),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_517),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_496),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

MAJx2_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_499),
.C(n_501),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_497),
.A2(n_498),
.B1(n_500),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_500),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_516),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_506),
.B(n_516),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_511),
.C(n_515),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_524),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.C(n_514),
.Y(n_511)
);

MAJx2_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_513),
.C(n_514),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_515),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_519),
.B(n_521),
.C(n_684),
.Y(n_683)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_570),
.B(n_681),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_529),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_SL g681 ( 
.A(n_527),
.B(n_529),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_532),
.C(n_542),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g676 ( 
.A(n_530),
.B(n_677),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_532),
.A2(n_543),
.B(n_678),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_533),
.B(n_543),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_541),
.Y(n_579)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_560),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_SL g658 ( 
.A(n_544),
.B(n_560),
.Y(n_658)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_551),
.Y(n_581)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_556),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_555),
.A2(n_578),
.B(n_580),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_555),
.B(n_581),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_555),
.B(n_647),
.Y(n_646)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_571),
.A2(n_675),
.B(n_680),
.Y(n_570)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_572),
.A2(n_655),
.B(n_674),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_573),
.A2(n_621),
.B(n_654),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_597),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_574),
.B(n_597),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_575),
.B(n_585),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_575),
.A2(n_576),
.B1(n_585),
.B2(n_586),
.Y(n_632)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_580),
.A2(n_591),
.B(n_594),
.Y(n_590)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_583),
.Y(n_616)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_592),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_598),
.B(n_613),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_598),
.B(n_615),
.C(n_619),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_599),
.A2(n_600),
.B1(n_609),
.B2(n_612),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_600),
.Y(n_631)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_603),
.Y(n_626)
);

INVx6_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_614),
.A2(n_615),
.B1(n_619),
.B2(n_620),
.Y(n_613)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_614),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_615),
.Y(n_620)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_617),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_622),
.A2(n_633),
.B(n_653),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_632),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_623),
.B(n_632),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_626),
.Y(n_638)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_634),
.A2(n_642),
.B(n_652),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_635),
.B(n_641),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_635),
.B(n_641),
.Y(n_652)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_643),
.B(n_645),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_R g645 ( 
.A(n_646),
.B(n_649),
.Y(n_645)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_656),
.B(n_657),
.Y(n_655)
);

NOR2x1_ASAP7_75t_SL g674 ( 
.A(n_656),
.B(n_657),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_658),
.B(n_659),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_658),
.B(n_670),
.C(n_673),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_660),
.A2(n_670),
.B1(n_672),
.B2(n_673),
.Y(n_659)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_660),
.Y(n_673)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_665),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_668),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_669),
.Y(n_668)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_670),
.Y(n_672)
);

NOR2x1_ASAP7_75t_SL g675 ( 
.A(n_676),
.B(n_679),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_676),
.B(n_679),
.Y(n_680)
);


endmodule