module fake_jpeg_22301_n_228 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_23),
.Y(n_49)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_29),
.B1(n_21),
.B2(n_22),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_25),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_25),
.B(n_18),
.C(n_36),
.D(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_22),
.B1(n_23),
.B2(n_21),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_26),
.C(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_30),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_36),
.B1(n_44),
.B2(n_37),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_94),
.B1(n_72),
.B2(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_96),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_33),
.B1(n_17),
.B2(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_10),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_118),
.B1(n_100),
.B2(n_83),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_63),
.C(n_51),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_114),
.C(n_73),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_54),
.B1(n_24),
.B2(n_68),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_62),
.B1(n_59),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_97),
.B1(n_81),
.B2(n_86),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_18),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_79),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_121),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_18),
.B1(n_62),
.B2(n_37),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_18),
.B(n_19),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_122),
.B(n_19),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_18),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_3),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_131),
.B1(n_138),
.B2(n_145),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_75),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_136),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_73),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_104),
.B1(n_107),
.B2(n_76),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_74),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_124),
.B(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_47),
.B1(n_44),
.B2(n_19),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_35),
.B1(n_47),
.B2(n_15),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_104),
.B(n_102),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_76),
.B1(n_35),
.B2(n_70),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_114),
.C(n_106),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_151),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_113),
.C(n_119),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_157),
.B1(n_130),
.B2(n_146),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_165),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_105),
.B(n_121),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_168),
.B(n_148),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_35),
.B(n_64),
.C(n_7),
.D(n_8),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_35),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_3),
.B(n_6),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_183),
.B1(n_185),
.B2(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_145),
.A3(n_138),
.B1(n_135),
.B2(n_126),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_167),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_153),
.C(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_127),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_139),
.B(n_129),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_170),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_6),
.B(n_7),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_154),
.C(n_151),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_187),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_155),
.C(n_176),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_189),
.C(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_152),
.C(n_157),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_204),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_150),
.C(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_173),
.B(n_171),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_10),
.B(n_12),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_160),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_196),
.B1(n_179),
.B2(n_160),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_179),
.B1(n_186),
.B2(n_185),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_158),
.B1(n_165),
.B2(n_99),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_206),
.B(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_200),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_212),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_199),
.C(n_12),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_13),
.B(n_7),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_209),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_219),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_6),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_215),
.B(n_13),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_225),
.B1(n_8),
.B2(n_122),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_220),
.B1(n_99),
.B2(n_8),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);


endmodule