module fake_ibex_1864_n_992 (n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_992);

input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_992;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_510;
wire n_193;
wire n_418;
wire n_845;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_959;
wire n_336;
wire n_930;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_158;
wire n_859;
wire n_470;
wire n_276;
wire n_339;
wire n_259;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_167;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_152;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_299;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_354;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_564;
wire n_506;
wire n_562;
wire n_444;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_947;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_921;
wire n_912;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_159;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_40),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_58),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_37),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_10),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_52),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_73),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_53),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_141),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_25),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_12),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_50),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_22),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_36),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_68),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_34),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_28),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_47),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_38),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_55),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_7),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_98),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_72),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_21),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_127),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_146),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_29),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_67),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_79),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_65),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_80),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_96),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_25),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_88),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_48),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_69),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_24),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_15),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_149),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_85),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_109),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_90),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_105),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_32),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_22),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_43),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_0),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_122),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_23),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_41),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_106),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_35),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_170),
.B(n_1),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_160),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_1),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_2),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_27),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_188),
.B(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_202),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_189),
.B(n_5),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_197),
.B(n_8),
.Y(n_268)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_171),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_168),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_184),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_157),
.B(n_8),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_193),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

NAND2x1p5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_84),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_237),
.B(n_83),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_156),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_10),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_156),
.B(n_11),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_215),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_161),
.B(n_91),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_164),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_172),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_12),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_174),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_174),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_176),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_176),
.Y(n_306)
);

AND3x2_ASAP7_75t_L g307 ( 
.A(n_164),
.B(n_13),
.C(n_15),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_217),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_217),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_229),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_165),
.B(n_13),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_165),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_167),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_151),
.Y(n_316)
);

BUFx8_ASAP7_75t_L g317 ( 
.A(n_154),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_155),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_181),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_243),
.B(n_16),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_159),
.B(n_17),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_162),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_243),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_213),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_187),
.B(n_17),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_180),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_183),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_200),
.Y(n_330)
);

BUFx8_ASAP7_75t_L g331 ( 
.A(n_185),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_186),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_190),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_205),
.B(n_18),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_210),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_194),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_211),
.B(n_19),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_195),
.Y(n_339)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_196),
.B(n_94),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_262),
.B(n_218),
.Y(n_343)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_276),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_253),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

OR2x6_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_225),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_324),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_284),
.B(n_198),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_254),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_264),
.B(n_232),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_291),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_283),
.B(n_178),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_340),
.B(n_199),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_253),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_254),
.B(n_207),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_280),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_212),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_254),
.A2(n_203),
.B1(n_177),
.B2(n_191),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_285),
.B(n_220),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_253),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_224),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_272),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_272),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_272),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_284),
.B(n_251),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_272),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_323),
.B(n_152),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_272),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_291),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_265),
.Y(n_392)
);

BUFx4f_ASAP7_75t_L g393 ( 
.A(n_286),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_300),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_337),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_252),
.B(n_226),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_300),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_252),
.B(n_227),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_340),
.B(n_228),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_304),
.B(n_233),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_294),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_251),
.B(n_235),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_294),
.Y(n_403)
);

INVx4_ASAP7_75t_SL g404 ( 
.A(n_308),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_284),
.B(n_238),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_266),
.B(n_240),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_255),
.B(n_166),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_279),
.Y(n_412)
);

NOR2x1p5_ASAP7_75t_L g413 ( 
.A(n_326),
.B(n_152),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_296),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_296),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_308),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_319),
.B(n_175),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_250),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_308),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_250),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_260),
.B(n_158),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_256),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_308),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_266),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_330),
.B(n_175),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_260),
.B(n_179),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_256),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g432 ( 
.A1(n_263),
.A2(n_208),
.B1(n_206),
.B2(n_182),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_267),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_267),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_286),
.B(n_150),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_270),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_270),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_287),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_287),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_288),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_281),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_271),
.B(n_219),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_L g443 ( 
.A(n_271),
.B(n_249),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_273),
.B(n_173),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_288),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_257),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_257),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_273),
.B(n_249),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_274),
.B(n_192),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_274),
.B(n_248),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_257),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_275),
.B(n_248),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_277),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_317),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_316),
.B(n_203),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_289),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_298),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_258),
.B(n_279),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_275),
.B(n_222),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_313),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_335),
.B(n_222),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_325),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_392),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_454),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_392),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_454),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_356),
.B(n_258),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_356),
.B(n_430),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_437),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_278),
.Y(n_473)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_368),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_387),
.B(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_365),
.A2(n_302),
.B1(n_268),
.B2(n_317),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_383),
.A2(n_405),
.B(n_357),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_428),
.B(n_302),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_378),
.B(n_352),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_429),
.B(n_461),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_437),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_414),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_365),
.A2(n_399),
.B1(n_393),
.B2(n_435),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_419),
.B(n_338),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_416),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_278),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_341),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_368),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_282),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_312),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_368),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_312),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_349),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_349),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_341),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_353),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_449),
.B(n_316),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_399),
.A2(n_268),
.B1(n_332),
.B2(n_339),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_438),
.Y(n_501)
);

AND2x6_ASAP7_75t_SL g502 ( 
.A(n_352),
.B(n_320),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_378),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_386),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_450),
.B(n_452),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_353),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_368),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_352),
.B(n_318),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_378),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_376),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_359),
.B(n_317),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_343),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_367),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_406),
.A2(n_339),
.B1(n_318),
.B2(n_322),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_367),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_377),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_377),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_346),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_411),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_438),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_439),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_322),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_452),
.B(n_332),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_396),
.B(n_331),
.Y(n_528)
);

AND2x4_ASAP7_75t_SL g529 ( 
.A(n_411),
.B(n_150),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_347),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_354),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_368),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_343),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_355),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_376),
.B(n_333),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_432),
.B(n_327),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_406),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_359),
.B(n_374),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_459),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_406),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_361),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_371),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_453),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_393),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_361),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_455),
.B(n_333),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_424),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_415),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_351),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_431),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_396),
.B(n_331),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_415),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_351),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_455),
.B(n_301),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_374),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_398),
.B(n_331),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_432),
.B(n_334),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_410),
.B(n_329),
.Y(n_566)
);

AOI221x1_ASAP7_75t_L g567 ( 
.A1(n_402),
.A2(n_290),
.B1(n_261),
.B2(n_321),
.C(n_315),
.Y(n_567)
);

NOR2x1_ASAP7_75t_L g568 ( 
.A(n_413),
.B(n_177),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_385),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_364),
.A2(n_191),
.B1(n_329),
.B2(n_336),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_436),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_445),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_406),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_463),
.B(n_364),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_467),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_463),
.A2(n_492),
.B1(n_509),
.B2(n_469),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_501),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_465),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_540),
.A2(n_564),
.B1(n_521),
.B2(n_509),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_466),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_472),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_506),
.B(n_382),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_497),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

O2A1O1Ixp33_ASAP7_75t_L g587 ( 
.A1(n_551),
.A2(n_560),
.B(n_524),
.C(n_525),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_481),
.A2(n_410),
.B1(n_443),
.B2(n_383),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_482),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_505),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_SL g591 ( 
.A(n_477),
.B(n_231),
.C(n_357),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_553),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_528),
.B(n_398),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_480),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_507),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_480),
.B(n_553),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_573),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_540),
.A2(n_231),
.B1(n_391),
.B2(n_395),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_515),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_489),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_480),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_516),
.A2(n_372),
.B1(n_373),
.B2(n_402),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_503),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_490),
.B(n_474),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_506),
.B(n_456),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_517),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_522),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_557),
.B(n_448),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_543),
.B(n_462),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_535),
.Y(n_616)
);

BUFx2_ASAP7_75t_SL g617 ( 
.A(n_489),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_562),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_540),
.A2(n_443),
.B1(n_405),
.B2(n_448),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_493),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_521),
.B(n_425),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_518),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_500),
.B(n_444),
.C(n_425),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_564),
.A2(n_460),
.B1(n_457),
.B2(n_360),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_519),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_493),
.B(n_444),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_479),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_514),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_370),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_537),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_510),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_475),
.B(n_370),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g634 ( 
.A1(n_564),
.A2(n_277),
.B1(n_400),
.B2(n_301),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_570),
.B(n_400),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_523),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_545),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_526),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_476),
.Y(n_640)
);

NOR2x1_ASAP7_75t_SL g641 ( 
.A(n_493),
.B(n_342),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_563),
.B(n_345),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_490),
.A2(n_543),
.B1(n_548),
.B2(n_504),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_464),
.Y(n_644)
);

AOI222xp33_ASAP7_75t_L g645 ( 
.A1(n_484),
.A2(n_277),
.B1(n_336),
.B2(n_305),
.C1(n_306),
.C2(n_309),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_548),
.B(n_369),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_493),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_539),
.B(n_434),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_520),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_524),
.A2(n_315),
.B1(n_305),
.B2(n_306),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_483),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_573),
.B(n_508),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_512),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_479),
.A2(n_303),
.B1(n_309),
.B2(n_297),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_471),
.B(n_485),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_468),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_471),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_502),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_525),
.A2(n_259),
.B(n_394),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_551),
.B(n_303),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_473),
.B(n_307),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_560),
.A2(n_201),
.B1(n_234),
.B2(n_239),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_508),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_SL g664 ( 
.A(n_508),
.B(n_344),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_530),
.Y(n_665)
);

AO21x1_ASAP7_75t_L g666 ( 
.A1(n_478),
.A2(n_259),
.B(n_363),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_473),
.B(n_427),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_566),
.B(n_344),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_549),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_542),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_499),
.B(n_427),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_474),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_486),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_531),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_487),
.B(n_422),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_508),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_538),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_536),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_587),
.A2(n_484),
.B1(n_541),
.B2(n_561),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_575),
.Y(n_681)
);

OAI222xp33_ASAP7_75t_L g682 ( 
.A1(n_602),
.A2(n_546),
.B1(n_568),
.B2(n_513),
.C1(n_544),
.C2(n_491),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_L g683 ( 
.A1(n_576),
.A2(n_494),
.B1(n_491),
.B2(n_487),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_609),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_655),
.B(n_494),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g686 ( 
.A1(n_666),
.A2(n_567),
.B(n_478),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_609),
.A2(n_499),
.B1(n_536),
.B2(n_572),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_627),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_614),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_587),
.A2(n_571),
.B1(n_552),
.B2(n_565),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_614),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_584),
.A2(n_536),
.B1(n_555),
.B2(n_556),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_615),
.A2(n_244),
.B1(n_532),
.B2(n_547),
.Y(n_693)
);

AOI221xp5_ASAP7_75t_L g694 ( 
.A1(n_597),
.A2(n_533),
.B1(n_534),
.B2(n_422),
.C(n_385),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_592),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_616),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_635),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_579),
.A2(n_584),
.B1(n_634),
.B2(n_660),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_634),
.A2(n_397),
.B1(n_292),
.B2(n_295),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_640),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_598),
.A2(n_474),
.B1(n_344),
.B2(n_350),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_600),
.B(n_495),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_586),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_657),
.B(n_495),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_651),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_SL g706 ( 
.A1(n_660),
.A2(n_381),
.B(n_380),
.C(n_366),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_612),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_673),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_591),
.A2(n_397),
.B1(n_559),
.B2(n_554),
.Y(n_709)
);

INVx6_ASAP7_75t_L g710 ( 
.A(n_598),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_643),
.B(n_19),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_633),
.B(n_344),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_659),
.A2(n_569),
.B(n_496),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_648),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_600),
.B(n_495),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_637),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_574),
.B(n_496),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_667),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_630),
.A2(n_281),
.B1(n_292),
.B2(n_295),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_639),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_596),
.A2(n_605),
.B1(n_621),
.B2(n_630),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_592),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_582),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_636),
.B(n_20),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_585),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_618),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_591),
.A2(n_496),
.B1(n_350),
.B2(n_366),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_667),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_662),
.A2(n_281),
.B1(n_292),
.B2(n_295),
.C(n_299),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_608),
.B(n_350),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_350),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_602),
.A2(n_628),
.B1(n_645),
.B2(n_613),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_618),
.B(n_20),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_630),
.A2(n_299),
.B1(n_381),
.B2(n_380),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_675),
.Y(n_736)
);

INVx6_ASAP7_75t_L g737 ( 
.A(n_621),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_631),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_588),
.B(n_21),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_645),
.B(n_23),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_644),
.B(n_299),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_621),
.B(n_404),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_661),
.B(n_348),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_601),
.B(n_404),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_624),
.A2(n_390),
.B1(n_358),
.B2(n_362),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_607),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_675),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_631),
.B(n_348),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_SL g749 ( 
.A1(n_658),
.A2(n_348),
.B1(n_388),
.B2(n_375),
.Y(n_749)
);

NAND2x1_ASAP7_75t_L g750 ( 
.A(n_664),
.B(n_348),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_623),
.A2(n_375),
.B1(n_379),
.B2(n_384),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_659),
.A2(n_389),
.B(n_423),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_646),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_661),
.A2(n_375),
.B1(n_379),
.B2(n_384),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_662),
.A2(n_408),
.B(n_421),
.C(n_407),
.Y(n_755)
);

BUFx2_ASAP7_75t_R g756 ( 
.A(n_632),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_646),
.A2(n_375),
.B1(n_388),
.B2(n_379),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_595),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_668),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_599),
.Y(n_760)
);

AOI21x1_ASAP7_75t_L g761 ( 
.A1(n_650),
.A2(n_606),
.B(n_626),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_671),
.A2(n_379),
.B1(n_384),
.B2(n_388),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_606),
.A2(n_384),
.B1(n_388),
.B2(n_423),
.Y(n_763)
);

BUFx12f_ASAP7_75t_L g764 ( 
.A(n_652),
.Y(n_764)
);

AOI221xp5_ASAP7_75t_L g765 ( 
.A1(n_650),
.A2(n_409),
.B1(n_441),
.B2(n_417),
.C(n_418),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_638),
.B(n_404),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_603),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_670),
.A2(n_441),
.B(n_418),
.C(n_417),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_611),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_629),
.A2(n_418),
.B1(n_417),
.B2(n_441),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_622),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_625),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_653),
.B(n_441),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_649),
.Y(n_774)
);

CKINVDCx6p67_ASAP7_75t_R g775 ( 
.A(n_669),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_617),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_619),
.A2(n_642),
.B1(n_670),
.B2(n_583),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_665),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_593),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_654),
.B(n_418),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_577),
.A2(n_417),
.B1(n_33),
.B2(n_39),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_592),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_674),
.Y(n_783)
);

AO22x1_ASAP7_75t_L g784 ( 
.A1(n_672),
.A2(n_31),
.B1(n_42),
.B2(n_44),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_677),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_577),
.A2(n_46),
.B1(n_49),
.B2(n_54),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_601),
.B(n_57),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_583),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_578),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_580),
.A2(n_64),
.B1(n_71),
.B2(n_74),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_581),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_589),
.A2(n_77),
.B1(n_81),
.B2(n_87),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_684),
.B(n_593),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_688),
.Y(n_794)
);

AOI221xp5_ASAP7_75t_L g795 ( 
.A1(n_683),
.A2(n_590),
.B1(n_610),
.B2(n_676),
.C(n_663),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_698),
.A2(n_663),
.B1(n_678),
.B2(n_676),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_696),
.B(n_727),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_706),
.A2(n_641),
.B(n_672),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_689),
.A2(n_652),
.B1(n_678),
.B2(n_679),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_691),
.A2(n_679),
.B1(n_647),
.B2(n_620),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_697),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_753),
.B(n_679),
.Y(n_802)
);

OA21x2_ASAP7_75t_L g803 ( 
.A1(n_752),
.A2(n_92),
.B(n_93),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_764),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_685),
.B(n_647),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_696),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_686),
.A2(n_95),
.B(n_97),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_724),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_733),
.A2(n_647),
.B1(n_620),
.B2(n_604),
.Y(n_809)
);

AOI222xp33_ASAP7_75t_L g810 ( 
.A1(n_682),
.A2(n_620),
.B1(n_604),
.B2(n_594),
.C1(n_102),
.C2(n_103),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_700),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_722),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_698),
.A2(n_604),
.B1(n_594),
.B2(n_101),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_725),
.B(n_594),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_SL g815 ( 
.A1(n_737),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_815)
);

AOI221xp5_ASAP7_75t_L g816 ( 
.A1(n_714),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.C(n_115),
.Y(n_816)
);

AO21x2_ASAP7_75t_L g817 ( 
.A1(n_763),
.A2(n_118),
.B(n_119),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_726),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_718),
.A2(n_123),
.B1(n_129),
.B2(n_130),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_705),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_760),
.Y(n_821)
);

INVx8_ASAP7_75t_L g822 ( 
.A(n_731),
.Y(n_822)
);

OAI21xp33_ASAP7_75t_L g823 ( 
.A1(n_734),
.A2(n_132),
.B(n_133),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_740),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_771),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_713),
.A2(n_143),
.B(n_144),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_738),
.B(n_772),
.Y(n_827)
);

AO21x2_ASAP7_75t_L g828 ( 
.A1(n_761),
.A2(n_757),
.B(n_690),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_708),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_SL g830 ( 
.A1(n_737),
.A2(n_711),
.B1(n_710),
.B2(n_776),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_729),
.A2(n_747),
.B1(n_736),
.B2(n_680),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_680),
.A2(n_690),
.B1(n_739),
.B2(n_759),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_742),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_695),
.B(n_723),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_758),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_693),
.B(n_712),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_L g837 ( 
.A1(n_721),
.A2(n_777),
.B1(n_728),
.B2(n_709),
.C(n_681),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_768),
.A2(n_751),
.B(n_750),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_767),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_769),
.B(n_746),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_759),
.A2(n_707),
.B1(n_720),
.B2(n_716),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_710),
.B(n_709),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_776),
.A2(n_719),
.B1(n_792),
.B2(n_687),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_775),
.A2(n_703),
.B1(n_742),
.B2(n_694),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_699),
.A2(n_692),
.B(n_719),
.C(n_735),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_699),
.A2(n_785),
.B1(n_704),
.B2(n_717),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_774),
.B(n_778),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_741),
.B(n_783),
.Y(n_848)
);

OAI211xp5_ASAP7_75t_L g849 ( 
.A1(n_730),
.A2(n_792),
.B(n_788),
.C(n_743),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_702),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_791),
.B(n_702),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_715),
.B(n_732),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_715),
.A2(n_787),
.B1(n_780),
.B2(n_779),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_731),
.B(n_732),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_787),
.B(n_695),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_701),
.A2(n_765),
.B1(n_770),
.B2(n_748),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_SL g857 ( 
.A1(n_789),
.A2(n_695),
.B1(n_723),
.B2(n_782),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_723),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_789),
.A2(n_773),
.B1(n_782),
.B2(n_749),
.Y(n_859)
);

BUFx4f_ASAP7_75t_SL g860 ( 
.A(n_744),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_766),
.B(n_744),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_754),
.A2(n_762),
.B1(n_781),
.B2(n_786),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_756),
.B(n_784),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_745),
.A2(n_540),
.B1(n_564),
.B2(n_521),
.Y(n_864)
);

BUFx4f_ASAP7_75t_SL g865 ( 
.A(n_755),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_745),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_836),
.A2(n_790),
.B1(n_837),
.B2(n_864),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_803),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_797),
.Y(n_869)
);

AND2x4_ASAP7_75t_SL g870 ( 
.A(n_804),
.B(n_855),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_SL g871 ( 
.A1(n_812),
.A2(n_860),
.B1(n_844),
.B2(n_864),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_810),
.B(n_824),
.C(n_796),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_855),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_794),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_840),
.B(n_806),
.Y(n_875)
);

OAI222xp33_ASAP7_75t_L g876 ( 
.A1(n_855),
.A2(n_863),
.B1(n_831),
.B2(n_796),
.C1(n_853),
.C2(n_865),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_843),
.A2(n_828),
.B(n_866),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_SL g878 ( 
.A1(n_830),
.A2(n_865),
.B1(n_860),
.B2(n_842),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_827),
.B(n_808),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_802),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_818),
.B(n_821),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_843),
.A2(n_846),
.B(n_828),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_831),
.B(n_832),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_832),
.A2(n_842),
.B1(n_809),
.B2(n_829),
.Y(n_884)
);

AOI33xp33_ASAP7_75t_L g885 ( 
.A1(n_801),
.A2(n_839),
.A3(n_835),
.B1(n_811),
.B2(n_820),
.B3(n_825),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_803),
.Y(n_886)
);

AOI33xp33_ASAP7_75t_L g887 ( 
.A1(n_841),
.A2(n_853),
.A3(n_815),
.B1(n_852),
.B2(n_824),
.B3(n_847),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_848),
.Y(n_888)
);

NAND3xp33_ASAP7_75t_L g889 ( 
.A(n_815),
.B(n_841),
.C(n_816),
.Y(n_889)
);

OAI22xp33_ASAP7_75t_L g890 ( 
.A1(n_813),
.A2(n_814),
.B1(n_793),
.B2(n_805),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_822),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_822),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_850),
.B(n_851),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_802),
.Y(n_894)
);

OAI322xp33_ASAP7_75t_L g895 ( 
.A1(n_854),
.A2(n_861),
.A3(n_833),
.B1(n_819),
.B2(n_856),
.C1(n_799),
.C2(n_800),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_833),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_849),
.A2(n_795),
.B1(n_822),
.B2(n_859),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_858),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_858),
.Y(n_899)
);

OAI31xp33_ASAP7_75t_L g900 ( 
.A1(n_823),
.A2(n_859),
.A3(n_862),
.B(n_798),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_845),
.B(n_857),
.C(n_834),
.Y(n_901)
);

OAI211xp5_ASAP7_75t_L g902 ( 
.A1(n_857),
.A2(n_862),
.B(n_807),
.C(n_826),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_845),
.A2(n_432),
.B1(n_597),
.B2(n_481),
.C(n_683),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_817),
.B(n_838),
.Y(n_904)
);

AOI221xp5_ASAP7_75t_L g905 ( 
.A1(n_817),
.A2(n_432),
.B1(n_597),
.B2(n_481),
.C(n_683),
.Y(n_905)
);

OAI22xp33_ASAP7_75t_L g906 ( 
.A1(n_855),
.A2(n_630),
.B1(n_621),
.B2(n_540),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_883),
.A2(n_903),
.B1(n_871),
.B2(n_867),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_SL g908 ( 
.A(n_891),
.B(n_892),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_868),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_879),
.B(n_883),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_877),
.B(n_874),
.Y(n_911)
);

NAND4xp25_ASAP7_75t_L g912 ( 
.A(n_905),
.B(n_878),
.C(n_884),
.D(n_897),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_888),
.B(n_885),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_877),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_885),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_872),
.A2(n_906),
.B1(n_889),
.B2(n_875),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_869),
.B(n_875),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_868),
.Y(n_918)
);

AOI221xp5_ASAP7_75t_L g919 ( 
.A1(n_876),
.A2(n_906),
.B1(n_884),
.B2(n_882),
.C(n_895),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_870),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_886),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_881),
.B(n_893),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_SL g923 ( 
.A1(n_870),
.A2(n_900),
.B(n_901),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_892),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_904),
.B(n_873),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_892),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_899),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_920),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_911),
.B(n_898),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_910),
.B(n_894),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_918),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_SL g932 ( 
.A(n_908),
.B(n_891),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_927),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_911),
.B(n_873),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_910),
.B(n_887),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_918),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_925),
.B(n_880),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_909),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_926),
.B(n_924),
.Y(n_939)
);

NAND4xp25_ASAP7_75t_SL g940 ( 
.A(n_916),
.B(n_887),
.C(n_902),
.D(n_892),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_921),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_940),
.A2(n_923),
.B(n_907),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_929),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_929),
.Y(n_944)
);

NAND2x1_ASAP7_75t_L g945 ( 
.A(n_931),
.B(n_926),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_938),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_938),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_934),
.B(n_927),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_937),
.B(n_925),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_935),
.B(n_915),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_928),
.B(n_912),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_933),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_931),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_952),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_949),
.B(n_937),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_942),
.A2(n_907),
.B1(n_912),
.B2(n_919),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_951),
.B(n_915),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_949),
.B(n_934),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_951),
.B(n_917),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_952),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_943),
.B(n_925),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_950),
.B(n_913),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_945),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_944),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_954),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_960),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_959),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_958),
.B(n_948),
.Y(n_968)
);

AOI221xp5_ASAP7_75t_L g969 ( 
.A1(n_957),
.A2(n_953),
.B1(n_930),
.B2(n_922),
.C(n_914),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_963),
.A2(n_932),
.B(n_939),
.Y(n_971)
);

OAI32xp33_ASAP7_75t_SL g972 ( 
.A1(n_956),
.A2(n_959),
.A3(n_957),
.B1(n_962),
.B2(n_955),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_955),
.B(n_932),
.Y(n_973)
);

XNOR2xp5_ASAP7_75t_L g974 ( 
.A(n_955),
.B(n_924),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_967),
.A2(n_914),
.B(n_890),
.C(n_896),
.Y(n_975)
);

OAI211xp5_ASAP7_75t_SL g976 ( 
.A1(n_973),
.A2(n_914),
.B(n_880),
.C(n_941),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_973),
.A2(n_961),
.B1(n_925),
.B2(n_946),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_965),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_978),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_977),
.Y(n_980)
);

OAI211xp5_ASAP7_75t_SL g981 ( 
.A1(n_975),
.A2(n_972),
.B(n_971),
.C(n_969),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_980),
.B(n_970),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_981),
.A2(n_976),
.B(n_966),
.C(n_968),
.Y(n_983)
);

NOR2x1p5_ASAP7_75t_L g984 ( 
.A(n_982),
.B(n_979),
.Y(n_984)
);

XNOR2xp5_ASAP7_75t_L g985 ( 
.A(n_983),
.B(n_974),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_984),
.Y(n_986)
);

OR3x1_ASAP7_75t_L g987 ( 
.A(n_985),
.B(n_941),
.C(n_936),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_986),
.Y(n_988)
);

XNOR2xp5_ASAP7_75t_L g989 ( 
.A(n_987),
.B(n_968),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_988),
.B(n_947),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_990),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_989),
.B1(n_890),
.B2(n_936),
.C(n_947),
.Y(n_992)
);


endmodule