module fake_jpeg_2809_n_231 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_231);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_83),
.Y(n_94)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_58),
.B1(n_70),
.B2(n_55),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_58),
.B1(n_70),
.B2(n_55),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_73),
.B(n_66),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_67),
.C(n_76),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_100),
.B(n_73),
.Y(n_140)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_59),
.B1(n_68),
.B2(n_80),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_112),
.Y(n_131)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_65),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_77),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_106),
.B1(n_105),
.B2(n_74),
.Y(n_123)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_129),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_89),
.B1(n_95),
.B2(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_130),
.B1(n_61),
.B2(n_64),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_89),
.B1(n_82),
.B2(n_59),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_140),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_89),
.C(n_54),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_4),
.C(n_6),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_62),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_77),
.B1(n_75),
.B2(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_63),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_26),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_144),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_147),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_68),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_34),
.Y(n_181)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_66),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_161),
.B(n_163),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_139),
.B1(n_122),
.B2(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_156),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_132),
.B1(n_10),
.B2(n_13),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_140),
.B(n_121),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_9),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_140),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_32),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_178),
.B1(n_179),
.B2(n_16),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_177),
.Y(n_190)
);

NOR2x1p5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_122),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_53),
.B(n_39),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_145),
.B1(n_148),
.B2(n_151),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_40),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_15),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_143),
.B(n_160),
.C(n_158),
.D(n_38),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_197),
.CI(n_48),
.CON(n_199),
.SN(n_199)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_185)
);

OAI22x1_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_164),
.B1(n_175),
.B2(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_189),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_36),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_194),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_17),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_19),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_42),
.B(n_51),
.Y(n_197)
);

AOI211xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_194),
.B(n_41),
.C(n_43),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_174),
.B1(n_167),
.B2(n_182),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_208),
.B1(n_192),
.B2(n_187),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_211),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_213),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_178),
.B1(n_184),
.B2(n_168),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.C(n_202),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_207),
.C(n_212),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_220),
.C(n_207),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_211),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_222),
.C(n_210),
.Y(n_226)
);

AOI31xp33_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_217),
.A3(n_198),
.B(n_205),
.Y(n_227)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_199),
.A3(n_24),
.B1(n_25),
.B2(n_27),
.C(n_29),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_44),
.B(n_47),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_229),
.B(n_49),
.Y(n_230)
);

AOI21x1_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_52),
.B(n_22),
.Y(n_231)
);


endmodule