module fake_jpeg_29686_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_38),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_1),
.CON(n_31),
.SN(n_31)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_23),
.Y(n_46)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_62),
.B1(n_39),
.B2(n_33),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_15),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_40),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_60),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_19),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_14),
.B1(n_19),
.B2(n_24),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_14),
.B1(n_37),
.B2(n_41),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_24),
.B1(n_12),
.B2(n_17),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_67),
.B(n_64),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_74),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_12),
.B1(n_17),
.B2(n_21),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_2),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_3),
.B1(n_58),
.B2(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_55),
.B(n_54),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_53),
.B(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_76),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_97),
.B(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_109),
.B1(n_90),
.B2(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_87),
.C(n_97),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_68),
.C(n_77),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_90),
.B(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_70),
.C(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_89),
.B1(n_96),
.B2(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_115),
.B(n_105),
.CI(n_112),
.CON(n_120),
.SN(n_120)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_108),
.B1(n_102),
.B2(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_103),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_123),
.B(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_124),
.C(n_125),
.Y(n_126)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.C(n_115),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_112),
.C(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_119),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_120),
.C(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_129),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_132),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_120),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_128),
.Y(n_138)
);


endmodule