module fake_netlist_6_527_n_1123 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1123);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1123;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_SL g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_143),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_29),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_105),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_133),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_109),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_87),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_122),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_60),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_97),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_131),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_180),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_40),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_178),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_132),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_77),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_93),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_106),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_139),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_2),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_84),
.Y(n_256)
);

BUFx8_ASAP7_75t_SL g257 ( 
.A(n_148),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_89),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_55),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_63),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_160),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_37),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_19),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_98),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_112),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_52),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_95),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_33),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_198),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_107),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_202),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_94),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_59),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_51),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_166),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_149),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_76),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_128),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_163),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_65),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_72),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_232),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_0),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_247),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_225),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_222),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_277),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_271),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_218),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_226),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_222),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_236),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_223),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_223),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_226),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_225),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_229),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_220),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_248),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_221),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_269),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_229),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_242),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_288),
.A2(n_249),
.B1(n_270),
.B2(n_237),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_242),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_238),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_253),
.B(n_282),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_334),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_238),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_217),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_291),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_337),
.A2(n_253),
.B(n_286),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_292),
.A2(n_281),
.B1(n_275),
.B2(n_237),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_316),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_294),
.A2(n_249),
.B1(n_270),
.B2(n_281),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g362 ( 
.A(n_298),
.B(n_295),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_224),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_303),
.B(n_227),
.Y(n_365)
);

BUFx8_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_294),
.A2(n_275),
.B1(n_278),
.B2(n_284),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_306),
.B(n_228),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_315),
.B(n_230),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_312),
.A2(n_287),
.B1(n_285),
.B2(n_283),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_315),
.A2(n_251),
.B1(n_273),
.B2(n_272),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_309),
.B(n_231),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_239),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_311),
.B(n_0),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_313),
.B(n_243),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_323),
.A2(n_245),
.B(n_244),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_290),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_293),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_301),
.A2(n_274),
.B1(n_268),
.B2(n_260),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_325),
.B(n_259),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_325),
.A2(n_258),
.B1(n_254),
.B2(n_250),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_246),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

CKINVDCx6p67_ASAP7_75t_R g402 ( 
.A(n_362),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_389),
.B(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_361),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_372),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

AO21x2_ASAP7_75t_L g413 ( 
.A1(n_346),
.A2(n_39),
.B(n_36),
.Y(n_413)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_343),
.A2(n_42),
.B(n_41),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_358),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_389),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_345),
.B(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_357),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_389),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_338),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_369),
.B(n_305),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_371),
.B(n_44),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_389),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_45),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_387),
.B(n_1),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_47),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_384),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_360),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_385),
.B(n_305),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_371),
.B(n_48),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_339),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_391),
.B(n_318),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_377),
.B(n_49),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_341),
.B(n_318),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_375),
.B(n_373),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_368),
.Y(n_460)
);

AND3x2_ASAP7_75t_L g461 ( 
.A(n_374),
.B(n_386),
.C(n_388),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_355),
.B(n_50),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_339),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_392),
.B(n_321),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_347),
.B(n_321),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_368),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_356),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_347),
.B(n_322),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_388),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_365),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_382),
.B(n_380),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_379),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_407),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_407),
.B(n_354),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_378),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_378),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_399),
.B(n_378),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_467),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_420),
.B(n_365),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_467),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_362),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_402),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_400),
.Y(n_494)
);

OR2x2_ASAP7_75t_SL g495 ( 
.A(n_436),
.B(n_383),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_440),
.A2(n_442),
.B(n_439),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_423),
.B(n_382),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_423),
.B(n_379),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_379),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_442),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_445),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_383),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_436),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_383),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_447),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_439),
.B(n_408),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_447),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_449),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_439),
.A2(n_380),
.B(n_381),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_432),
.B(n_381),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_431),
.B(n_322),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_443),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_430),
.B(n_380),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_443),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_430),
.B(n_390),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_444),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_438),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_444),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_455),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_408),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_431),
.B(n_376),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_437),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_408),
.A2(n_376),
.B(n_339),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_418),
.B(n_339),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_458),
.B(n_366),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_468),
.B(n_1),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_444),
.B(n_366),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_412),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_450),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_394),
.B(n_366),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_398),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_402),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_R g549 ( 
.A(n_422),
.B(n_53),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_417),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_421),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_513),
.B(n_433),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_490),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_505),
.B(n_516),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_491),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_422),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_481),
.B(n_451),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_505),
.B(n_454),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_492),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_503),
.B(n_418),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_516),
.A2(n_435),
.B(n_418),
.C(n_462),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_394),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_513),
.B(n_433),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_483),
.B(n_461),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_526),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_521),
.B(n_433),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_533),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_535),
.B(n_433),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_518),
.A2(n_456),
.B1(n_466),
.B2(n_424),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_541),
.B(n_454),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

AO22x1_ASAP7_75t_L g574 ( 
.A1(n_524),
.A2(n_433),
.B1(n_456),
.B2(n_339),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_475),
.B(n_421),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_535),
.B(n_433),
.Y(n_577)
);

NOR2xp67_ASAP7_75t_SL g578 ( 
.A(n_471),
.B(n_473),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_487),
.B(n_433),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_474),
.A2(n_460),
.B1(n_452),
.B2(n_453),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_533),
.B(n_452),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_507),
.A2(n_413),
.B1(n_404),
.B2(n_411),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_500),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_474),
.A2(n_460),
.B1(n_453),
.B2(n_466),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_538),
.B(n_454),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_528),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_482),
.B(n_424),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_482),
.B(n_409),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_507),
.A2(n_413),
.B1(n_409),
.B2(n_411),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_524),
.A2(n_463),
.B1(n_457),
.B2(n_448),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_547),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_499),
.B(n_469),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_476),
.A2(n_413),
.B1(n_395),
.B2(n_397),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_477),
.B(n_478),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_479),
.B(n_396),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_470),
.B(n_463),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_480),
.B(n_396),
.Y(n_599)
);

INVx8_ASAP7_75t_L g600 ( 
.A(n_521),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_545),
.B(n_506),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_551),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_539),
.B(n_396),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_484),
.A2(n_395),
.B1(n_397),
.B2(n_463),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_470),
.B(n_396),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_501),
.B(n_396),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_496),
.B(n_401),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_534),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_527),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_529),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_546),
.B(n_54),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_510),
.B(n_485),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_530),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_472),
.B(n_426),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_470),
.B(n_401),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_523),
.A2(n_457),
.B1(n_448),
.B2(n_429),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_502),
.B(n_426),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_504),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_567),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_567),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

OR2x6_ASAP7_75t_SL g623 ( 
.A(n_576),
.B(n_519),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_556),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_575),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_554),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_575),
.B(n_531),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_SL g629 ( 
.A(n_557),
.B(n_549),
.C(n_532),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_502),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_578),
.B(n_525),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_SL g632 ( 
.A(n_557),
.B(n_489),
.C(n_540),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_617),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_608),
.B(n_495),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_609),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_600),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_586),
.B(n_485),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_598),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_601),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_558),
.A2(n_546),
.B1(n_488),
.B2(n_486),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_597),
.A2(n_536),
.B(n_520),
.C(n_522),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_566),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_566),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_609),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_600),
.B(n_536),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

HAxp5_ASAP7_75t_L g648 ( 
.A(n_601),
.B(n_493),
.CON(n_648),
.SN(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_573),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_R g650 ( 
.A(n_562),
.B(n_548),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_579),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_597),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_R g653 ( 
.A(n_553),
.B(n_537),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_611),
.B(n_508),
.Y(n_655)
);

CKINVDCx8_ASAP7_75t_R g656 ( 
.A(n_598),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_594),
.B(n_509),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_612),
.B(n_512),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_569),
.B(n_514),
.Y(n_660)
);

AND3x1_ASAP7_75t_SL g661 ( 
.A(n_588),
.B(n_542),
.C(n_515),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_598),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_610),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_596),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_564),
.B(n_543),
.Y(n_665)
);

BUFx4f_ASAP7_75t_L g666 ( 
.A(n_613),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_587),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_544),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_580),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_602),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_617),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_603),
.A2(n_552),
.B(n_550),
.C(n_537),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_616),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_570),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_498),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_555),
.B(n_511),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_599),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_577),
.A2(n_457),
.B(n_448),
.C(n_429),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_582),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_555),
.B(n_2),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_590),
.B(n_3),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_637),
.A2(n_563),
.B(n_559),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_624),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_640),
.B(n_592),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_636),
.Y(n_686)
);

OAI22x1_ASAP7_75t_L g687 ( 
.A1(n_681),
.A2(n_581),
.B1(n_585),
.B2(n_559),
.Y(n_687)
);

AOI21x1_ASAP7_75t_L g688 ( 
.A1(n_641),
.A2(n_574),
.B(n_589),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_675),
.A2(n_572),
.B(n_571),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_649),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_664),
.B(n_607),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_625),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_635),
.B(n_662),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_660),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_680),
.B(n_604),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

OAI22x1_ASAP7_75t_L g697 ( 
.A1(n_681),
.A2(n_414),
.B1(n_614),
.B2(n_591),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_677),
.A2(n_414),
.B(n_595),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_620),
.Y(n_699)
);

NOR2x1_ASAP7_75t_L g700 ( 
.A(n_633),
.B(n_401),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_640),
.B(n_643),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_L g702 ( 
.A1(n_632),
.A2(n_591),
.B(n_583),
.Y(n_702)
);

CKINVDCx8_ASAP7_75t_R g703 ( 
.A(n_645),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_657),
.B(n_401),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_632),
.B(n_415),
.C(n_401),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_669),
.A2(n_429),
.B(n_415),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_665),
.A2(n_429),
.B(n_415),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_634),
.B(n_415),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_635),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_652),
.B(n_429),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_630),
.B(n_448),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_650),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_631),
.A2(n_457),
.B(n_448),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_636),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_665),
.A2(n_457),
.B(n_426),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_619),
.Y(n_716)
);

AO31x2_ASAP7_75t_L g717 ( 
.A1(n_679),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

AND2x2_ASAP7_75t_SL g719 ( 
.A(n_673),
.B(n_4),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_652),
.B(n_5),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_658),
.A2(n_426),
.B(n_61),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_682),
.A2(n_426),
.B(n_7),
.C(n_8),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_647),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_629),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_724)
);

AOI21x1_ASAP7_75t_L g725 ( 
.A1(n_641),
.A2(n_62),
.B(n_58),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_621),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_658),
.A2(n_66),
.B(n_64),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_666),
.B(n_6),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_672),
.A2(n_68),
.B(n_67),
.Y(n_729)
);

NOR2x1_ASAP7_75t_R g730 ( 
.A(n_644),
.B(n_69),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_655),
.A2(n_73),
.B(n_71),
.Y(n_731)
);

AO21x1_ASAP7_75t_L g732 ( 
.A1(n_673),
.A2(n_9),
.B(n_10),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_678),
.A2(n_135),
.B(n_215),
.Y(n_733)
);

BUFx4f_ASAP7_75t_SL g734 ( 
.A(n_647),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_627),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_642),
.A2(n_134),
.B(n_214),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_L g737 ( 
.A1(n_629),
.A2(n_10),
.B(n_12),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_630),
.B(n_74),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_674),
.B(n_12),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_735),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_SL g741 ( 
.A(n_703),
.B(n_638),
.Y(n_741)
);

AOI21x1_ASAP7_75t_L g742 ( 
.A1(n_688),
.A2(n_646),
.B(n_676),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_736),
.A2(n_729),
.B(n_702),
.C(n_694),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_734),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_706),
.A2(n_671),
.B(n_633),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_SL g746 ( 
.A(n_730),
.B(n_656),
.Y(n_746)
);

CKINVDCx6p67_ASAP7_75t_R g747 ( 
.A(n_686),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_684),
.Y(n_748)
);

OA21x2_ASAP7_75t_L g749 ( 
.A1(n_698),
.A2(n_670),
.B(n_676),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_737),
.A2(n_666),
.B(n_651),
.C(n_639),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

AO31x2_ASAP7_75t_L g752 ( 
.A1(n_697),
.A2(n_661),
.A3(n_663),
.B(n_667),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_691),
.A2(n_638),
.B(n_646),
.Y(n_753)
);

OA21x2_ASAP7_75t_L g754 ( 
.A1(n_707),
.A2(n_668),
.B(n_661),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_683),
.A2(n_638),
.B(n_671),
.Y(n_755)
);

BUFx12f_ASAP7_75t_L g756 ( 
.A(n_712),
.Y(n_756)
);

OAI21x1_ASAP7_75t_L g757 ( 
.A1(n_713),
.A2(n_622),
.B(n_626),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_709),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_724),
.A2(n_728),
.B(n_722),
.C(n_720),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_SL g760 ( 
.A1(n_685),
.A2(n_695),
.B(n_739),
.C(n_689),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_721),
.A2(n_668),
.B(n_628),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_701),
.B(n_628),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_727),
.A2(n_626),
.B(n_622),
.C(n_654),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_719),
.A2(n_653),
.B1(n_647),
.B2(n_648),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_686),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_686),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_708),
.A2(n_705),
.B(n_731),
.C(n_738),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_725),
.A2(n_653),
.B(n_140),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_693),
.B(n_623),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_687),
.A2(n_216),
.B(n_136),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_693),
.B(n_75),
.Y(n_771)
);

AO31x2_ASAP7_75t_L g772 ( 
.A1(n_732),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_690),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_696),
.Y(n_774)
);

CKINVDCx11_ASAP7_75t_R g775 ( 
.A(n_714),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_715),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_704),
.A2(n_17),
.B(n_18),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_726),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_710),
.A2(n_144),
.B(n_213),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_SL g780 ( 
.A(n_714),
.B(n_718),
.Y(n_780)
);

O2A1O1Ixp5_ASAP7_75t_L g781 ( 
.A1(n_716),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_716),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_733),
.A2(n_20),
.B(n_21),
.Y(n_783)
);

CKINVDCx11_ASAP7_75t_R g784 ( 
.A(n_714),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_699),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_738),
.A2(n_145),
.B(n_211),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_718),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_700),
.A2(n_142),
.B(n_210),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_711),
.B(n_22),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_717),
.A2(n_23),
.A3(n_24),
.B(n_25),
.Y(n_790)
);

OAI22x1_ASAP7_75t_L g791 ( 
.A1(n_711),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_718),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_723),
.B(n_26),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_723),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_706),
.A2(n_141),
.B(n_206),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_736),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_797)
);

AOI21x1_ASAP7_75t_SL g798 ( 
.A1(n_720),
.A2(n_30),
.B(n_31),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_694),
.A2(n_151),
.B(n_205),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_719),
.B(n_30),
.Y(n_800)
);

AO21x1_ASAP7_75t_L g801 ( 
.A1(n_729),
.A2(n_31),
.B(n_32),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_684),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_694),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_803)
);

AO32x2_ASAP7_75t_L g804 ( 
.A1(n_732),
.A2(n_34),
.A3(n_35),
.B1(n_78),
.B2(n_79),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_724),
.A2(n_35),
.B(n_80),
.C(n_81),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_764),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_782),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_801),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_740),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_748),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_800),
.A2(n_92),
.B1(n_96),
.B2(n_99),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_751),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_777),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_803),
.A2(n_103),
.B1(n_104),
.B2(n_108),
.Y(n_814)
);

INVx6_ASAP7_75t_L g815 ( 
.A(n_744),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_785),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_773),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_746),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_774),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_802),
.Y(n_820)
);

INVx6_ASAP7_75t_L g821 ( 
.A(n_744),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_790),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_790),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_790),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_789),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_791),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_SL g827 ( 
.A1(n_783),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_762),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_792),
.Y(n_829)
);

CKINVDCx6p67_ASAP7_75t_R g830 ( 
.A(n_775),
.Y(n_830)
);

BUFx10_ASAP7_75t_L g831 ( 
.A(n_787),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_SL g832 ( 
.A1(n_795),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_756),
.A2(n_129),
.B1(n_138),
.B2(n_147),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_769),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_784),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_758),
.Y(n_836)
);

CKINVDCx6p67_ASAP7_75t_R g837 ( 
.A(n_747),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_765),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_776),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_761),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_797),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_743),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_760),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_750),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_844)
);

HB1xp67_ASAP7_75t_SL g845 ( 
.A(n_793),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_752),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_765),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_765),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_770),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_849)
);

INVx4_ASAP7_75t_SL g850 ( 
.A(n_772),
.Y(n_850)
);

INVx6_ASAP7_75t_L g851 ( 
.A(n_780),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_759),
.B(n_179),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_766),
.B(n_181),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_794),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_767),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_771),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_754),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_745),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_772),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_772),
.Y(n_860)
);

CKINVDCx11_ASAP7_75t_R g861 ( 
.A(n_741),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_798),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_753),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_749),
.Y(n_864)
);

BUFx4f_ASAP7_75t_SL g865 ( 
.A(n_786),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_822),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_823),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_858),
.B(n_742),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_863),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_830),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_864),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_807),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_857),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_810),
.B(n_804),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_820),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_839),
.A2(n_768),
.B(n_796),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_846),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_824),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_817),
.B(n_804),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_819),
.B(n_859),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_847),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_860),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_828),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_842),
.A2(n_805),
.B(n_841),
.C(n_808),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_816),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_855),
.A2(n_755),
.B(n_749),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_850),
.B(n_804),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_850),
.B(n_754),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_843),
.A2(n_757),
.B(n_799),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_809),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_829),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_862),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_829),
.B(n_763),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_854),
.B(n_778),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_862),
.Y(n_896)
);

CKINVDCx11_ASAP7_75t_R g897 ( 
.A(n_835),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_845),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_865),
.A2(n_779),
.B1(n_788),
.B2(n_781),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_843),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_852),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_844),
.A2(n_189),
.B(n_190),
.Y(n_902)
);

INVx4_ASAP7_75t_SL g903 ( 
.A(n_851),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_808),
.A2(n_192),
.B(n_193),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_836),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_842),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_851),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_861),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_840),
.A2(n_194),
.B(n_195),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_853),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_907),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_871),
.B(n_848),
.Y(n_912)
);

NAND4xp25_ASAP7_75t_L g913 ( 
.A(n_895),
.B(n_841),
.C(n_826),
.D(n_813),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_893),
.A2(n_806),
.B(n_853),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_871),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_873),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_L g917 ( 
.A(n_885),
.B(n_827),
.C(n_814),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_871),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_874),
.B(n_812),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_886),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_880),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_880),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_874),
.B(n_838),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_873),
.B(n_835),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_892),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_883),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_877),
.B(n_838),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_882),
.Y(n_928)
);

BUFx4f_ASAP7_75t_SL g929 ( 
.A(n_905),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_882),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_877),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_884),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_893),
.A2(n_887),
.B(n_868),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_866),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_879),
.B(n_835),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_877),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_890),
.A2(n_825),
.B(n_834),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_878),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_866),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_867),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_886),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_887),
.A2(n_837),
.B(n_849),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_872),
.B(n_867),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_916),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_918),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_916),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_915),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_915),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_918),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_935),
.B(n_919),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_936),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_926),
.B(n_901),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_932),
.B(n_921),
.Y(n_953)
);

AND2x4_ASAP7_75t_SL g954 ( 
.A(n_912),
.B(n_894),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_918),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_936),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_929),
.B(n_869),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_943),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_925),
.B(n_919),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_911),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_935),
.B(n_888),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_936),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_936),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_923),
.B(n_888),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_943),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_911),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_931),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_931),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_931),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_920),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_964),
.B(n_923),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_959),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_946),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_958),
.B(n_908),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_951),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_964),
.B(n_924),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_965),
.B(n_911),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_944),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_966),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_947),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_961),
.B(n_924),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_947),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_944),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_950),
.B(n_953),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_948),
.Y(n_985)
);

INVx4_ASAP7_75t_SL g986 ( 
.A(n_944),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_951),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_974),
.B(n_869),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_980),
.B(n_970),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_972),
.B(n_950),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_961),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_982),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_981),
.B(n_946),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_982),
.B(n_948),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_983),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_985),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_978),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_985),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_976),
.B(n_954),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_973),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_990),
.B(n_984),
.Y(n_1001)
);

NOR2x1_ASAP7_75t_L g1002 ( 
.A(n_988),
.B(n_983),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_1000),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_999),
.B(n_976),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_991),
.B(n_973),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_995),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_993),
.B(n_977),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_992),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_989),
.B(n_997),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_1006),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_989),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1009),
.B(n_971),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_1004),
.Y(n_1013)
);

OAI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_1005),
.A2(n_900),
.B1(n_917),
.B2(n_978),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_1008),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_1012),
.B(n_1001),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1015),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1011),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_1007),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1014),
.B(n_996),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1010),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_1010),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1012),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_1012),
.B(n_998),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_1013),
.A2(n_913),
.B1(n_906),
.B2(n_900),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1022),
.B(n_978),
.Y(n_1026)
);

OAI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_1022),
.A2(n_979),
.B1(n_957),
.B2(n_908),
.C(n_898),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1017),
.B(n_986),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_1018),
.B(n_897),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_1021),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1024),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_908),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1019),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1031),
.B(n_1016),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1027),
.A2(n_1023),
.B(n_1025),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1028),
.B(n_1029),
.Y(n_1036)
);

AOI211xp5_ASAP7_75t_L g1037 ( 
.A1(n_1033),
.A2(n_908),
.B(n_870),
.C(n_818),
.Y(n_1037)
);

AND2x2_ASAP7_75t_SL g1038 ( 
.A(n_1026),
.B(n_908),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_SL g1039 ( 
.A(n_1032),
.B(n_908),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_869),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1035),
.A2(n_904),
.B(n_907),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1038),
.A2(n_994),
.B(n_904),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1034),
.A2(n_906),
.B(n_994),
.C(n_833),
.Y(n_1043)
);

AOI221xp5_ASAP7_75t_L g1044 ( 
.A1(n_1039),
.A2(n_899),
.B1(n_811),
.B2(n_896),
.C(n_960),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1040),
.Y(n_1045)
);

INVxp33_ASAP7_75t_SL g1046 ( 
.A(n_1045),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1041),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1044),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1043),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1042),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1045),
.Y(n_1051)
);

OAI322xp33_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_1036),
.A3(n_1037),
.B1(n_987),
.B2(n_975),
.C1(n_953),
.C2(n_986),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_1048),
.B(n_832),
.C(n_831),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_1049),
.B(n_831),
.C(n_896),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_L g1055 ( 
.A(n_1050),
.B(n_1047),
.Y(n_1055)
);

OAI211xp5_ASAP7_75t_L g1056 ( 
.A1(n_1050),
.A2(n_1046),
.B(n_856),
.C(n_942),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1051),
.B(n_971),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_1056),
.B(n_1055),
.C(n_1054),
.Y(n_1058)
);

AOI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_1052),
.A2(n_960),
.B1(n_896),
.B2(n_987),
.C(n_975),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_1053),
.B(n_815),
.C(n_821),
.Y(n_1060)
);

AND4x1_ASAP7_75t_L g1061 ( 
.A(n_1057),
.B(n_821),
.C(n_815),
.D(n_986),
.Y(n_1061)
);

OAI211xp5_ASAP7_75t_L g1062 ( 
.A1(n_1056),
.A2(n_960),
.B(n_986),
.C(n_942),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_1058),
.B(n_901),
.C(n_969),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1060),
.A2(n_903),
.B1(n_954),
.B2(n_901),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_L g1065 ( 
.A(n_1062),
.B(n_914),
.C(n_902),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1061),
.B(n_968),
.Y(n_1066)
);

NAND4xp25_ASAP7_75t_SL g1067 ( 
.A(n_1059),
.B(n_910),
.C(n_951),
.D(n_956),
.Y(n_1067)
);

NAND4xp75_ASAP7_75t_L g1068 ( 
.A(n_1059),
.B(n_910),
.C(n_963),
.D(n_956),
.Y(n_1068)
);

AOI221xp5_ASAP7_75t_L g1069 ( 
.A1(n_1058),
.A2(n_954),
.B1(n_969),
.B2(n_967),
.C(n_955),
.Y(n_1069)
);

NAND4xp25_ASAP7_75t_L g1070 ( 
.A(n_1058),
.B(n_881),
.C(n_894),
.D(n_912),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_1068),
.Y(n_1071)
);

NAND4xp75_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_956),
.C(n_963),
.D(n_903),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_1070),
.B(n_197),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_1066),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1064),
.A2(n_914),
.B(n_894),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1063),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_L g1077 ( 
.A(n_1067),
.B(n_902),
.C(n_909),
.Y(n_1077)
);

AOI221x1_ASAP7_75t_L g1078 ( 
.A1(n_1065),
.A2(n_963),
.B1(n_967),
.B2(n_955),
.C(n_962),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_L g1079 ( 
.A(n_1070),
.B(n_909),
.C(n_937),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1074),
.Y(n_1080)
);

NAND4xp75_ASAP7_75t_L g1081 ( 
.A(n_1073),
.B(n_199),
.C(n_200),
.D(n_201),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1071),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1079),
.A2(n_894),
.B1(n_912),
.B2(n_903),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_1075),
.B(n_203),
.Y(n_1084)
);

AND3x4_ASAP7_75t_L g1085 ( 
.A(n_1077),
.B(n_881),
.C(n_912),
.Y(n_1085)
);

NAND4xp75_ASAP7_75t_L g1086 ( 
.A(n_1078),
.B(n_1076),
.C(n_1072),
.D(n_207),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1076),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_1074),
.B(n_881),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1071),
.Y(n_1089)
);

AND3x4_ASAP7_75t_L g1090 ( 
.A(n_1073),
.B(n_927),
.C(n_903),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_1071),
.B(n_937),
.C(n_933),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_1071),
.B(n_933),
.C(n_890),
.Y(n_1092)
);

AOI222xp33_ASAP7_75t_L g1093 ( 
.A1(n_1087),
.A2(n_903),
.B1(n_968),
.B2(n_949),
.C1(n_945),
.C2(n_872),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_1088),
.Y(n_1094)
);

AOI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1082),
.A2(n_968),
.B1(n_949),
.B2(n_945),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_1089),
.B(n_891),
.C(n_876),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1081),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1084),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1080),
.B(n_962),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1090),
.A2(n_938),
.B1(n_927),
.B2(n_868),
.Y(n_1100)
);

OAI22x1_ASAP7_75t_L g1101 ( 
.A1(n_1094),
.A2(n_1085),
.B1(n_1086),
.B2(n_1083),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_1098),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1097),
.A2(n_1092),
.B1(n_1091),
.B2(n_938),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1099),
.A2(n_938),
.B1(n_927),
.B2(n_868),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1095),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1100),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1102),
.A2(n_1093),
.B1(n_1096),
.B2(n_938),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1101),
.A2(n_938),
.B1(n_927),
.B2(n_875),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1105),
.B(n_891),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1108),
.A2(n_1103),
.B1(n_1106),
.B2(n_1107),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1110),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1111),
.B(n_1109),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_1104),
.B1(n_938),
.B2(n_922),
.Y(n_1114)
);

AO22x2_ASAP7_75t_L g1115 ( 
.A1(n_1112),
.A2(n_939),
.B1(n_930),
.B2(n_934),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1113),
.A2(n_922),
.B1(n_921),
.B2(n_868),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1114),
.A2(n_875),
.B(n_876),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_930),
.B(n_939),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_879),
.Y(n_1119)
);

NOR3xp33_ASAP7_75t_L g1120 ( 
.A(n_1117),
.B(n_889),
.C(n_940),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1119),
.A2(n_934),
.B(n_940),
.Y(n_1121)
);

AOI22x1_ASAP7_75t_SL g1122 ( 
.A1(n_1120),
.A2(n_1118),
.B1(n_928),
.B2(n_941),
.Y(n_1122)
);

AOI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_889),
.C(n_928),
.Y(n_1123)
);


endmodule