module fake_netlist_1_6965_n_37 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
BUFx2_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
BUFx3_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_9), .B(n_0), .Y(n_20) );
NAND2xp33_ASAP7_75t_R g21 ( .A(n_20), .B(n_11), .Y(n_21) );
NAND2xp33_ASAP7_75t_R g22 ( .A(n_19), .B(n_11), .Y(n_22) );
NAND2x1p5_ASAP7_75t_L g23 ( .A(n_18), .B(n_12), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_17), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_16), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
OAI321xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_27), .A3(n_15), .B1(n_21), .B2(n_0), .C(n_2), .Y(n_30) );
O2A1O1Ixp33_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_2), .B(n_15), .C(n_6), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_31), .B(n_15), .Y(n_32) );
CKINVDCx14_ASAP7_75t_R g33 ( .A(n_30), .Y(n_33) );
BUFx2_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
INVx3_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_37) );
endmodule