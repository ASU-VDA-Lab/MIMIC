module fake_jpeg_31223_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_49),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_13),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_54),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_0),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_21),
.C(n_19),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_17),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_64),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_23),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_11),
.Y(n_65)
);

INVx2_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_66),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_27),
.Y(n_74)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_81),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_83),
.B1(n_99),
.B2(n_108),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_26),
.B1(n_38),
.B2(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_100),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_115),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_71),
.B1(n_55),
.B2(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_107),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_38),
.B1(n_40),
.B2(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_21),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_7),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_7),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_43),
.A2(n_38),
.B1(n_19),
.B2(n_18),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_18),
.B1(n_17),
.B2(n_3),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_121),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_63),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_132),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_89),
.B1(n_97),
.B2(n_84),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_105),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_136),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_11),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_145),
.Y(n_167)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_102),
.B(n_116),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_97),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_130),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_94),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_103),
.C(n_82),
.Y(n_154)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_149),
.B1(n_133),
.B2(n_125),
.Y(n_178)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_83),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_131),
.B(n_122),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_148),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_84),
.B1(n_105),
.B2(n_91),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_96),
.B1(n_75),
.B2(n_112),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_167),
.B1(n_152),
.B2(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_124),
.B(n_79),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_89),
.B1(n_79),
.B2(n_114),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_122),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_131),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_117),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_118),
.B(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_120),
.B(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_173),
.Y(n_179)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_194),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_193),
.B(n_196),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_153),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_197),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_153),
.C(n_175),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_161),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_159),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_184),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_154),
.C(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_218),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_183),
.B1(n_160),
.B2(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_164),
.Y(n_218)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_199),
.B1(n_200),
.B2(n_211),
.C(n_188),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_224),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_195),
.A3(n_181),
.B1(n_192),
.B2(n_158),
.C1(n_183),
.C2(n_174),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_221),
.B(n_206),
.C(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_152),
.B1(n_159),
.B2(n_193),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_225),
.B(n_150),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_151),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_222),
.C(n_213),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_205),
.B1(n_201),
.B2(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_233),
.B1(n_226),
.B2(n_216),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_205),
.B1(n_201),
.B2(n_166),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_222),
.C(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_229),
.C(n_194),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_232),
.B(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_235),
.B1(n_227),
.B2(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_131),
.B1(n_179),
.B2(n_209),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_241),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_238),
.A3(n_229),
.B1(n_244),
.B2(n_239),
.C1(n_182),
.C2(n_189),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_209),
.B(n_186),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_SL g257 ( 
.A(n_254),
.B(n_247),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_250),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_260),
.A3(n_246),
.B1(n_185),
.B2(n_156),
.C1(n_168),
.C2(n_134),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_247),
.B(n_248),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_261),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_168),
.A3(n_179),
.B1(n_134),
.B2(n_128),
.C1(n_122),
.C2(n_123),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);


endmodule