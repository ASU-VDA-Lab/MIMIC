module fake_jpeg_9127_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_23),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_32),
.B1(n_16),
.B2(n_30),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_30),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_32),
.B1(n_16),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_18),
.B1(n_19),
.B2(n_2),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_29),
.B1(n_22),
.B2(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_47),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_28),
.C(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2x1_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_23),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_64),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_68),
.B1(n_76),
.B2(n_78),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_70),
.B1(n_73),
.B2(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_68)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_83),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_54),
.B1(n_60),
.B2(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_0),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_4),
.B(n_5),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_3),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_59),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_46),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_4),
.B(n_6),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_7),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_7),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_80),
.B1(n_67),
.B2(n_11),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_72),
.C(n_78),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_107),
.C(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_108),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_81),
.C(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_92),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_70),
.B1(n_79),
.B2(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_117),
.B1(n_102),
.B2(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_120),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_71),
.C(n_69),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_118),
.A2(n_95),
.B(n_87),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_130),
.B(n_118),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_90),
.C(n_87),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_133),
.C(n_135),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_93),
.B(n_101),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_98),
.C(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_136),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_84),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_111),
.C(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_135),
.C(n_129),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_146),
.B(n_119),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_89),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_100),
.A3(n_121),
.B1(n_120),
.B2(n_103),
.C1(n_119),
.C2(n_9),
.Y(n_147)
);

AOI321xp33_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.C(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_155),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_141),
.B(n_89),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_124),
.B1(n_133),
.B2(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_143),
.B1(n_138),
.B2(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_88),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_124),
.B1(n_145),
.B2(n_140),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_163),
.B(n_164),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_168),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_10),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.C(n_163),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_159),
.C(n_158),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_158),
.B(n_77),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_174),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_173),
.Y(n_178)
);


endmodule