module fake_jpeg_15855_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_53),
.B1(n_24),
.B2(n_26),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_20),
.B1(n_27),
.B2(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_15),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_26),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_60),
.B1(n_67),
.B2(n_72),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_15),
.C(n_28),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_79),
.C(n_6),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_36),
.B1(n_21),
.B2(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_25),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_55),
.B1(n_44),
.B2(n_25),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_0),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_30),
.B1(n_29),
.B2(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_30),
.C(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NOR4xp25_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_3),
.C(n_4),
.D(n_6),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_4),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_4),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_83),
.B(n_64),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_77),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_116),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_114),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_76),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_60),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_80),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_122),
.B(n_99),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_67),
.B(n_79),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_125),
.B(n_100),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_14),
.C(n_8),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_128),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_78),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_106),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_133),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_126),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_88),
.B(n_91),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_114),
.B(n_115),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_87),
.B1(n_91),
.B2(n_107),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_145),
.B1(n_147),
.B2(n_116),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_109),
.C(n_107),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_151),
.C(n_153),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_94),
.B1(n_105),
.B2(n_108),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_108),
.B1(n_105),
.B2(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_94),
.B1(n_109),
.B2(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_99),
.C(n_74),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_84),
.C(n_106),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_133),
.B(n_130),
.C(n_132),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_112),
.B(n_124),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_119),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_166),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_167),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_117),
.B1(n_106),
.B2(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_180),
.B1(n_135),
.B2(n_129),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_110),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_139),
.B(n_146),
.C(n_140),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_169),
.B(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_173),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_178),
.B1(n_151),
.B2(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_175),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_143),
.C(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_190),
.C(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_142),
.C(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_142),
.C(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_175),
.B1(n_158),
.B2(n_178),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_165),
.C(n_180),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_198),
.C(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_174),
.C(n_160),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_163),
.C(n_177),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_150),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_206),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_168),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_186),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_152),
.B1(n_168),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_168),
.B1(n_140),
.B2(n_156),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_193),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_187),
.B(n_168),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_SL g211 ( 
.A(n_208),
.B(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_186),
.C(n_185),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_218),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_201),
.A2(n_156),
.B1(n_182),
.B2(n_194),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_203),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_213),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_230),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_210),
.B1(n_212),
.B2(n_208),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_156),
.C(n_171),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_222),
.B(n_225),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_113),
.A3(n_90),
.B1(n_11),
.B2(n_12),
.C1(n_7),
.C2(n_10),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_225),
.B1(n_90),
.B2(n_113),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_238),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_10),
.B(n_12),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_235),
.C(n_84),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_13),
.Y(n_243)
);


endmodule