module fake_jpeg_3279_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_47),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_34),
.Y(n_79)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_61),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_36),
.B1(n_46),
.B2(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_39),
.B1(n_38),
.B2(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_3),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_52),
.C(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_34),
.Y(n_85)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_43),
.B1(n_44),
.B2(n_39),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_69),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_43),
.B(n_39),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_88),
.B1(n_76),
.B2(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_5),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_7),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_7),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_8),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_102),
.B1(n_103),
.B2(n_109),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_76),
.B(n_78),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_23),
.B(n_25),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_75),
.C(n_70),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.C(n_15),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_13),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_116),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_115),
.B1(n_102),
.B2(n_106),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_28),
.C(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_115),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_119),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_100),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_118),
.B(n_101),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_111),
.C(n_110),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_97),
.Y(n_128)
);


endmodule