module fake_jpeg_13610_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_21),
.C(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_76),
.C(n_72),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_19),
.B(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_79),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_50),
.C(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_0),
.Y(n_110)
);

INVx13_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_81),
.B1(n_80),
.B2(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_95),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_55),
.B1(n_68),
.B2(n_61),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_53),
.B1(n_65),
.B2(n_57),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_52),
.B(n_60),
.C(n_69),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_93),
.B(n_96),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_55),
.B1(n_68),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_72),
.B1(n_53),
.B2(n_67),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_58),
.B1(n_63),
.B2(n_52),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_51),
.B(n_54),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_64),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_103),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_114),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_93),
.B1(n_88),
.B2(n_94),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_73),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_64),
.B1(n_39),
.B2(n_37),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_1),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_124),
.B1(n_115),
.B2(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_64),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_1),
.B(n_4),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_132),
.B(n_14),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_36),
.C(n_35),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_135),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_5),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_138),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_6),
.B(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_34),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_32),
.C(n_31),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_29),
.C(n_28),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_27),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_144)
);

BUFx12f_ASAP7_75t_SL g145 ( 
.A(n_125),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_146),
.B(n_147),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_15),
.B(n_16),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_16),
.B(n_17),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_152),
.B(n_136),
.Y(n_158)
);

XNOR2x2_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_17),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_146),
.C(n_147),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_156),
.B(n_149),
.C(n_133),
.D(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

AO221x1_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_134),
.B1(n_150),
.B2(n_137),
.C(n_145),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_126),
.C(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_162),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_164),
.B(n_159),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_138),
.A3(n_139),
.B1(n_157),
.B2(n_154),
.C1(n_119),
.C2(n_152),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_157),
.C(n_137),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_119),
.Y(n_169)
);


endmodule