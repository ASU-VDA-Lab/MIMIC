module fake_jpeg_16159_n_291 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_291);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_18),
.B1(n_23),
.B2(n_16),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_23),
.B1(n_16),
.B2(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_19),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_14),
.B1(n_18),
.B2(n_20),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_39),
.B1(n_49),
.B2(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_14),
.B1(n_39),
.B2(n_20),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_25),
.B(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_65),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_16),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_86),
.B1(n_56),
.B2(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_84),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_82),
.B(n_77),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_21),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_19),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_11),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_50),
.A3(n_69),
.B1(n_54),
.B2(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_42),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_100),
.B1(n_73),
.B2(n_90),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_51),
.B1(n_58),
.B2(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_99),
.B1(n_102),
.B2(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_51),
.C(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_110),
.B(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_63),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_61),
.B1(n_68),
.B2(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_61),
.B1(n_45),
.B2(n_67),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_45),
.B1(n_28),
.B2(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_74),
.B1(n_42),
.B2(n_40),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_75),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_60),
.B1(n_45),
.B2(n_17),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_85),
.B(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_40),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_71),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_71),
.B(n_19),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_125),
.B(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_72),
.A3(n_83),
.B1(n_82),
.B2(n_78),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_72),
.B1(n_83),
.B2(n_76),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_121),
.B1(n_92),
.B2(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_76),
.B1(n_80),
.B2(n_86),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_130),
.B(n_102),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_85),
.B1(n_76),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_94),
.B1(n_103),
.B2(n_29),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_17),
.B1(n_13),
.B2(n_15),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_42),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_154),
.B1(n_155),
.B2(n_160),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_95),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_146),
.C(n_133),
.Y(n_163)
);

NAND2xp67_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_125),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_153),
.B(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_147),
.B1(n_131),
.B2(n_127),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_121),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_94),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_30),
.B1(n_74),
.B2(n_40),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_40),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_26),
.B(n_15),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_30),
.B1(n_40),
.B2(n_19),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_19),
.B1(n_36),
.B2(n_24),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_8),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_8),
.B(n_12),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_8),
.B1(n_11),
.B2(n_2),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_167),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_133),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_163),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_118),
.Y(n_171)
);

NOR4xp25_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_176),
.C(n_183),
.D(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_114),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_144),
.B1(n_149),
.B2(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_115),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_111),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_148),
.B(n_138),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_111),
.C(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_181),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_159),
.C(n_160),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_8),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_26),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_7),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_184),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_26),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_7),
.Y(n_184)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_199),
.B1(n_170),
.B2(n_173),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_166),
.B1(n_184),
.B2(n_163),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_194),
.B(n_171),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_144),
.B1(n_141),
.B2(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_206),
.B1(n_7),
.B2(n_11),
.Y(n_218)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_142),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_181),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_153),
.Y(n_205)
);

AOI211xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_13),
.B(n_24),
.C(n_2),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_155),
.B1(n_154),
.B2(n_2),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_221),
.Y(n_231)
);

XOR2x2_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_183),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_186),
.B(n_208),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_178),
.B1(n_173),
.B2(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_210),
.B(n_222),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_162),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_219),
.C(n_187),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_15),
.C(n_13),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_188),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_6),
.B1(n_10),
.B2(n_2),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_191),
.B1(n_199),
.B2(n_201),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_198),
.C(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_236),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_196),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_24),
.C(n_5),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_216),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_5),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_211),
.B1(n_209),
.B2(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_207),
.B1(n_190),
.B2(n_219),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_190),
.B1(n_9),
.B2(n_3),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_227),
.B(n_5),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_250),
.B(n_239),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_240),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_264),
.C(n_265),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_234),
.B1(n_231),
.B2(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_254),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_231),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_24),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_247),
.B(n_9),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_252),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_24),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_242),
.B1(n_245),
.B2(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_272),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_268),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_24),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_271),
.Y(n_276)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_260),
.C(n_257),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_3),
.B(n_4),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_273),
.B(n_274),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_3),
.B(n_4),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_280),
.C(n_275),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_11),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.C(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_282),
.C(n_4),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_10),
.B(n_0),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_0),
.Y(n_290)
);

OAI31xp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_1),
.A3(n_10),
.B(n_283),
.Y(n_291)
);


endmodule