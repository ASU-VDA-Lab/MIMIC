module fake_netlist_6_2635_n_785 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_785);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_785;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_38),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_24),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_27),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_74),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_86),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_35),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_25),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_51),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_8),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_21),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_61),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_6),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_26),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_45),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_149),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_57),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_56),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_50),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_60),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_112),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_22),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_49),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_130),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_106),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_7),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_87),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

OAI22x1_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_0),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_1),
.B(n_2),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_199),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_170),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_227)
);

BUFx8_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_19),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_188),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_20),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g236 ( 
.A1(n_161),
.A2(n_10),
.B(n_11),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_164),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

OAI21x1_ASAP7_75t_L g246 ( 
.A1(n_190),
.A2(n_12),
.B(n_13),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_198),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_160),
.Y(n_249)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_23),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

BUFx8_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_187),
.B(n_15),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_R g259 ( 
.A(n_218),
.B(n_171),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_224),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_253),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_253),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_249),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_172),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_R g270 ( 
.A(n_223),
.B(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

BUFx6f_ASAP7_75t_SL g275 ( 
.A(n_222),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_252),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_256),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_256),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_248),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_248),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_248),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_248),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_248),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_238),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_238),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_238),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_228),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_228),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_228),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_244),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_244),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_223),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_240),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_216),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_229),
.B(n_177),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_216),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_254),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_233),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_232),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_239),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_280),
.C(n_279),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_230),
.B(n_233),
.C(n_246),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_281),
.B(n_230),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_241),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_258),
.B(n_251),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_303),
.B(n_250),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_178),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_234),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_229),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

AO221x1_ASAP7_75t_L g328 ( 
.A1(n_274),
.A2(n_242),
.B1(n_246),
.B2(n_236),
.C(n_243),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_229),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_217),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_301),
.B(n_180),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_243),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_289),
.B(n_181),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_217),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_217),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_217),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_217),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_267),
.B(n_243),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_269),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_243),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_257),
.B(n_234),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_237),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_259),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_237),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_295),
.B(n_182),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_261),
.B(n_220),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_263),
.B(n_220),
.Y(n_350)
);

BUFx2_ASAP7_75t_R g351 ( 
.A(n_260),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_275),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_264),
.B(n_220),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_265),
.B(n_220),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_275),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_260),
.B(n_207),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_266),
.B(n_226),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_266),
.B(n_183),
.Y(n_359)
);

BUFx8_ASAP7_75t_L g360 ( 
.A(n_275),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_259),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_301),
.B(n_191),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_192),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_259),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_301),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_300),
.A2(n_227),
.B1(n_225),
.B2(n_208),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_194),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_346),
.B(n_361),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_306),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_311),
.B(n_196),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_365),
.B(n_197),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_310),
.B(n_200),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_310),
.B(n_202),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_340),
.B(n_203),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_206),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_327),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_322),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_209),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_221),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_213),
.Y(n_389)
);

BUFx4f_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_319),
.B(n_221),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_328),
.A2(n_236),
.B1(n_215),
.B2(n_17),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_28),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

NOR3xp33_ASAP7_75t_SL g396 ( 
.A(n_335),
.B(n_15),
.C(n_16),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_16),
.Y(n_397)
);

NAND2x1p5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_29),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_319),
.B(n_30),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_314),
.B(n_31),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_17),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_312),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_364),
.A2(n_98),
.B(n_34),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_371),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_336),
.B(n_37),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_309),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_323),
.A2(n_18),
.B1(n_39),
.B2(n_40),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_323),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_313),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_314),
.B(n_44),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_320),
.B(n_47),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_315),
.B(n_52),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_344),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_417)
);

AND3x1_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_358),
.C(n_320),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_360),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_321),
.A2(n_59),
.B1(n_63),
.B2(n_65),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_366),
.B(n_335),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_333),
.A2(n_362),
.B1(n_318),
.B2(n_331),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_362),
.Y(n_426)
);

BUFx8_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_SL g429 ( 
.A(n_359),
.B(n_348),
.C(n_332),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_349),
.B(n_67),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_326),
.B(n_68),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_350),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

AND3x2_ASAP7_75t_SL g438 ( 
.A(n_359),
.B(n_69),
.C(n_70),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_324),
.B(n_71),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_404),
.B(n_423),
.Y(n_441)
);

NOR2x1_ASAP7_75t_SL g442 ( 
.A(n_392),
.B(n_348),
.Y(n_442)
);

O2A1O1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_397),
.A2(n_401),
.B(n_420),
.C(n_407),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_373),
.Y(n_445)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_418),
.B(n_330),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_424),
.A2(n_339),
.B(n_338),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_391),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_337),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_72),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_414),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_372),
.B(n_79),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_430),
.B(n_80),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_432),
.B(n_81),
.Y(n_456)
);

O2A1O1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_388),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_88),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_375),
.A2(n_89),
.B(n_90),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_395),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_92),
.Y(n_462)
);

A2O1A1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_425),
.A2(n_93),
.B(n_94),
.C(n_95),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_97),
.C(n_100),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_400),
.A2(n_101),
.B(n_102),
.C(n_104),
.Y(n_465)
);

NAND2x1p5_ASAP7_75t_L g466 ( 
.A(n_390),
.B(n_107),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_108),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_391),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_433),
.A2(n_399),
.B1(n_415),
.B2(n_413),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_431),
.A2(n_379),
.B1(n_378),
.B2(n_414),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_109),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_110),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_435),
.A2(n_389),
.B(n_416),
.Y(n_475)
);

O2A1O1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_376),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_427),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_L g478 ( 
.A1(n_384),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_381),
.B(n_387),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_406),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_122),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_SL g482 ( 
.A1(n_411),
.A2(n_123),
.B(n_124),
.C(n_126),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_380),
.A2(n_434),
.B(n_386),
.Y(n_483)
);

OAI22x1_ASAP7_75t_L g484 ( 
.A1(n_437),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_390),
.B(n_412),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_410),
.B(n_132),
.Y(n_486)
);

INVx3_ASAP7_75t_SL g487 ( 
.A(n_419),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_383),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_393),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_490)
);

BUFx8_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_398),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_138),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_410),
.B(n_139),
.Y(n_494)
);

O2A1O1Ixp33_ASAP7_75t_SL g495 ( 
.A1(n_422),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_398),
.B(n_408),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

BUFx4f_ASAP7_75t_SL g498 ( 
.A(n_427),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_394),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_475),
.A2(n_403),
.B(n_405),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_405),
.B(n_422),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_471),
.A2(n_409),
.B(n_417),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_470),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_450),
.A2(n_417),
.B(n_402),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

INVx8_ASAP7_75t_L g507 ( 
.A(n_452),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_444),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_450),
.A2(n_394),
.B(n_438),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_394),
.Y(n_510)
);

OAI21x1_ASAP7_75t_SL g511 ( 
.A1(n_442),
.A2(n_396),
.B(n_145),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_460),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_451),
.A2(n_143),
.B(n_147),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_148),
.B(n_150),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_454),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_462),
.A2(n_152),
.B(n_153),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_443),
.B(n_154),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_458),
.A2(n_155),
.B(n_467),
.Y(n_520)
);

AOI22x1_ASAP7_75t_L g521 ( 
.A1(n_447),
.A2(n_496),
.B1(n_492),
.B2(n_469),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_479),
.A2(n_474),
.B(n_448),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_464),
.A2(n_473),
.B(n_462),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_463),
.A2(n_482),
.B(n_455),
.Y(n_524)
);

AO21x2_ASAP7_75t_L g525 ( 
.A1(n_456),
.A2(n_495),
.B(n_472),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g526 ( 
.A1(n_465),
.A2(n_481),
.B(n_459),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_460),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_480),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_466),
.Y(n_530)
);

AOI21x1_ASAP7_75t_L g531 ( 
.A1(n_441),
.A2(n_494),
.B(n_493),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_487),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_488),
.Y(n_534)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_457),
.A2(n_476),
.B(n_478),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_485),
.A2(n_489),
.B(n_486),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_468),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_499),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_453),
.A2(n_490),
.B(n_484),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_477),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_491),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_498),
.A2(n_471),
.B(n_475),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_475),
.A2(n_483),
.B(n_386),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_452),
.B(n_460),
.Y(n_547)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_547),
.B(n_506),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_542),
.A2(n_502),
.B1(n_519),
.B2(n_523),
.Y(n_550)
);

BUFx2_ASAP7_75t_R g551 ( 
.A(n_532),
.Y(n_551)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_514),
.A2(n_505),
.B(n_501),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_529),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_507),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_517),
.A2(n_503),
.B1(n_511),
.B2(n_541),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_516),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_534),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_532),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_546),
.A2(n_520),
.B(n_521),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_541),
.A2(n_517),
.B1(n_511),
.B2(n_535),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_536),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_504),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_539),
.A2(n_541),
.B1(n_540),
.B2(n_533),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_539),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_517),
.A2(n_503),
.B1(n_541),
.B2(n_505),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_507),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_533),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_507),
.Y(n_570)
);

INVx4_ASAP7_75t_SL g571 ( 
.A(n_547),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_543),
.A2(n_530),
.B1(n_508),
.B2(n_538),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_500),
.A2(n_501),
.B(n_531),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_507),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_540),
.B(n_536),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_547),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_522),
.A2(n_515),
.B(n_509),
.Y(n_578)
);

NOR2x1_ASAP7_75t_SL g579 ( 
.A(n_545),
.B(n_525),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_517),
.A2(n_535),
.B1(n_540),
.B2(n_530),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_545),
.A2(n_530),
.B1(n_543),
.B2(n_525),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_527),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_512),
.Y(n_586)
);

NAND2x1p5_ASAP7_75t_L g587 ( 
.A(n_509),
.B(n_515),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_528),
.Y(n_588)
);

AO21x1_ASAP7_75t_L g589 ( 
.A1(n_510),
.A2(n_526),
.B(n_524),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_554),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_512),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_564),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_580),
.A2(n_510),
.B1(n_513),
.B2(n_528),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_568),
.Y(n_595)
);

CKINVDCx11_ASAP7_75t_R g596 ( 
.A(n_583),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_563),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_584),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_585),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_585),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_588),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_512),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_549),
.B(n_545),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_559),
.B(n_518),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_566),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_SL g611 ( 
.A(n_568),
.B(n_525),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_582),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_559),
.B(n_518),
.Y(n_613)
);

NOR3xp33_ASAP7_75t_SL g614 ( 
.A(n_560),
.B(n_544),
.C(n_548),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_510),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_582),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_558),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_549),
.B(n_507),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_551),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_568),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_575),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_549),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_524),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_572),
.B(n_526),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_589),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_586),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_550),
.A2(n_504),
.B1(n_548),
.B2(n_567),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_586),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_577),
.B(n_562),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

AND2x4_ASAP7_75t_SL g633 ( 
.A(n_568),
.B(n_570),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_552),
.A2(n_557),
.B1(n_568),
.B2(n_570),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_571),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_608),
.B(n_587),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_609),
.B(n_579),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_609),
.B(n_579),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_613),
.B(n_587),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_626),
.B(n_587),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_591),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_598),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_622),
.B(n_571),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_613),
.B(n_552),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_602),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_602),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_622),
.B(n_571),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_615),
.B(n_578),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_603),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_603),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_617),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_625),
.B(n_578),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_623),
.B(n_560),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_615),
.B(n_631),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_631),
.B(n_578),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_590),
.B(n_571),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_627),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_606),
.B(n_556),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_596),
.B(n_620),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_601),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_591),
.Y(n_662)
);

AOI221xp5_ASAP7_75t_L g663 ( 
.A1(n_629),
.A2(n_556),
.B1(n_574),
.B2(n_570),
.C(n_573),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_573),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_599),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_600),
.Y(n_666)
);

NOR2x1_ASAP7_75t_L g667 ( 
.A(n_619),
.B(n_574),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_600),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_632),
.B(n_561),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_627),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_601),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_649),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_641),
.B(n_604),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_649),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_650),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_650),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_654),
.B(n_625),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_641),
.B(n_604),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_654),
.B(n_624),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_645),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_671),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_651),
.B(n_657),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_663),
.B(n_591),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_642),
.B(n_597),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_605),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_661),
.B(n_610),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_658),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_662),
.B(n_638),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_645),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_639),
.B(n_607),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_653),
.B(n_634),
.C(n_614),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_646),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_639),
.B(n_607),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_637),
.B(n_635),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_661),
.B(n_612),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_656),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_646),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_667),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_658),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_664),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_670),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_688),
.B(n_637),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_682),
.B(n_648),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_688),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_688),
.B(n_638),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_691),
.B(n_660),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_681),
.B(n_684),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_700),
.B(n_648),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_685),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_700),
.B(n_655),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_694),
.B(n_677),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_694),
.B(n_669),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_699),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_694),
.B(n_655),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_679),
.B(n_636),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_680),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_701),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_687),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_685),
.B(n_686),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_672),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_687),
.Y(n_721)
);

NAND4xp25_ASAP7_75t_L g722 ( 
.A(n_706),
.B(n_683),
.C(n_695),
.D(n_659),
.Y(n_722)
);

NAND2x1_ASAP7_75t_L g723 ( 
.A(n_704),
.B(n_718),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_718),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_707),
.B(n_592),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_719),
.A2(n_683),
.B(n_698),
.C(n_593),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_703),
.B(n_644),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_721),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_721),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_709),
.A2(n_678),
.B1(n_673),
.B2(n_696),
.Y(n_730)
);

NOR4xp25_ASAP7_75t_L g731 ( 
.A(n_713),
.B(n_698),
.C(n_676),
.D(n_675),
.Y(n_731)
);

AOI31xp33_ASAP7_75t_L g732 ( 
.A1(n_725),
.A2(n_711),
.A3(n_702),
.B(n_705),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_723),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_724),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_722),
.A2(n_720),
.B(n_717),
.C(n_715),
.Y(n_735)
);

AOI21xp33_ASAP7_75t_L g736 ( 
.A1(n_726),
.A2(n_685),
.B(n_678),
.Y(n_736)
);

AOI321xp33_ASAP7_75t_L g737 ( 
.A1(n_735),
.A2(n_731),
.A3(n_730),
.B1(n_729),
.B2(n_728),
.C(n_711),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_734),
.B(n_727),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_736),
.Y(n_739)
);

AOI211xp5_ASAP7_75t_SL g740 ( 
.A1(n_732),
.A2(n_704),
.B(n_678),
.C(n_673),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_733),
.Y(n_741)
);

AOI21xp33_ASAP7_75t_L g742 ( 
.A1(n_733),
.A2(n_673),
.B(n_640),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_702),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_738),
.B(n_596),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_742),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_737),
.B(n_741),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_741),
.B1(n_704),
.B2(n_712),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_746),
.A2(n_743),
.B1(n_716),
.B2(n_674),
.C(n_692),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_716),
.B1(n_689),
.B2(n_697),
.C(n_705),
.Y(n_749)
);

NAND5xp2_ASAP7_75t_L g750 ( 
.A(n_746),
.B(n_618),
.C(n_690),
.D(n_693),
.E(n_714),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_748),
.A2(n_656),
.B1(n_712),
.B2(n_647),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_749),
.A2(n_656),
.B1(n_712),
.B2(n_647),
.Y(n_752)
);

NOR2x1p5_ASAP7_75t_L g753 ( 
.A(n_750),
.B(n_570),
.Y(n_753)
);

OAI211xp5_ASAP7_75t_SL g754 ( 
.A1(n_748),
.A2(n_667),
.B(n_636),
.C(n_644),
.Y(n_754)
);

AO22x2_ASAP7_75t_L g755 ( 
.A1(n_750),
.A2(n_670),
.B1(n_714),
.B2(n_680),
.Y(n_755)
);

NOR2x1_ASAP7_75t_L g756 ( 
.A(n_750),
.B(n_570),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_750),
.B(n_708),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_SL g758 ( 
.A(n_751),
.B(n_611),
.C(n_616),
.Y(n_758)
);

AOI211xp5_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_621),
.B(n_611),
.C(n_628),
.Y(n_759)
);

NAND2x1_ASAP7_75t_L g760 ( 
.A(n_756),
.B(n_647),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_753),
.B(n_757),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_755),
.B(n_708),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_752),
.B(n_710),
.Y(n_763)
);

OAI221xp5_ASAP7_75t_L g764 ( 
.A1(n_756),
.A2(n_595),
.B1(n_640),
.B2(n_621),
.C(n_652),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_758),
.A2(n_643),
.B1(n_607),
.B2(n_621),
.C(n_710),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_760),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_762),
.Y(n_768)
);

CKINVDCx6p67_ASAP7_75t_R g769 ( 
.A(n_763),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_765),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_767),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_764),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_769),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_766),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_773),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_771),
.B(n_759),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_772),
.A2(n_595),
.B1(n_633),
.B2(n_621),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_770),
.Y(n_778)
);

AOI22x1_ASAP7_75t_L g779 ( 
.A1(n_775),
.A2(n_774),
.B1(n_574),
.B2(n_621),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_778),
.A2(n_595),
.B1(n_633),
.B2(n_643),
.Y(n_780)
);

XNOR2xp5_ASAP7_75t_L g781 ( 
.A(n_779),
.B(n_776),
.Y(n_781)
);

AOI21xp33_ASAP7_75t_SL g782 ( 
.A1(n_781),
.A2(n_777),
.B(n_780),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_782),
.A2(n_619),
.B1(n_630),
.B2(n_643),
.Y(n_783)
);

XNOR2xp5_ASAP7_75t_L g784 ( 
.A(n_783),
.B(n_619),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_784),
.A2(n_668),
.B1(n_666),
.B2(n_665),
.Y(n_785)
);


endmodule