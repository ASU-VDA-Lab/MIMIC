module real_jpeg_13552_n_12 (n_5, n_4, n_8, n_0, n_261, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_261;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_2),
.A2(n_44),
.B1(n_62),
.B2(n_63),
.Y(n_122)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_28),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_28),
.B1(n_62),
.B2(n_63),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_6),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_100),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_6),
.B(n_25),
.C(n_38),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_6),
.B(n_29),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_37),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_63),
.B(n_73),
.C(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_59),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_68),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_68),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_33),
.B1(n_55),
.B2(n_56),
.Y(n_105)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_126),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_125),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_106),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_16),
.B(n_106),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.C(n_89),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_19),
.B(n_50),
.C(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_20),
.B(n_35),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_21),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_23),
.A2(n_30),
.B(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_23),
.B(n_34),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_25),
.B(n_157),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_28),
.A2(n_41),
.B(n_74),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_28),
.B(n_60),
.C(n_63),
.Y(n_211)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_32),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_30),
.B(n_137),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_30),
.A2(n_31),
.B(n_92),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_31),
.B(n_169),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_34),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_34),
.B(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B(n_45),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_36),
.A2(n_86),
.B(n_98),
.Y(n_224)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_37),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_37),
.B(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_37),
.B(n_142),
.Y(n_152)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_42),
.B(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_45),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_45),
.B(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_46),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_69),
.B2(n_70),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_64),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_54),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_54),
.B(n_115),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_55),
.B(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_67),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_59),
.B(n_105),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_63),
.B1(n_73),
.B2(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_64),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_71),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_75),
.B(n_79),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_77),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_81),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_79),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_81),
.B(n_100),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_82),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_84),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_83),
.A2(n_84),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_84),
.B(n_181),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_89),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.C(n_101),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_90),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_91),
.B(n_95),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_94),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_94),
.B(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_99),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_103),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_121),
.B(n_124),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_120),
.B(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_123),
.B(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_252),
.B(n_257),
.Y(n_126)
);

AOI321xp33_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_226),
.A3(n_245),
.B1(n_250),
.B2(n_251),
.C(n_261),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_202),
.B(n_225),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_185),
.B(n_201),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_172),
.B(n_184),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_153),
.B(n_171),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_147),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_147),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_146),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_144),
.C(n_146),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_165),
.B(n_170),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_161),
.B(n_164),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_168),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_174),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_200),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_200),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_192),
.B1(n_193),
.B2(n_199),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.C(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_193),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.CI(n_196),
.CON(n_193),
.SN(n_193)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.C(n_196),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_204),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_214),
.B2(n_215),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_208),
.C(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_221),
.C(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_240),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_240),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_236),
.C(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_234),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_231),
.CI(n_234),
.CON(n_242),
.SN(n_242)
);

NAND2x1_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_242),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_249),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);


endmodule