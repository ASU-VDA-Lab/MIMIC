module fake_jpeg_23659_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_39),
.Y(n_53)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_30),
.B1(n_28),
.B2(n_23),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_49),
.B1(n_54),
.B2(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_28),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_55),
.Y(n_76)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_29),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_24),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_26),
.C(n_18),
.Y(n_80)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_23),
.B1(n_19),
.B2(n_32),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_70),
.B1(n_78),
.B2(n_54),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_18),
.C(n_17),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_79),
.B(n_29),
.Y(n_110)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_22),
.B(n_19),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_71),
.C(n_84),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_48),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_44),
.B1(n_48),
.B2(n_58),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_92),
.B1(n_95),
.B2(n_108),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_48),
.B1(n_58),
.B2(n_50),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_48),
.B1(n_58),
.B2(n_50),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_54),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_31),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_102),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_10),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_26),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_109),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_46),
.C(n_38),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_51),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_52),
.B1(n_46),
.B2(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_42),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_29),
.B(n_31),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_83),
.B1(n_77),
.B2(n_75),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_117),
.B1(n_119),
.B2(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_66),
.B1(n_46),
.B2(n_91),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_126),
.B(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_52),
.B1(n_42),
.B2(n_57),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_84),
.B1(n_71),
.B2(n_74),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_96),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_132),
.C(n_108),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_29),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_46),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_36),
.C(n_40),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_73),
.B1(n_72),
.B2(n_11),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_40),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_98),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_147),
.C(n_151),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_96),
.A3(n_95),
.B1(n_102),
.B2(n_98),
.C(n_36),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_101),
.C(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_101),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_27),
.B(n_1),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_88),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_88),
.B1(n_104),
.B2(n_38),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_160),
.B1(n_114),
.B2(n_113),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_122),
.C(n_29),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_104),
.B1(n_31),
.B2(n_27),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_29),
.C(n_27),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_8),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_176),
.B1(n_185),
.B2(n_7),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_165),
.B(n_0),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_125),
.B1(n_120),
.B2(n_134),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_173),
.B1(n_178),
.B2(n_0),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_4),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_115),
.B(n_136),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_171),
.B(n_179),
.Y(n_198)
);

AOI22x1_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_140),
.B1(n_151),
.B2(n_136),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_122),
.B1(n_132),
.B2(n_115),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_0),
.C(n_2),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_150),
.B1(n_146),
.B2(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_143),
.B1(n_137),
.B2(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_139),
.B1(n_144),
.B2(n_145),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_158),
.A3(n_157),
.B1(n_160),
.B2(n_159),
.C1(n_27),
.C2(n_153),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_200),
.A3(n_202),
.B1(n_187),
.B2(n_203),
.C1(n_190),
.C2(n_196),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_27),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_196),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_190),
.C(n_193),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_197),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_8),
.C(n_14),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_204),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_174),
.C(n_167),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_202),
.C(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_176),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_15),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_181),
.B1(n_182),
.B2(n_177),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_3),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_185),
.B(n_170),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_207),
.A2(n_211),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_169),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_179),
.B(n_184),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_217),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_216),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_195),
.B(n_193),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_207),
.B(n_208),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_209),
.B1(n_211),
.B2(n_215),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_7),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_9),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_229),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_9),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_9),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_213),
.C(n_218),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_233),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_225),
.B(n_229),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_207),
.C(n_11),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_10),
.B(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_15),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_13),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_224),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_14),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_234),
.B(n_237),
.C(n_15),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_250),
.B(n_240),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_250),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_251),
.B(n_255),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_242),
.Y(n_257)
);


endmodule