module real_jpeg_4456_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_0),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_0),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_1),
.Y(n_134)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_1),
.Y(n_350)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_1),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_2),
.A2(n_49),
.B1(n_250),
.B2(n_332),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_2),
.A2(n_49),
.B1(n_309),
.B2(n_409),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_2),
.A2(n_49),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_3),
.Y(n_528)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_4),
.Y(n_352)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_4),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_5),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_5),
.A2(n_56),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_5),
.A2(n_56),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_5),
.A2(n_56),
.B1(n_412),
.B2(n_414),
.Y(n_411)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_6),
.Y(n_525)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_9),
.A2(n_144),
.B1(n_145),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_9),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_9),
.A2(n_113),
.B1(n_144),
.B2(n_297),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_9),
.A2(n_144),
.B1(n_275),
.B2(n_392),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_9),
.A2(n_144),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_10),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_12),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_87),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_12),
.A2(n_87),
.B1(n_223),
.B2(n_242),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_12),
.A2(n_87),
.B1(n_306),
.B2(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_13),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_13),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_13),
.A2(n_186),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_13),
.A2(n_39),
.B1(n_186),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_13),
.A2(n_186),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_14),
.A2(n_201),
.B1(n_207),
.B2(n_208),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_14),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_14),
.A2(n_120),
.B1(n_207),
.B2(n_274),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_14),
.A2(n_207),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_14),
.A2(n_53),
.B1(n_147),
.B2(n_207),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_15),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_15),
.A2(n_201),
.B1(n_230),
.B2(n_250),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_15),
.A2(n_65),
.B1(n_230),
.B2(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_15),
.A2(n_54),
.B1(n_133),
.B2(n_230),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_16),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_16),
.A2(n_94),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_16),
.A2(n_94),
.B1(n_115),
.B2(n_242),
.Y(n_406)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_18),
.A2(n_123),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_18),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_18),
.B(n_194),
.C(n_197),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_18),
.B(n_73),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_18),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_18),
.B(n_118),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_18),
.B(n_288),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_523),
.B(n_526),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_165),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_163),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_135),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_23),
.B(n_135),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_124),
.B2(n_125),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_57),
.C(n_95),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_26),
.B(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_27),
.A2(n_43),
.B1(n_50),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_27),
.A2(n_380),
.B(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_27),
.A2(n_50),
.B1(n_426),
.B2(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_28),
.A2(n_378),
.B(n_379),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_28),
.B(n_381),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_36)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_38),
.Y(n_285)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_38),
.Y(n_292)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_40),
.Y(n_421)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_50),
.B(n_179),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_50),
.A2(n_445),
.B(n_467),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_51),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_51),
.B(n_143),
.Y(n_466)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_57),
.A2(n_95),
.B1(n_96),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_57)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_58),
.A2(n_81),
.B1(n_88),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_58),
.A2(n_88),
.B1(n_323),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_58),
.A2(n_88),
.B1(n_419),
.B2(n_422),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g302 ( 
.A1(n_60),
.A2(n_287),
.A3(n_303),
.B1(n_306),
.B2(n_308),
.Y(n_302)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_69),
.Y(n_312)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

AOI22x1_ASAP7_75t_L g446 ( 
.A1(n_73),
.A2(n_127),
.B1(n_327),
.B2(n_447),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_73),
.A2(n_127),
.B1(n_156),
.B2(n_455),
.Y(n_454)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_77),
.Y(n_233)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_77),
.Y(n_278)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_82),
.Y(n_389)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_88),
.B(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_88),
.A2(n_323),
.B(n_326),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_141),
.C(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_95),
.A2(n_96),
.B1(n_153),
.B2(n_154),
.Y(n_512)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_117),
.B(n_119),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_97),
.A2(n_175),
.B(n_180),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_97),
.A2(n_117),
.B1(n_227),
.B2(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_97),
.A2(n_180),
.B(n_273),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_97),
.A2(n_117),
.B1(n_391),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_98),
.B(n_181),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_98),
.A2(n_118),
.B1(n_408),
.B2(n_411),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_98),
.A2(n_118),
.B1(n_411),
.B2(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_98),
.A2(n_118),
.B1(n_430),
.B2(n_458),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_109),
.Y(n_310)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_110),
.A2(n_227),
.B(n_234),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_117),
.A2(n_234),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_118),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_119),
.Y(n_458)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_122),
.Y(n_392)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_122),
.Y(n_416)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_127),
.A2(n_281),
.B(n_289),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_127),
.B(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_127),
.A2(n_289),
.B(n_480),
.Y(n_479)
);

OAI21xp33_ASAP7_75t_SL g378 ( 
.A1(n_132),
.A2(n_179),
.B(n_359),
.Y(n_378)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.C(n_151),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_518)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_140),
.A2(n_141),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_151),
.A2(n_152),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_159),
.Y(n_388)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_506),
.B(n_520),
.Y(n_166)
);

OAI311xp33_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_395),
.A3(n_482),
.B1(n_500),
.C1(n_501),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_337),
.B(n_394),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_314),
.B(n_336),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_267),
.B(n_313),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_237),
.B(n_266),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_198),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_173),
.B(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_189),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_174),
.A2(n_189),
.B1(n_190),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_178),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_211),
.B(n_217),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g281 ( 
.A1(n_179),
.A2(n_282),
.B(n_286),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_179),
.B(n_349),
.Y(n_359)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_185),
.Y(n_433)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_224),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_199),
.B(n_225),
.C(n_236),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_211),
.B(n_217),
.Y(n_199)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_200),
.Y(n_262)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_211),
.A2(n_362),
.B1(n_363),
.B2(n_366),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_211),
.A2(n_401),
.B1(n_402),
.B2(n_406),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_211),
.A2(n_404),
.B(n_406),
.Y(n_434)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_221),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_212),
.A2(n_255),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_212),
.A2(n_296),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_212),
.A2(n_367),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_220),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_220),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_235),
.B2(n_236),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_259),
.B(n_265),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_247),
.B(n_258),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_243),
.Y(n_371)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_257),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_254),
.B(n_256),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_252),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_256),
.A2(n_295),
.B(n_300),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_263),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_269),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_293),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_279),
.B2(n_280),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_279),
.C(n_293),
.Y(n_315)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_277),
.Y(n_410)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_282),
.Y(n_423)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_302),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx4_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_315),
.B(n_316),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_321),
.B2(n_335),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_320),
.C(n_335),
.Y(n_338)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_328),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_329),
.C(n_330),
.Y(n_372)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_338),
.B(n_339),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_375),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_340)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_360),
.B2(n_361),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_343),
.B(n_360),
.Y(n_478)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_347),
.A3(n_351),
.B1(n_353),
.B2(n_359),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_372),
.B(n_373),
.C(n_375),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_385),
.B2(n_393),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_376),
.B(n_386),
.C(n_390),
.Y(n_491)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_390),
.Y(n_385)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

INVx11_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_468),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_SL g501 ( 
.A1(n_396),
.A2(n_468),
.B(n_502),
.C(n_505),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_448),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_397),
.B(n_448),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_427),
.C(n_436),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_398),
.B(n_427),
.CI(n_436),
.CON(n_481),
.SN(n_481)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_417),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_418),
.C(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_407),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_400),
.B(n_407),
.Y(n_474)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx8_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

INVx8_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.Y(n_417)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_419),
.Y(n_447)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_434),
.B2(n_435),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_434),
.Y(n_462)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_434),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_434),
.A2(n_435),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_434),
.A2(n_462),
.B(n_465),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_443),
.C(n_446),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_438),
.B(n_440),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_443),
.A2(n_444),
.B1(n_446),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_449),
.B(n_452),
.C(n_460),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_460),
.B2(n_461),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_456),
.B(n_459),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_457),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_459),
.B(n_511),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_459),
.B(n_509),
.C(n_511),
.Y(n_519)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_481),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_481),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_474),
.C(n_475),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_471),
.B1(n_474),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.C(n_479),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_476),
.A2(n_477),
.B1(n_479),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_479),
.Y(n_488)
);

BUFx24_ASAP7_75t_SL g530 ( 
.A(n_481),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_495),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_503),
.B(n_504),
.Y(n_502)
);

NOR2x1_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_492),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_492),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.C(n_491),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_498),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_490),
.B1(n_491),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_491),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_497),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_497),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_515),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_508),
.B(n_514),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_514),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_510),
.Y(n_508)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_512),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_515),
.A2(n_521),
.B(n_522),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_519),
.Y(n_522)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_524),
.Y(n_527)
);

INVx13_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_528),
.Y(n_526)
);


endmodule