module fake_jpeg_3711_n_656 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_656);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_656;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_612;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_58),
.Y(n_191)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_59),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_10),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_71),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_83),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_100),
.Y(n_137)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_92),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_95),
.Y(n_194)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_96),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_23),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_99),
.B(n_15),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_29),
.B(n_10),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_35),
.Y(n_108)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_33),
.Y(n_111)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_41),
.B(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_118),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_55),
.A2(n_11),
.B1(n_18),
.B2(n_17),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_23),
.B1(n_48),
.B2(n_46),
.Y(n_131)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_40),
.B(n_11),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_40),
.B(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_124),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_32),
.Y(n_123)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_47),
.B(n_8),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_131),
.A2(n_172),
.B1(n_175),
.B2(n_181),
.Y(n_297)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_60),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_142),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_61),
.B(n_48),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_146),
.B(n_161),
.Y(n_250)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_147),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_30),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_152),
.B(n_169),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_73),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_79),
.A2(n_30),
.B1(n_50),
.B2(n_31),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_162),
.A2(n_199),
.B1(n_200),
.B2(n_215),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_44),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_46),
.B1(n_39),
.B2(n_52),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_129),
.A2(n_50),
.B1(n_39),
.B2(n_22),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_123),
.A2(n_50),
.B1(n_71),
.B2(n_88),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_78),
.B(n_13),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_86),
.B(n_101),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_89),
.A2(n_13),
.B(n_19),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_192),
.B(n_3),
.Y(n_273)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_90),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_65),
.A2(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_91),
.B(n_7),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_92),
.Y(n_211)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_81),
.B(n_7),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_84),
.A2(n_70),
.B1(n_69),
.B2(n_72),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_217),
.A2(n_200),
.B1(n_192),
.B2(n_220),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_222),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_93),
.A2(n_8),
.B1(n_17),
.B2(n_15),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_220),
.A2(n_226),
.B1(n_152),
.B2(n_169),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_110),
.B(n_12),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_81),
.B(n_12),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_223),
.B(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_115),
.Y(n_225)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_109),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_231),
.Y(n_315)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_175),
.A2(n_77),
.B1(n_181),
.B2(n_149),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_235),
.A2(n_268),
.B1(n_284),
.B2(n_309),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_145),
.A2(n_95),
.B1(n_122),
.B2(n_119),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_237),
.A2(n_240),
.B1(n_244),
.B2(n_252),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_238),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_152),
.A2(n_130),
.B1(n_107),
.B2(n_14),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_241),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_145),
.A2(n_97),
.B(n_18),
.C(n_15),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_242),
.B(n_288),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_148),
.B(n_97),
.C(n_18),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_245),
.B(n_307),
.C(n_229),
.Y(n_314)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_246),
.Y(n_327)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_159),
.Y(n_247)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_249),
.Y(n_373)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_162),
.A2(n_156),
.B1(n_153),
.B2(n_206),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

BUFx4f_ASAP7_75t_L g362 ( 
.A(n_255),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_133),
.B(n_2),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_256),
.B(n_280),
.Y(n_328)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_140),
.Y(n_257)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_257),
.Y(n_344)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_258),
.Y(n_359)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_151),
.Y(n_267)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_198),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_268)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_269),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_165),
.Y(n_270)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_165),
.Y(n_271)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_271),
.Y(n_342)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_273),
.B(n_274),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_133),
.B(n_3),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_170),
.Y(n_276)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_177),
.Y(n_277)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_277),
.Y(n_370)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_150),
.Y(n_278)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_278),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_279),
.A2(n_244),
.B1(n_252),
.B2(n_302),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_180),
.B(n_5),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_137),
.B(n_5),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_283),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_180),
.A2(n_5),
.B1(n_208),
.B2(n_137),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_282),
.A2(n_304),
.B(n_279),
.Y(n_367)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_168),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_285),
.B(n_289),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_138),
.A2(n_158),
.B1(n_221),
.B2(n_218),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_286),
.A2(n_287),
.B1(n_294),
.B2(n_312),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_191),
.A2(n_143),
.B1(n_202),
.B2(n_182),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_182),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_168),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_290),
.Y(n_316)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_292),
.Y(n_348)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_160),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_295),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_223),
.A2(n_201),
.B1(n_136),
.B2(n_210),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_135),
.B(n_144),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_141),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_298),
.Y(n_364)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_178),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_170),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_301),
.Y(n_368)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_174),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_303),
.B(n_305),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_147),
.A2(n_194),
.B1(n_205),
.B2(n_227),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_164),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_196),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_306),
.B(n_308),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_166),
.B(n_187),
.C(n_194),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_134),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_217),
.A2(n_134),
.B1(n_189),
.B2(n_209),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_228),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_310),
.Y(n_357)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_189),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_243),
.B(n_209),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_313),
.B(n_322),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_247),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_226),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_317),
.B(n_326),
.C(n_337),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_239),
.B(n_171),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_229),
.B(n_179),
.C(n_171),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_281),
.A2(n_139),
.B(n_179),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_332),
.A2(n_354),
.B(n_371),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_139),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_242),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_139),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_250),
.B(n_245),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_358),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_265),
.A2(n_294),
.B(n_240),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_254),
.A2(n_302),
.B1(n_235),
.B2(n_297),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_356),
.A2(n_362),
.B1(n_358),
.B2(n_346),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_295),
.B(n_307),
.Y(n_358)
);

AOI32xp33_ASAP7_75t_L g360 ( 
.A1(n_297),
.A2(n_259),
.A3(n_236),
.B1(n_263),
.B2(n_266),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_257),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_367),
.B(n_350),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_297),
.B(n_234),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_369),
.B(n_337),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_268),
.B1(n_262),
.B2(n_267),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_309),
.B1(n_304),
.B2(n_287),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_374),
.A2(n_378),
.B1(n_394),
.B2(n_401),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_348),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_375),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_377),
.Y(n_452)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_311),
.C(n_230),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_379),
.B(n_380),
.C(n_383),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_314),
.B(n_271),
.C(n_270),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_276),
.B1(n_299),
.B2(n_296),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_384),
.A2(n_385),
.B1(n_390),
.B2(n_412),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_290),
.B1(n_233),
.B2(n_241),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_286),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_405),
.Y(n_428)
);

OA21x2_ASAP7_75t_SL g389 ( 
.A1(n_339),
.A2(n_249),
.B(n_238),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_403),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_333),
.A2(n_298),
.B1(n_306),
.B2(n_260),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_362),
.A2(n_338),
.B1(n_349),
.B2(n_313),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_392),
.A2(n_365),
.B1(n_343),
.B2(n_321),
.Y(n_424)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_338),
.A2(n_249),
.B1(n_269),
.B2(n_322),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_336),
.A2(n_317),
.B(n_367),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_373),
.B(n_321),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_397),
.A2(n_399),
.B(n_400),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_398),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_326),
.B1(n_332),
.B2(n_341),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_363),
.A2(n_329),
.B1(n_370),
.B2(n_352),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_411),
.B1(n_420),
.B2(n_391),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_324),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_328),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_393),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g410 ( 
.A(n_363),
.B(n_353),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_325),
.A2(n_357),
.B1(n_316),
.B2(n_364),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_318),
.A2(n_342),
.B1(n_361),
.B2(n_344),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_368),
.A2(n_318),
.B1(n_361),
.B2(n_342),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_413),
.A2(n_365),
.B1(n_335),
.B2(n_331),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_315),
.B(n_319),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_417),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_315),
.B(n_319),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_415),
.B(n_418),
.Y(n_443)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_419),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_327),
.B(n_330),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_334),
.B(n_359),
.C(n_330),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_334),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_347),
.A2(n_320),
.B1(n_327),
.B2(n_359),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_335),
.Y(n_421)
);

OAI21xp33_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_345),
.B(n_320),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_421),
.Y(n_422)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_424),
.A2(n_427),
.B(n_449),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_414),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_431),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_399),
.A2(n_331),
.B(n_345),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_435),
.B(n_420),
.Y(n_479)
);

OAI21xp33_ASAP7_75t_L g440 ( 
.A1(n_396),
.A2(n_323),
.B(n_386),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_440),
.A2(n_454),
.B(n_459),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_417),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_456),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_376),
.B(n_323),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_445),
.C(n_410),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_376),
.B(n_386),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_377),
.A2(n_388),
.B(n_382),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_385),
.B(n_382),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_455),
.B(n_402),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_401),
.A2(n_394),
.B(n_411),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_374),
.A2(n_409),
.B1(n_406),
.B2(n_375),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_421),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_458),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_379),
.B(n_410),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_383),
.A2(n_408),
.B(n_404),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_462),
.Y(n_488)
);

INVx3_ASAP7_75t_SL g464 ( 
.A(n_432),
.Y(n_464)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_464),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_383),
.C(n_408),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_465),
.B(n_491),
.C(n_498),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_467),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_460),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_423),
.A2(n_384),
.B1(n_378),
.B2(n_390),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_468),
.A2(n_477),
.B1(n_439),
.B2(n_499),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_473),
.Y(n_527)
);

OAI32xp33_ASAP7_75t_L g474 ( 
.A1(n_461),
.A2(n_429),
.A3(n_458),
.B1(n_433),
.B2(n_452),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_423),
.A2(n_380),
.B1(n_405),
.B2(n_395),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_475),
.A2(n_477),
.B1(n_487),
.B2(n_490),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_476),
.A2(n_484),
.B(n_492),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_423),
.A2(n_403),
.B1(n_387),
.B2(n_381),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_426),
.Y(n_478)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_445),
.B(n_442),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_481),
.Y(n_525)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_482),
.Y(n_535)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_483),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_452),
.A2(n_407),
.B1(n_398),
.B2(n_416),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_436),
.Y(n_485)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_455),
.A2(n_412),
.B1(n_407),
.B2(n_415),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_486),
.A2(n_499),
.B1(n_468),
.B2(n_492),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_431),
.A2(n_418),
.B1(n_454),
.B2(n_430),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_489),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_460),
.B(n_438),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_450),
.A2(n_453),
.B1(n_427),
.B2(n_440),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_428),
.B(n_446),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_434),
.A2(n_449),
.B(n_431),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_428),
.B(n_446),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_493),
.B(n_497),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_460),
.B(n_450),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_494),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_434),
.A2(n_431),
.B(n_453),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_495),
.A2(n_496),
.B(n_425),
.Y(n_520)
);

OAI32xp33_ASAP7_75t_L g496 ( 
.A1(n_428),
.A2(n_446),
.A3(n_438),
.B1(n_431),
.B2(n_457),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_428),
.B(n_443),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_443),
.B(n_444),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_457),
.A2(n_424),
.B1(n_456),
.B2(n_439),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_422),
.C(n_462),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_505),
.B(n_523),
.C(n_497),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_466),
.B(n_447),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_508),
.B(n_516),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_509),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_447),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_510),
.B(n_518),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_511),
.A2(n_524),
.B1(n_536),
.B2(n_521),
.Y(n_554)
);

AO21x2_ASAP7_75t_SL g512 ( 
.A1(n_469),
.A2(n_495),
.B(n_496),
.Y(n_512)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_512),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_488),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_513),
.B(n_526),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_464),
.Y(n_515)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_432),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_448),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

XNOR2x1_ASAP7_75t_L g549 ( 
.A(n_520),
.B(n_521),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_486),
.A2(n_448),
.B1(n_451),
.B2(n_441),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_451),
.C(n_437),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_487),
.A2(n_435),
.B1(n_437),
.B2(n_432),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_480),
.B(n_475),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_481),
.A2(n_484),
.B1(n_469),
.B2(n_470),
.Y(n_529)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_529),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_500),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_530),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_497),
.B(n_498),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_531),
.B(n_502),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_470),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_532),
.B(n_514),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_489),
.Y(n_539)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_539),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_509),
.Y(n_574)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_527),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_556),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_517),
.B(n_498),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_545),
.B(n_548),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_503),
.B(n_471),
.C(n_500),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_553),
.C(n_555),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_511),
.A2(n_467),
.B1(n_476),
.B2(n_463),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_547),
.A2(n_563),
.B1(n_501),
.B2(n_528),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_517),
.B(n_471),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_518),
.B(n_474),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g577 ( 
.A(n_550),
.B(n_562),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_534),
.B(n_478),
.Y(n_551)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_551),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_503),
.B(n_472),
.C(n_482),
.Y(n_553)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_554),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_505),
.B(n_472),
.C(n_483),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_SL g556 ( 
.A(n_506),
.B(n_512),
.C(n_534),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_464),
.C(n_523),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_558),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_502),
.B(n_531),
.C(n_507),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_544),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_560),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_520),
.A2(n_536),
.B1(n_512),
.B2(n_524),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_564),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_539),
.B(n_522),
.Y(n_567)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_567),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_506),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_568),
.B(n_575),
.Y(n_592)
);

XOR2x1_ASAP7_75t_SL g571 ( 
.A(n_562),
.B(n_530),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_574),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_522),
.Y(n_572)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_572),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_504),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_563),
.A2(n_557),
.B1(n_547),
.B2(n_552),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_578),
.A2(n_579),
.B1(n_576),
.B2(n_566),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_537),
.A2(n_504),
.B(n_512),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_580),
.A2(n_587),
.B(n_567),
.Y(n_602)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_582),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_561),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_588),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_586),
.B(n_555),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_549),
.A2(n_530),
.B(n_509),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_584),
.B(n_558),
.C(n_541),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_589),
.B(n_596),
.C(n_598),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_593),
.B(n_601),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_579),
.A2(n_552),
.B1(n_538),
.B2(n_542),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_594),
.A2(n_595),
.B1(n_572),
.B2(n_605),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_574),
.B(n_559),
.C(n_544),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_554),
.C(n_550),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g600 ( 
.A(n_571),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_600),
.B(n_575),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_573),
.B(n_549),
.Y(n_601)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_602),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_573),
.B(n_565),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_603),
.B(n_604),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_583),
.B(n_535),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_568),
.B(n_542),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_605),
.B(n_587),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_580),
.A2(n_556),
.B(n_565),
.Y(n_607)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_607),
.Y(n_609)
);

A2O1A1Ixp33_ASAP7_75t_SL g631 ( 
.A1(n_611),
.A2(n_577),
.B(n_590),
.C(n_600),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_SL g634 ( 
.A(n_612),
.B(n_577),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_607),
.A2(n_569),
.B1(n_599),
.B2(n_597),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_614),
.B(n_616),
.Y(n_628)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_591),
.Y(n_615)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_615),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_589),
.B(n_578),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_597),
.B(n_593),
.Y(n_617)
);

NOR2x1_ASAP7_75t_L g627 ( 
.A(n_617),
.B(n_619),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_597),
.B(n_585),
.Y(n_619)
);

BUFx24_ASAP7_75t_SL g620 ( 
.A(n_592),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_620),
.B(n_622),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_570),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_621),
.B(n_596),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_606),
.A2(n_566),
.B1(n_576),
.B2(n_582),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_623),
.B(n_600),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_614),
.A2(n_602),
.B(n_598),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_625),
.A2(n_629),
.B(n_633),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_626),
.A2(n_630),
.B(n_628),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_618),
.B(n_594),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_590),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_SL g637 ( 
.A(n_631),
.B(n_634),
.Y(n_637)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_632),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_613),
.B(n_585),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_627),
.B(n_610),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_636),
.B(n_639),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_621),
.Y(n_638)
);

AOI21xp33_ASAP7_75t_L g648 ( 
.A1(n_638),
.A2(n_631),
.B(n_612),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_L g640 ( 
.A(n_624),
.B(n_608),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_640),
.A2(n_635),
.B(n_609),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_635),
.B(n_616),
.C(n_608),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_623),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_644),
.B(n_645),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_642),
.B(n_641),
.Y(n_645)
);

OAI211xp5_ASAP7_75t_L g649 ( 
.A1(n_646),
.A2(n_648),
.B(n_640),
.C(n_637),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_649),
.B(n_651),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_647),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_650),
.C(n_581),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_653),
.A2(n_581),
.B(n_519),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_654),
.B(n_515),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_655),
.A2(n_533),
.B(n_645),
.Y(n_656)
);


endmodule