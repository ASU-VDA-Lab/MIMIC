module fake_jpeg_2507_n_676 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_676);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_676;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_75),
.Y(n_137)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g153 ( 
.A(n_65),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_10),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_87),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_71),
.Y(n_169)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_74),
.B(n_49),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_80),
.Y(n_141)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_33),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_0),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_79),
.B(n_67),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_82),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_21),
.B(n_10),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_84),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_85),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_86),
.B(n_91),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_10),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_89),
.Y(n_227)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_41),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_92),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_36),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_104),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_98),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_101),
.A2(n_130),
.B1(n_26),
.B2(n_27),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_25),
.B(n_12),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_115),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_25),
.B(n_12),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_27),
.Y(n_148)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g110 ( 
.A(n_44),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_110),
.Y(n_229)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_44),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_39),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_13),
.B1(n_1),
.B2(n_3),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_37),
.Y(n_131)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_49),
.B1(n_37),
.B2(n_56),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_134),
.A2(n_152),
.B1(n_155),
.B2(n_162),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_148),
.B(n_186),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_150),
.B(n_17),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_85),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_152)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_79),
.B(n_52),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_154),
.B(n_161),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_74),
.A2(n_57),
.B1(n_52),
.B2(n_50),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_158),
.A2(n_173),
.B1(n_210),
.B2(n_220),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_79),
.A2(n_26),
.B1(n_51),
.B2(n_48),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_57),
.B1(n_22),
.B2(n_47),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_96),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_176),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_177),
.B(n_113),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_100),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_178),
.B(n_193),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_111),
.A2(n_52),
.B1(n_50),
.B2(n_47),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_183),
.A2(n_211),
.B1(n_120),
.B2(n_114),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_84),
.B(n_39),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_88),
.B(n_46),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_61),
.Y(n_194)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_89),
.B(n_43),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_195),
.B(n_196),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_72),
.B(n_43),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_68),
.Y(n_199)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_67),
.B(n_34),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_216),
.Y(n_257)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_60),
.A2(n_34),
.B1(n_32),
.B2(n_50),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_62),
.A2(n_132),
.B1(n_128),
.B2(n_121),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_100),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_215),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_64),
.B(n_22),
.Y(n_216)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_71),
.A2(n_47),
.B1(n_22),
.B2(n_35),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_117),
.B(n_14),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_221),
.B(n_19),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_73),
.A2(n_35),
.B1(n_3),
.B2(n_5),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_223),
.A2(n_226),
.B1(n_146),
.B2(n_175),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_126),
.A2(n_35),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_225),
.A2(n_119),
.B1(n_112),
.B2(n_98),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_83),
.A2(n_35),
.B1(n_0),
.B2(n_6),
.Y(n_226)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_142),
.B(n_110),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_232),
.B(n_233),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_110),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_153),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_236),
.B(n_268),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_129),
.B1(n_102),
.B2(n_118),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_238),
.A2(n_242),
.B1(n_288),
.B2(n_225),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_140),
.B(n_77),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_240),
.B(n_253),
.Y(n_340)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_241),
.Y(n_330)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_147),
.B(n_77),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_249),
.B(n_254),
.Y(n_347)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_250),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_0),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_177),
.B(n_93),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_255),
.B(n_256),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_137),
.A2(n_65),
.B(n_59),
.C(n_103),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_0),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_258),
.B(n_271),
.Y(n_358)
);

BUFx12_ASAP7_75t_L g259 ( 
.A(n_163),
.Y(n_259)
);

INVx13_ASAP7_75t_L g343 ( 
.A(n_259),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_106),
.C(n_99),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_261),
.B(n_293),
.C(n_295),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_141),
.B(n_70),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_263),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_171),
.B(n_69),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_168),
.Y(n_264)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_264),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_97),
.B1(n_92),
.B2(n_127),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_265),
.A2(n_314),
.B1(n_155),
.B2(n_247),
.Y(n_322)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_156),
.Y(n_267)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_269),
.A2(n_300),
.B1(n_309),
.B2(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_181),
.B(n_5),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_153),
.B(n_95),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_272),
.B(n_275),
.Y(n_329)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_138),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_273),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_153),
.B(n_90),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_167),
.A2(n_124),
.B1(n_7),
.B2(n_9),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_277),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_167),
.A2(n_6),
.B1(n_9),
.B2(n_14),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_136),
.B(n_15),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_282),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_15),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_143),
.Y(n_284)
);

INVx4_ASAP7_75t_SL g351 ( 
.A(n_284),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_218),
.A2(n_139),
.B1(n_192),
.B2(n_166),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

BUFx12_ASAP7_75t_L g287 ( 
.A(n_163),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_152),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_133),
.B(n_184),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_151),
.B(n_18),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_296),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_202),
.B(n_19),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_189),
.B(n_19),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_209),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_185),
.B(n_19),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_298),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_185),
.B(n_202),
.Y(n_298)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_144),
.Y(n_299)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_187),
.A2(n_170),
.B1(n_190),
.B2(n_145),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_143),
.B(n_135),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_306),
.Y(n_360)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_138),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_135),
.Y(n_303)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_144),
.Y(n_304)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

BUFx12_ASAP7_75t_L g305 ( 
.A(n_145),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_157),
.B(n_165),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_170),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_308),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_190),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_134),
.A2(n_149),
.B1(n_182),
.B2(n_188),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_157),
.B(n_165),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_149),
.A2(n_182),
.B1(n_180),
.B2(n_162),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_172),
.B(n_191),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_172),
.Y(n_316)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_318),
.B(n_288),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_322),
.A2(n_332),
.B1(n_348),
.B2(n_374),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_164),
.B1(n_224),
.B2(n_146),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_324),
.A2(n_331),
.B1(n_344),
.B2(n_304),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_266),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_339),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_164),
.B1(n_224),
.B2(n_207),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_314),
.A2(n_159),
.B1(n_160),
.B2(n_197),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g338 ( 
.A(n_268),
.B(n_180),
.C(n_191),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_268),
.C(n_256),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_266),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_242),
.A2(n_207),
.B1(n_205),
.B2(n_169),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_244),
.A2(n_159),
.B1(n_160),
.B2(n_212),
.Y(n_348)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_248),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_359),
.Y(n_404)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_243),
.Y(n_370)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_245),
.Y(n_372)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_233),
.A2(n_308),
.B1(n_307),
.B2(n_290),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_373),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_251),
.A2(n_197),
.B1(n_212),
.B2(n_169),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_250),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_251),
.A2(n_232),
.B(n_240),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_376),
.A2(n_236),
.B(n_280),
.Y(n_428)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_264),
.Y(n_377)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_270),
.Y(n_378)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_252),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_258),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_386),
.B(n_363),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_345),
.B(n_252),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_387),
.B(n_389),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_388),
.A2(n_413),
.B1(n_414),
.B2(n_422),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_254),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_291),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_393),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_325),
.B(n_246),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_392),
.B(n_409),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_253),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_291),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_394),
.B(n_396),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_325),
.B(n_257),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_355),
.A2(n_366),
.B(n_363),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_398),
.A2(n_356),
.B(n_353),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_400),
.A2(n_411),
.B1(n_416),
.B2(n_417),
.Y(n_436)
);

A2O1A1O1Ixp25_ASAP7_75t_L g401 ( 
.A1(n_355),
.A2(n_251),
.B(n_234),
.C(n_255),
.D(n_249),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_401),
.A2(n_428),
.B(n_368),
.Y(n_449)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_364),
.B(n_271),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_405),
.B(n_418),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_323),
.A2(n_284),
.B1(n_277),
.B2(n_316),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_234),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_420),
.C(n_369),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_324),
.A2(n_331),
.B1(n_318),
.B2(n_334),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_340),
.B(n_282),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_412),
.B(n_415),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_322),
.A2(n_261),
.B1(n_295),
.B2(n_281),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_344),
.A2(n_293),
.B1(n_298),
.B2(n_294),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_340),
.B(n_293),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_334),
.A2(n_175),
.B1(n_205),
.B2(n_204),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_326),
.A2(n_204),
.B1(n_304),
.B2(n_237),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_278),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_349),
.B(n_278),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_419),
.B(n_423),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_365),
.B(n_237),
.C(n_239),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_365),
.A2(n_299),
.B1(n_239),
.B2(n_313),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_350),
.B(n_319),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_321),
.A2(n_299),
.B1(n_313),
.B2(n_260),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_424),
.A2(n_425),
.B1(n_351),
.B2(n_362),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_332),
.A2(n_280),
.B1(n_260),
.B2(n_286),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_347),
.B(n_337),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_427),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_329),
.B(n_235),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_347),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_429),
.B(n_433),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_418),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_447),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_432),
.B(n_448),
.C(n_455),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_360),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_411),
.A2(n_348),
.B1(n_374),
.B2(n_346),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_437),
.A2(n_451),
.B1(n_464),
.B2(n_425),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_380),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_444),
.B(n_450),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_399),
.A2(n_338),
.B1(n_323),
.B2(n_346),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_446),
.A2(n_453),
.B1(n_470),
.B2(n_398),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_380),
.Y(n_447)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_387),
.C(n_384),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_449),
.A2(n_467),
.B(n_468),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_396),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_357),
.B1(n_366),
.B2(n_372),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_399),
.A2(n_357),
.B1(n_328),
.B2(n_370),
.Y(n_453)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_328),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_381),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_466),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_459),
.A2(n_383),
.B1(n_390),
.B2(n_395),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_463),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_394),
.B(n_320),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_400),
.A2(n_320),
.B1(n_369),
.B2(n_362),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_378),
.C(n_377),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_382),
.A2(n_351),
.B1(n_354),
.B2(n_330),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_413),
.A2(n_367),
.B1(n_356),
.B2(n_353),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_472),
.A2(n_476),
.B1(n_485),
.B2(n_491),
.Y(n_513)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_439),
.Y(n_473)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_473),
.Y(n_514)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_439),
.Y(n_474)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_474),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_405),
.Y(n_477)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_460),
.A2(n_386),
.B(n_424),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_479),
.A2(n_478),
.B(n_476),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_436),
.A2(n_423),
.B1(n_391),
.B2(n_388),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_481),
.A2(n_508),
.B1(n_466),
.B2(n_437),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_458),
.Y(n_482)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_482),
.Y(n_530)
);

XOR2x1_ASAP7_75t_SL g483 ( 
.A(n_448),
.B(n_401),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_483),
.B(n_463),
.Y(n_527)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_484),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_414),
.B1(n_419),
.B2(n_389),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_390),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_496),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

INVx13_ASAP7_75t_L g542 ( 
.A(n_489),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_453),
.A2(n_393),
.B1(n_395),
.B2(n_407),
.Y(n_491)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_493),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_494),
.A2(n_498),
.B1(n_461),
.B2(n_438),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_431),
.A2(n_410),
.B1(n_403),
.B2(n_383),
.Y(n_495)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_495),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_430),
.B(n_402),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_454),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_497),
.B(n_501),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_470),
.A2(n_412),
.B1(n_417),
.B2(n_415),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_503),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_441),
.B(n_336),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_469),
.A2(n_397),
.B(n_402),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_502),
.A2(n_404),
.B(n_379),
.Y(n_541)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_468),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_504),
.Y(n_537)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_506),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_457),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_464),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_507),
.B(n_509),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_436),
.A2(n_397),
.B1(n_421),
.B2(n_342),
.Y(n_508)
);

AO22x1_ASAP7_75t_L g509 ( 
.A1(n_446),
.A2(n_416),
.B1(n_379),
.B2(n_367),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_492),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_510),
.B(n_531),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_478),
.A2(n_449),
.B(n_460),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_511),
.A2(n_524),
.B(n_479),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_512),
.A2(n_516),
.B1(n_521),
.B2(n_522),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_481),
.A2(n_434),
.B1(n_440),
.B2(n_442),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_462),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_519),
.B(n_528),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_432),
.C(n_429),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_520),
.B(n_534),
.C(n_535),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_485),
.A2(n_434),
.B1(n_442),
.B2(n_440),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_507),
.A2(n_461),
.B1(n_455),
.B2(n_451),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_523),
.A2(n_540),
.B1(n_544),
.B2(n_509),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_527),
.B(n_529),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_490),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_490),
.B(n_433),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g531 ( 
.A(n_471),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_487),
.B(n_443),
.C(n_317),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_480),
.B(n_317),
.C(n_354),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_483),
.B(n_471),
.C(n_477),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_539),
.B(n_545),
.C(n_546),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_508),
.A2(n_457),
.B1(n_467),
.B2(n_404),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_491),
.A2(n_342),
.B1(n_341),
.B2(n_351),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_486),
.B(n_333),
.C(n_302),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_333),
.C(n_286),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_493),
.Y(n_548)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_548),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_502),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_560),
.Y(n_579)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_551),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_552),
.A2(n_577),
.B1(n_512),
.B2(n_538),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_525),
.B(n_498),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_553),
.B(n_557),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_515),
.B(n_473),
.Y(n_554)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_554),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_518),
.Y(n_555)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_555),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_530),
.B(n_488),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_539),
.B(n_488),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_558),
.B(n_561),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_475),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_517),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_518),
.B(n_499),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_563),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_532),
.B(n_505),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_520),
.B(n_475),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g591 ( 
.A(n_565),
.B(n_533),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_566),
.A2(n_511),
.B(n_524),
.Y(n_578)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_514),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_568),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_522),
.B(n_503),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_569),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_528),
.B(n_474),
.C(n_335),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_572),
.C(n_575),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_529),
.B(n_509),
.Y(n_572)
);

INVxp33_ASAP7_75t_L g573 ( 
.A(n_540),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_573),
.B(n_541),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_521),
.B(n_516),
.Y(n_574)
);

AOI221xp5_ASAP7_75t_L g589 ( 
.A1(n_574),
.A2(n_543),
.B1(n_544),
.B2(n_532),
.C(n_533),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_523),
.B(n_371),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_526),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_576),
.Y(n_590)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_536),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_578),
.A2(n_585),
.B(n_559),
.Y(n_617)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_582),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_564),
.B(n_535),
.C(n_513),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_586),
.B(n_591),
.Y(n_622)
);

A2O1A1O1Ixp25_ASAP7_75t_L g588 ( 
.A1(n_549),
.A2(n_527),
.B(n_543),
.C(n_546),
.D(n_545),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_600),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_589),
.Y(n_611)
);

INVx13_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_592),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_573),
.A2(n_506),
.B1(n_484),
.B2(n_489),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_595),
.A2(n_552),
.B1(n_571),
.B2(n_563),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_564),
.B(n_506),
.C(n_371),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_596),
.B(n_547),
.C(n_550),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_549),
.A2(n_542),
.B1(n_341),
.B2(n_359),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_597),
.A2(n_580),
.B1(n_590),
.B2(n_585),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_556),
.A2(n_542),
.B1(n_361),
.B2(n_303),
.Y(n_600)
);

XOR2x2_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_343),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_602),
.B(n_560),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_603),
.A2(n_583),
.B1(n_598),
.B2(n_594),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_604),
.B(n_617),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_565),
.C(n_570),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_605),
.B(n_609),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_581),
.A2(n_599),
.B(n_601),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_608),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_596),
.B(n_547),
.C(n_567),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_579),
.B(n_567),
.C(n_571),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_610),
.B(n_613),
.C(n_616),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_579),
.B(n_566),
.C(n_575),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_593),
.A2(n_554),
.B1(n_562),
.B2(n_548),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_598),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_591),
.B(n_274),
.Y(n_615)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_615),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_584),
.B(n_559),
.C(n_274),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_580),
.B(n_274),
.Y(n_618)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_618),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_273),
.C(n_296),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_619),
.B(n_604),
.C(n_616),
.Y(n_631)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_620),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_601),
.A2(n_241),
.B1(n_267),
.B2(n_343),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_623),
.A2(n_595),
.B1(n_583),
.B2(n_587),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_611),
.A2(n_612),
.B(n_585),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g641 ( 
.A1(n_624),
.A2(n_607),
.B(n_617),
.Y(n_641)
);

INVxp33_ASAP7_75t_L g642 ( 
.A(n_626),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_611),
.B(n_590),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_639),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_629),
.A2(n_636),
.B1(n_638),
.B2(n_305),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_631),
.B(n_619),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_607),
.A2(n_621),
.B1(n_612),
.B2(n_578),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_632),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_620),
.B(n_587),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_605),
.B(n_602),
.C(n_597),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_623),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_640),
.B(n_588),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_646),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_643),
.B(n_647),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_610),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_627),
.B(n_609),
.C(n_622),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_630),
.B(n_613),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_648),
.B(n_651),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_649),
.A2(n_650),
.B(n_625),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_630),
.B(n_592),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_627),
.B(n_343),
.C(n_305),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_305),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_652),
.B(n_653),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_645),
.A2(n_632),
.B1(n_637),
.B2(n_629),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_654),
.A2(n_660),
.B1(n_641),
.B2(n_259),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_648),
.B(n_624),
.Y(n_657)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_657),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g664 ( 
.A(n_659),
.B(n_642),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_642),
.A2(n_625),
.B1(n_636),
.B2(n_633),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_644),
.A2(n_634),
.B(n_639),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_662),
.A2(n_647),
.B(n_645),
.Y(n_663)
);

OAI31xp33_ASAP7_75t_SL g670 ( 
.A1(n_663),
.A2(n_668),
.A3(n_259),
.B(n_287),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_664),
.A2(n_657),
.B(n_654),
.Y(n_669)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_661),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_L g671 ( 
.A(n_666),
.B(n_667),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_655),
.A2(n_259),
.B(n_287),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_669),
.A2(n_670),
.B(n_665),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_672),
.B(n_673),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_671),
.B(n_658),
.C(n_656),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_674),
.A2(n_656),
.B(n_658),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_675),
.B(n_287),
.Y(n_676)
);


endmodule