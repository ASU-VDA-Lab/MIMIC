module fake_netlist_6_2461_n_1728 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1728);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1728;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_62),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_18),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_17),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_65),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_61),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_64),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_19),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_38),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_95),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_1),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_142),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_78),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_87),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_59),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_77),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_118),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_35),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_101),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_26),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_33),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_153),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_27),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_86),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_99),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_102),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_72),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_10),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_116),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_42),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_113),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_93),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_89),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_70),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_158),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_22),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_17),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_6),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_14),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_107),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_32),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_129),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_31),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_10),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_34),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_55),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_2),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_83),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_98),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_122),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_151),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_157),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_23),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_140),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_136),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_23),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_159),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_126),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_143),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_167),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_55),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_161),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_71),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_41),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_54),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_51),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_108),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_160),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_20),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_47),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_19),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_128),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_52),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_26),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_13),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_35),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_8),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_12),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_60),
.Y(n_310)
);

BUFx8_ASAP7_75t_SL g311 ( 
.A(n_14),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_7),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_47),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_73),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_88),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_155),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_31),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_51),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_85),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_124),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_37),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_131),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_48),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_149),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_46),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_21),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_16),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_119),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_94),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_5),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_92),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_68),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_21),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_52),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_30),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_154),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_8),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_114),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_24),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_82),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_33),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_3),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_30),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_74),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_112),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_197),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_311),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_178),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_181),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_174),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_294),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_281),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_242),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_219),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_207),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_334),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_210),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_180),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_213),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_244),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_241),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_222),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_181),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_217),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_205),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_209),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_178),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_228),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_184),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_237),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_240),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_230),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_250),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_254),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_278),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_232),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_280),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_284),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_221),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_290),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_319),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_184),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_295),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_296),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_257),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_299),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_308),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_330),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_223),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_196),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_188),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_292),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_225),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_182),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_178),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_188),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_235),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_178),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_175),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_236),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_175),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_186),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_182),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_178),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_211),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_211),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_257),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_316),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_422),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_422),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_316),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_364),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_348),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_186),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_387),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_373),
.B(n_234),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_234),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_349),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_400),
.B(n_268),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_355),
.A2(n_335),
.B1(n_344),
.B2(n_343),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_268),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_384),
.A2(n_190),
.B1(n_344),
.B2(n_343),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_352),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_176),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_352),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_356),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_191),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_356),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_359),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_351),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_359),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_357),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_357),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

AND3x2_ASAP7_75t_L g474 ( 
.A(n_406),
.B(n_302),
.C(n_204),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_358),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_377),
.A2(n_265),
.B1(n_342),
.B2(n_203),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_362),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_363),
.A2(n_195),
.B1(n_342),
.B2(n_190),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_358),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_420),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_432),
.B(n_196),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_351),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_351),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_360),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_433),
.B(n_201),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_362),
.B(n_206),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_351),
.B(n_187),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_360),
.Y(n_488)
);

BUFx8_ASAP7_75t_L g489 ( 
.A(n_417),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_366),
.B(n_208),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_351),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_366),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_367),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_424),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_385),
.B(n_196),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_434),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_431),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_431),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_367),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_379),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_371),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_361),
.B(n_215),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_427),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_350),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_385),
.B(n_315),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_393),
.B(n_315),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_371),
.B(n_226),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_393),
.B(n_229),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_372),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_468),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_444),
.B(n_415),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_441),
.B(n_415),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_451),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_418),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_454),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_468),
.Y(n_523)
);

INVx8_ASAP7_75t_L g524 ( 
.A(n_490),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_187),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_470),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_470),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_481),
.B(n_368),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_469),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_481),
.B(n_368),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_374),
.C(n_372),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_490),
.A2(n_417),
.B1(n_353),
.B2(n_374),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_SL g538 ( 
.A(n_499),
.B(n_509),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_469),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_456),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_476),
.A2(n_305),
.B1(n_258),
.B2(n_252),
.Y(n_545)
);

AOI21x1_ASAP7_75t_L g546 ( 
.A1(n_461),
.A2(n_428),
.B(n_426),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_452),
.A2(n_233),
.B(n_231),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_476),
.A2(n_478),
.B1(n_489),
.B2(n_398),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_477),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_490),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_469),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_464),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_510),
.Y(n_557)
);

AND3x2_ASAP7_75t_L g558 ( 
.A(n_499),
.B(n_423),
.C(n_403),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_453),
.B(n_243),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_510),
.A2(n_429),
.B1(n_428),
.B2(n_426),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_440),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_460),
.A2(n_247),
.B1(n_337),
.B2(n_333),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_443),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_457),
.B(n_315),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_446),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_459),
.B(n_429),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_482),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_447),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_482),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_478),
.B(n_193),
.Y(n_573)
);

NOR2x1p5_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_193),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_480),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_445),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_510),
.A2(n_370),
.B1(n_187),
.B2(n_288),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_466),
.A2(n_275),
.B(n_255),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_482),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_482),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_437),
.B(n_404),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_498),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_449),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_438),
.Y(n_588)
);

NOR2x1p5_ASAP7_75t_L g589 ( 
.A(n_437),
.B(n_195),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_510),
.A2(n_187),
.B1(n_212),
.B2(n_288),
.Y(n_591)
);

BUFx10_ASAP7_75t_L g592 ( 
.A(n_496),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_498),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_439),
.B(n_345),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_R g595 ( 
.A(n_506),
.B(n_177),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_467),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_455),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_503),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_SL g600 ( 
.A(n_508),
.B(n_203),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_485),
.B(n_437),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_504),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_467),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_473),
.B(n_397),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_471),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_463),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_508),
.B(n_345),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_471),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_458),
.B(n_416),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_489),
.B(n_345),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_489),
.B(n_177),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_473),
.B(n_279),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_489),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_473),
.B(n_179),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_486),
.A2(n_324),
.B1(n_331),
.B2(n_338),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_463),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_472),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_L g619 ( 
.A(n_487),
.B(n_187),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_475),
.A2(n_261),
.B1(n_259),
.B2(n_256),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_475),
.B(n_325),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_479),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_486),
.B(n_179),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_479),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_435),
.B(n_285),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_435),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_435),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_435),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_484),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_504),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_484),
.B(n_402),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_488),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_486),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_488),
.B(n_494),
.C(n_492),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_492),
.B(n_411),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_486),
.B(n_183),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_483),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_R g639 ( 
.A(n_494),
.B(n_238),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_502),
.B(n_183),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_512),
.B(n_185),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_474),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_512),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_487),
.B(n_212),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_504),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_493),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_504),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_504),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_504),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_483),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_483),
.B(n_185),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_493),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_487),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_483),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_497),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_501),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_483),
.B(n_189),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_500),
.B(n_329),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_487),
.A2(n_324),
.B1(n_331),
.B2(n_338),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_491),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_483),
.B(n_189),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_633),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_585),
.B(n_593),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_515),
.B(n_491),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_515),
.B(n_491),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_513),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_583),
.B(n_404),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_614),
.B(n_416),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_521),
.B(n_339),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_529),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g676 ( 
.A(n_588),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_585),
.B(n_239),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_621),
.A2(n_410),
.B(n_413),
.C(n_405),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_627),
.B(n_192),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_559),
.A2(n_298),
.B1(n_310),
.B2(n_314),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_529),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_552),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_518),
.B(n_491),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_627),
.B(n_192),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_601),
.B(n_500),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_517),
.B(n_194),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_589),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_631),
.B(n_194),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_537),
.B(n_198),
.Y(n_689)
);

AND2x6_ASAP7_75t_SL g690 ( 
.A(n_604),
.B(n_386),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_552),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_513),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_626),
.B(n_500),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_524),
.B(n_245),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_595),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_626),
.B(n_500),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_639),
.B(n_198),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_628),
.B(n_557),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_628),
.A2(n_495),
.B(n_321),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_635),
.B(n_419),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_514),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_557),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_542),
.B(n_199),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_565),
.B(n_199),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_589),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_518),
.B(n_287),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_557),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_528),
.B(n_532),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_600),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_607),
.B(n_200),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_574),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_524),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_614),
.B(n_419),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_576),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_524),
.B(n_246),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_574),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_654),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_579),
.A2(n_288),
.B1(n_212),
.B2(n_487),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_654),
.B(n_212),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_519),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_648),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_662),
.B(n_200),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_566),
.B(n_569),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_519),
.B(n_495),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_533),
.B(n_248),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_520),
.B(n_495),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_594),
.B(n_202),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_616),
.B(n_262),
.C(n_269),
.Y(n_728)
);

INVxp33_ASAP7_75t_L g729 ( 
.A(n_609),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_662),
.B(n_202),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_522),
.B(n_495),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_522),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_538),
.B(n_386),
.C(n_388),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_615),
.B(n_332),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_535),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_559),
.B(n_332),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_540),
.B(n_544),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_578),
.B(n_616),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_559),
.A2(n_303),
.B1(n_263),
.B2(n_260),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_559),
.B(n_341),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_514),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_524),
.B(n_249),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_559),
.B(n_341),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_625),
.B(n_346),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_625),
.B(n_410),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_625),
.A2(n_251),
.B1(n_291),
.B2(n_289),
.Y(n_746)
);

INVx8_ASAP7_75t_L g747 ( 
.A(n_613),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_640),
.B(n_346),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_544),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_524),
.A2(n_495),
.B(n_212),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_625),
.B(n_270),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_579),
.A2(n_288),
.B1(n_487),
.B2(n_257),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_661),
.B(n_271),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_549),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_549),
.B(n_495),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_533),
.B(n_272),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_523),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_L g758 ( 
.A(n_591),
.B(n_273),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_526),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_620),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_609),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_623),
.A2(n_323),
.B1(n_297),
.B2(n_286),
.Y(n_762)
);

INVx8_ASAP7_75t_L g763 ( 
.A(n_613),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_556),
.A2(n_276),
.B1(n_283),
.B2(n_320),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_556),
.B(n_216),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_637),
.A2(n_547),
.B1(n_525),
.B2(n_613),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_646),
.A2(n_413),
.B(n_396),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_649),
.B(n_388),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_568),
.B(n_487),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_527),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_568),
.B(n_389),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_516),
.B(n_389),
.Y(n_772)
);

AND2x2_ASAP7_75t_SL g773 ( 
.A(n_545),
.B(n_643),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_577),
.B(n_391),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_596),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_653),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_596),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_597),
.B(n_391),
.Y(n_778)
);

CKINVDCx16_ASAP7_75t_R g779 ( 
.A(n_592),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_531),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_547),
.A2(n_412),
.B1(n_409),
.B2(n_408),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_579),
.A2(n_322),
.B1(n_218),
.B2(n_313),
.Y(n_782)
);

AOI221xp5_ASAP7_75t_L g783 ( 
.A1(n_573),
.A2(n_545),
.B1(n_564),
.B2(n_550),
.C(n_266),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_597),
.B(n_392),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_592),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_547),
.A2(n_322),
.B1(n_220),
.B2(n_317),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_536),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_599),
.B(n_392),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_603),
.B(n_394),
.Y(n_789)
);

CKINVDCx11_ASAP7_75t_R g790 ( 
.A(n_592),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_642),
.B(n_224),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_605),
.B(n_394),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_605),
.B(n_395),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_608),
.B(n_395),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_558),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_610),
.B(n_412),
.C(n_409),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_643),
.B(n_396),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_608),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_613),
.A2(n_408),
.B1(n_407),
.B2(n_405),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_611),
.B(n_253),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_536),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_612),
.B(n_399),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_612),
.A2(n_322),
.B1(n_264),
.B2(n_301),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_618),
.B(n_267),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_618),
.B(n_399),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_622),
.B(n_307),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_622),
.B(n_306),
.Y(n_807)
);

AND2x2_ASAP7_75t_SL g808 ( 
.A(n_619),
.B(n_407),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_629),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_629),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_641),
.B(n_300),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_SL g812 ( 
.A(n_575),
.B(n_318),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_641),
.A2(n_293),
.B1(n_274),
.B2(n_277),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_576),
.B(n_401),
.C(n_282),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_624),
.B(n_401),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_380),
.C(n_378),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_575),
.B(n_654),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_632),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_575),
.B(n_380),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_632),
.B(n_378),
.Y(n_820)
);

AND2x6_ASAP7_75t_SL g821 ( 
.A(n_613),
.B(n_376),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_564),
.A2(n_376),
.B1(n_375),
.B2(n_146),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_564),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_644),
.B(n_375),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_717),
.B(n_654),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_673),
.B(n_644),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_818),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_738),
.A2(n_564),
.B1(n_634),
.B2(n_562),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_737),
.B(n_647),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_783),
.A2(n_571),
.B1(n_561),
.B2(n_562),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_776),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_720),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_722),
.A2(n_567),
.B1(n_571),
.B2(n_563),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_717),
.A2(n_698),
.B(n_696),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_737),
.B(n_647),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_717),
.B(n_575),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_774),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_698),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_700),
.B(n_592),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_732),
.B(n_646),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_776),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_788),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_703),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_735),
.B(n_650),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_717),
.B(n_649),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_760),
.A2(n_560),
.B1(n_663),
.B2(n_650),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_729),
.A2(n_567),
.B1(n_563),
.B2(n_554),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_712),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_749),
.B(n_663),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_712),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_SL g851 ( 
.A(n_728),
.B(n_664),
.C(n_659),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_675),
.B(n_602),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_675),
.B(n_602),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_761),
.B(n_652),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_712),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_754),
.B(n_541),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_775),
.B(n_548),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_777),
.B(n_548),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_797),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_730),
.A2(n_561),
.B1(n_580),
.B2(n_555),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_675),
.B(n_602),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_688),
.A2(n_555),
.B(n_580),
.C(n_554),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_798),
.B(n_551),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_702),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_702),
.B(n_602),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_809),
.B(n_551),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_810),
.B(n_539),
.Y(n_867)
);

INVx5_ASAP7_75t_L g868 ( 
.A(n_780),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_723),
.A2(n_630),
.B1(n_658),
.B2(n_660),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_790),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_667),
.B(n_539),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_671),
.B(n_539),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_708),
.A2(n_630),
.B1(n_658),
.B2(n_660),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_823),
.A2(n_586),
.B1(n_587),
.B2(n_590),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_668),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_714),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_721),
.B(n_586),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_676),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_804),
.B(n_584),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_665),
.B(n_587),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_797),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_702),
.B(n_630),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_745),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_674),
.B(n_584),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_681),
.B(n_584),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_693),
.A2(n_630),
.B(n_531),
.Y(n_886)
);

BUFx12f_ASAP7_75t_SL g887 ( 
.A(n_672),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_711),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_745),
.B(n_590),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_682),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_670),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_687),
.B(n_598),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_668),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_766),
.B(n_531),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_691),
.B(n_584),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_707),
.B(n_638),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_822),
.B(n_695),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_734),
.B(n_771),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_692),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_812),
.B(n_531),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_669),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_771),
.B(n_638),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_669),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_683),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_701),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_683),
.Y(n_906)
);

O2A1O1Ixp5_ASAP7_75t_L g907 ( 
.A1(n_753),
.A2(n_657),
.B(n_656),
.C(n_546),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_779),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_704),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_716),
.B(n_666),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_778),
.B(n_638),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_820),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_709),
.B(n_780),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_780),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_778),
.B(n_638),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_736),
.A2(n_656),
.B1(n_598),
.B2(n_606),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_718),
.A2(n_606),
.B1(n_617),
.B2(n_657),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_765),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_820),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_705),
.B(n_617),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_SL g921 ( 
.A(n_786),
.B(n_655),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_784),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_747),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_824),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_824),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_685),
.A2(n_655),
.B(n_651),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_726),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_784),
.B(n_570),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_719),
.A2(n_715),
.B(n_694),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_789),
.B(n_570),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_789),
.B(n_570),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_773),
.B(n_572),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_672),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_726),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_785),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_740),
.A2(n_572),
.B1(n_534),
.B2(n_543),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_741),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_769),
.B(n_655),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_731),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_686),
.B(n_546),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_792),
.B(n_572),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_817),
.B(n_553),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_731),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_792),
.B(n_581),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_755),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_793),
.B(n_581),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_806),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_769),
.B(n_655),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_755),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_793),
.B(n_581),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_815),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_747),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_757),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_724),
.Y(n_954)
);

BUFx2_ASAP7_75t_SL g955 ( 
.A(n_772),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_679),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_794),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_794),
.B(n_553),
.Y(n_958)
);

AND2x6_ASAP7_75t_SL g959 ( 
.A(n_800),
.B(n_0),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_802),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_807),
.Y(n_961)
);

INVxp67_ASAP7_75t_SL g962 ( 
.A(n_802),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_725),
.B(n_655),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_689),
.B(n_543),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_743),
.A2(n_553),
.B1(n_534),
.B2(n_636),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_805),
.B(n_543),
.Y(n_966)
);

NOR2x1p5_ASAP7_75t_L g967 ( 
.A(n_805),
.B(n_636),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_690),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_759),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_756),
.B(n_651),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_796),
.B(n_636),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_770),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_787),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_672),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_801),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_795),
.B(n_651),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_811),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_819),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_733),
.B(n_582),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_713),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_719),
.Y(n_981)
);

AO22x1_ASAP7_75t_L g982 ( 
.A1(n_727),
.A2(n_582),
.B1(n_534),
.B2(n_530),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_706),
.B(n_582),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_748),
.B(n_791),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_747),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_710),
.B(n_530),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_781),
.B(n_530),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_684),
.B(n_651),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_SL g989 ( 
.A(n_814),
.B(n_2),
.C(n_3),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_697),
.B(n_645),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_SL g991 ( 
.A(n_763),
.B(n_651),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_782),
.B(n_531),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_744),
.B(n_4),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_677),
.B(n_6),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_768),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_803),
.B(n_11),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_768),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_808),
.B(n_12),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_984),
.B(n_746),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_825),
.A2(n_742),
.B(n_763),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_922),
.B(n_799),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_897),
.A2(n_993),
.B(n_898),
.C(n_998),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_993),
.A2(n_957),
.B(n_960),
.C(n_897),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_839),
.B(n_813),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_832),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_825),
.A2(n_763),
.B(n_750),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_843),
.A2(n_909),
.B1(n_932),
.B2(n_956),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_842),
.B(n_764),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_989),
.A2(n_680),
.B(n_678),
.C(n_751),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_929),
.A2(n_758),
.B(n_699),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_899),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_883),
.B(n_739),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_878),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_837),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_962),
.B(n_762),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_883),
.B(n_752),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_962),
.A2(n_816),
.B1(n_767),
.B2(n_821),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_951),
.B(n_15),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_981),
.A2(n_145),
.B(n_144),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_935),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_900),
.A2(n_141),
.B(n_139),
.C(n_135),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_994),
.A2(n_15),
.B(n_20),
.C(n_22),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_912),
.B(n_24),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_952),
.B(n_132),
.Y(n_1024)
);

BUFx4_ASAP7_75t_SL g1025 ( 
.A(n_876),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_923),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_838),
.B(n_120),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_SL g1028 ( 
.A(n_848),
.B(n_850),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_952),
.B(n_117),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_877),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_932),
.A2(n_111),
.B1(n_105),
.B2(n_104),
.Y(n_1031)
);

NOR2xp67_ASAP7_75t_L g1032 ( 
.A(n_888),
.B(n_100),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_996),
.A2(n_25),
.B(n_28),
.C(n_29),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_919),
.B(n_25),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_910),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_905),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_908),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_924),
.B(n_36),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_828),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_828),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_838),
.B(n_91),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_968),
.B(n_43),
.C(n_44),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_981),
.A2(n_894),
.B(n_834),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_925),
.B(n_43),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_848),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_910),
.B(n_920),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_848),
.Y(n_1047)
);

AOI21x1_ASAP7_75t_L g1048 ( 
.A1(n_982),
.A2(n_970),
.B(n_963),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_854),
.B(n_45),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_894),
.A2(n_914),
.B(n_868),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_978),
.B(n_45),
.Y(n_1051)
);

BUFx4f_ASAP7_75t_SL g1052 ( 
.A(n_870),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_826),
.B(n_875),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_848),
.B(n_57),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_905),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_893),
.B(n_46),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_923),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_859),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_901),
.B(n_50),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_918),
.B(n_63),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_947),
.B(n_58),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_920),
.B(n_76),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_937),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_903),
.B(n_79),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_856),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_889),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_868),
.A2(n_914),
.B(n_835),
.Y(n_1067)
);

AO22x1_ASAP7_75t_L g1068 ( 
.A1(n_974),
.A2(n_53),
.B1(n_81),
.B2(n_881),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_887),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_880),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_847),
.A2(n_913),
.B(n_900),
.C(n_992),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_868),
.A2(n_914),
.B(n_829),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_868),
.A2(n_914),
.B(n_861),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_830),
.A2(n_906),
.B1(n_904),
.B2(n_874),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_923),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_850),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_850),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_852),
.A2(n_853),
.B(n_861),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_961),
.B(n_977),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_864),
.B(n_933),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_980),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_830),
.A2(n_874),
.B1(n_927),
.B2(n_949),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_964),
.A2(n_889),
.B1(n_979),
.B2(n_967),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_934),
.B(n_939),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_985),
.B(n_892),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_964),
.A2(n_851),
.B(n_988),
.C(n_921),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_943),
.A2(n_945),
.B1(n_860),
.B2(n_833),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_852),
.A2(n_865),
.B(n_853),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_954),
.B(n_827),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_865),
.A2(n_882),
.B(n_845),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_963),
.A2(n_970),
.B(n_862),
.C(n_913),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_938),
.A2(n_948),
.B(n_862),
.C(n_995),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_882),
.A2(n_845),
.B(n_879),
.Y(n_1093)
);

AND2x4_ASAP7_75t_SL g1094 ( 
.A(n_985),
.B(n_850),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_955),
.B(n_933),
.Y(n_1095)
);

OR2x6_ASAP7_75t_SL g1096 ( 
.A(n_846),
.B(n_872),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_847),
.A2(n_940),
.B(n_987),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_890),
.B(n_902),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_851),
.A2(n_979),
.B(n_986),
.C(n_907),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_985),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_864),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_926),
.A2(n_886),
.B(n_915),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_840),
.A2(n_844),
.B(n_849),
.C(n_871),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_911),
.A2(n_866),
.B(n_863),
.C(n_858),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_928),
.A2(n_941),
.B(n_946),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_855),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_855),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_973),
.B(n_836),
.Y(n_1108)
);

BUFx2_ASAP7_75t_R g1109 ( 
.A(n_836),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_857),
.A2(n_931),
.B(n_944),
.C(n_950),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_971),
.B(n_953),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_855),
.B(n_971),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_930),
.B(n_966),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_831),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_959),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_991),
.B(n_841),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_990),
.B(n_976),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_891),
.B(n_975),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_997),
.A2(n_958),
.B(n_916),
.C(n_983),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_867),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_969),
.B(n_972),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_997),
.A2(n_833),
.B(n_860),
.C(n_972),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_942),
.B(n_895),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_942),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_884),
.A2(n_885),
.B(n_896),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_936),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_873),
.A2(n_869),
.B(n_917),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_917),
.A2(n_984),
.B1(n_962),
.B2(n_957),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_L g1129 ( 
.A1(n_984),
.A2(n_900),
.B(n_688),
.C(n_898),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_922),
.B(n_984),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_922),
.B(n_984),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_984),
.A2(n_993),
.B(n_898),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_984),
.A2(n_962),
.B1(n_957),
.B2(n_960),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_832),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_899),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1053),
.B(n_1084),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1020),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1132),
.B(n_1130),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_1062),
.B(n_1024),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1005),
.Y(n_1140)
);

AOI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1048),
.A2(n_1093),
.B(n_1043),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1010),
.A2(n_1105),
.B(n_1102),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1078),
.A2(n_1088),
.B(n_1090),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1025),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1099),
.A2(n_1129),
.B(n_1002),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1113),
.A2(n_1110),
.B(n_1103),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_1037),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1013),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_1133),
.A2(n_1003),
.A3(n_1128),
.B(n_1087),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1050),
.A2(n_1006),
.B(n_1125),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1013),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1104),
.A2(n_1000),
.B(n_1015),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1131),
.B(n_1065),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1030),
.A2(n_1074),
.B1(n_1082),
.B2(n_1040),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1074),
.B(n_1082),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1091),
.A2(n_1071),
.B(n_1119),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1127),
.A2(n_1117),
.B(n_999),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1033),
.B(n_1008),
.C(n_1066),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1016),
.A2(n_1098),
.B(n_1120),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_SL g1160 ( 
.A1(n_1039),
.A2(n_1097),
.B(n_1116),
.C(n_1012),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1030),
.B(n_1004),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_1035),
.B(n_1007),
.Y(n_1162)
);

AOI211x1_ASAP7_75t_L g1163 ( 
.A1(n_1018),
.A2(n_1038),
.B(n_1044),
.C(n_1034),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1097),
.A2(n_1087),
.B(n_1092),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_R g1165 ( 
.A(n_1069),
.B(n_1046),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1026),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1122),
.A2(n_1108),
.A3(n_1017),
.B(n_1064),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1009),
.B(n_1022),
.C(n_1083),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1126),
.A2(n_1064),
.B(n_1017),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1073),
.A2(n_1072),
.B(n_1067),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1026),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1134),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1089),
.B(n_1070),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1096),
.A2(n_1001),
.B1(n_1023),
.B2(n_1056),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1070),
.B(n_1111),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1026),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1036),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_1014),
.B(n_1095),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1135),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1057),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1123),
.A2(n_1124),
.B(n_1121),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1114),
.B(n_1085),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1114),
.B(n_1085),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1062),
.A2(n_1079),
.B1(n_1112),
.B2(n_1061),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_1028),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1057),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1021),
.A2(n_1059),
.B(n_1019),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1112),
.B(n_1063),
.Y(n_1188)
);

AOI31xp67_ASAP7_75t_L g1189 ( 
.A1(n_1027),
.A2(n_1041),
.A3(n_1060),
.B(n_1055),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1042),
.A2(n_1051),
.B(n_1080),
.C(n_1049),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1054),
.A2(n_1076),
.B(n_1077),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1024),
.B(n_1029),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1029),
.A2(n_1031),
.B(n_1075),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1081),
.A2(n_1068),
.B1(n_1115),
.B2(n_1058),
.C(n_1118),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1057),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1077),
.B(n_1101),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1075),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1107),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1107),
.B(n_1045),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_1075),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1052),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1094),
.A2(n_1045),
.B(n_1047),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1032),
.A2(n_1109),
.B(n_1106),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1100),
.A2(n_717),
.B(n_929),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1010),
.A2(n_717),
.B(n_929),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1025),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_1028),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1002),
.A2(n_984),
.B(n_688),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1030),
.B(n_842),
.Y(n_1209)
);

OAI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1007),
.A2(n_545),
.B1(n_984),
.B2(n_993),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1091),
.A2(n_1086),
.B(n_1099),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1005),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1005),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1026),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1002),
.A2(n_984),
.B(n_1132),
.C(n_1129),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1026),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1053),
.B(n_957),
.Y(n_1217)
);

CKINVDCx11_ASAP7_75t_R g1218 ( 
.A(n_1020),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1015),
.A2(n_984),
.B(n_994),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1030),
.B(n_839),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1086),
.A2(n_1099),
.B(n_1129),
.Y(n_1221)
);

OAI22x1_ASAP7_75t_L g1222 ( 
.A1(n_1007),
.A2(n_545),
.B1(n_984),
.B2(n_993),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1223)
);

AND2x6_ASAP7_75t_L g1224 ( 
.A(n_1062),
.B(n_923),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1007),
.B(n_843),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1030),
.B(n_842),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1005),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1046),
.B(n_1085),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1007),
.B(n_843),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1046),
.B(n_1085),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1026),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1102),
.A2(n_1043),
.B(n_1078),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1013),
.Y(n_1237)
);

BUFx4_ASAP7_75t_SL g1238 ( 
.A(n_1037),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1025),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1020),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1130),
.B(n_1131),
.Y(n_1241)
);

O2A1O1Ixp5_ASAP7_75t_SL g1242 ( 
.A1(n_1132),
.A2(n_1040),
.B(n_1039),
.C(n_984),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1102),
.A2(n_1043),
.B(n_1078),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1053),
.B(n_957),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1026),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1011),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1053),
.A2(n_984),
.B1(n_962),
.B2(n_1084),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1008),
.A2(n_984),
.B1(n_363),
.B2(n_379),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1046),
.B(n_1085),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1053),
.B(n_957),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1013),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1030),
.B(n_842),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1053),
.A2(n_984),
.B1(n_962),
.B2(n_1084),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1013),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1048),
.A2(n_894),
.B(n_1093),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1053),
.A2(n_984),
.B1(n_962),
.B2(n_1084),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1013),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1008),
.A2(n_984),
.B1(n_363),
.B2(n_379),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1086),
.A2(n_1099),
.B(n_1129),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1053),
.B(n_957),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1247),
.B(n_1253),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1148),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1190),
.A2(n_1174),
.B(n_1208),
.C(n_1158),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1158),
.A2(n_1222),
.B1(n_1210),
.B2(n_1168),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_SL g1266 ( 
.A(n_1144),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1208),
.A2(n_1157),
.B(n_1169),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1192),
.B(n_1191),
.Y(n_1268)
);

OAI211xp5_ASAP7_75t_L g1269 ( 
.A1(n_1248),
.A2(n_1258),
.B(n_1169),
.C(n_1163),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1164),
.A2(n_1156),
.B(n_1146),
.C(n_1145),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1145),
.A2(n_1259),
.B(n_1221),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1200),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1242),
.B(n_1174),
.C(n_1215),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1154),
.A2(n_1230),
.B1(n_1225),
.B2(n_1156),
.C(n_1221),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1180),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1151),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1154),
.A2(n_1155),
.B1(n_1138),
.B2(n_1256),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1251),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1139),
.B(n_1229),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_1159),
.B(n_1152),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1136),
.A2(n_1139),
.B1(n_1244),
.B2(n_1260),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1235),
.A2(n_1243),
.B(n_1143),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1237),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1255),
.A2(n_1170),
.B(n_1204),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1219),
.A2(n_1181),
.B(n_1187),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1217),
.A2(n_1260),
.A3(n_1250),
.B(n_1244),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1171),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1237),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1136),
.B(n_1223),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1217),
.A2(n_1250),
.B(n_1193),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1194),
.B(n_1184),
.C(n_1220),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1218),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1139),
.A2(n_1162),
.B1(n_1241),
.B2(n_1231),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1246),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1227),
.B(n_1233),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1211),
.A2(n_1188),
.B(n_1177),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1161),
.B(n_1236),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1188),
.A2(n_1179),
.B(n_1202),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1203),
.A2(n_1196),
.B(n_1228),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1229),
.B(n_1232),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1196),
.A2(n_1172),
.B(n_1213),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1153),
.A2(n_1173),
.B1(n_1254),
.B2(n_1175),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1149),
.A2(n_1167),
.A3(n_1212),
.B(n_1153),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1182),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1167),
.Y(n_1305)
);

AOI22x1_ASAP7_75t_L g1306 ( 
.A1(n_1185),
.A2(n_1207),
.B1(n_1180),
.B2(n_1234),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1209),
.A2(n_1226),
.B1(n_1252),
.B2(n_1257),
.Y(n_1307)
);

NOR2x1_ASAP7_75t_R g1308 ( 
.A(n_1206),
.B(n_1239),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1178),
.A2(n_1183),
.B(n_1249),
.C(n_1232),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1199),
.A2(n_1198),
.B(n_1186),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1249),
.B(n_1224),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1166),
.A2(n_1197),
.B(n_1216),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1166),
.A2(n_1197),
.B(n_1216),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1189),
.A2(n_1224),
.B(n_1186),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1195),
.A2(n_1224),
.B(n_1234),
.Y(n_1315)
);

BUFx2_ASAP7_75t_R g1316 ( 
.A(n_1201),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1171),
.A2(n_1214),
.B(n_1245),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1171),
.B(n_1214),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1176),
.A2(n_1245),
.B(n_1165),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1176),
.B(n_1147),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1238),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1137),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1240),
.B(n_1136),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1161),
.B(n_1237),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1161),
.B(n_1237),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1225),
.B(n_984),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1225),
.B(n_984),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1210),
.A2(n_714),
.B(n_576),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1136),
.B(n_1223),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1158),
.A2(n_812),
.B1(n_984),
.B2(n_489),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1161),
.B(n_1237),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1145),
.A2(n_1259),
.B(n_1221),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1142),
.A2(n_1146),
.B(n_1152),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1238),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1140),
.Y(n_1339)
);

BUFx4f_ASAP7_75t_SL g1340 ( 
.A(n_1137),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1136),
.B(n_1223),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1169),
.A2(n_984),
.B(n_1002),
.C(n_1132),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1158),
.A2(n_1210),
.B1(n_1222),
.B2(n_1132),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1148),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1148),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1248),
.A2(n_984),
.B1(n_1258),
.B2(n_1136),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1148),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1158),
.A2(n_1210),
.B1(n_1222),
.B2(n_1132),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1238),
.Y(n_1349)
);

BUFx10_ASAP7_75t_L g1350 ( 
.A(n_1144),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1140),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1169),
.A2(n_984),
.B(n_1002),
.C(n_1132),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1248),
.A2(n_984),
.B1(n_363),
.B2(n_379),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1158),
.A2(n_1210),
.B1(n_1222),
.B2(n_1132),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1225),
.B(n_984),
.Y(n_1356)
);

OAI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1248),
.A2(n_984),
.B1(n_538),
.B2(n_550),
.C(n_688),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1161),
.B(n_1237),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_L g1360 ( 
.A(n_1158),
.B(n_984),
.C(n_688),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1248),
.A2(n_984),
.B1(n_1258),
.B2(n_812),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1237),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1150),
.A2(n_1141),
.B(n_1205),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_1147),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1248),
.A2(n_984),
.B1(n_363),
.B2(n_379),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1140),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1279),
.B(n_1301),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1283),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1270),
.A2(n_1290),
.B(n_1274),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1357),
.A2(n_1361),
.B(n_1346),
.C(n_1342),
.Y(n_1370)
);

OA22x2_ASAP7_75t_L g1371 ( 
.A1(n_1269),
.A2(n_1293),
.B1(n_1323),
.B2(n_1341),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1326),
.A2(n_1327),
.B1(n_1356),
.B2(n_1265),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1297),
.B(n_1326),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1279),
.B(n_1301),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1327),
.B(n_1356),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1289),
.B(n_1329),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1304),
.B(n_1307),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1330),
.A2(n_1265),
.B1(n_1355),
.B2(n_1348),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1307),
.B(n_1300),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1324),
.B(n_1325),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1270),
.A2(n_1290),
.B(n_1309),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1332),
.B(n_1358),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1295),
.B(n_1302),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_R g1384 ( 
.A(n_1337),
.B(n_1349),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1353),
.A2(n_1365),
.B1(n_1291),
.B2(n_1360),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1302),
.B(n_1281),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1309),
.A2(n_1352),
.B(n_1342),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1279),
.B(n_1343),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1343),
.B(n_1348),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1314),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1336),
.A2(n_1280),
.B(n_1273),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1288),
.B(n_1355),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1264),
.A2(n_1352),
.B(n_1267),
.C(n_1261),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1362),
.B(n_1286),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1285),
.A2(n_1262),
.B(n_1363),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1292),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1277),
.A2(n_1345),
.B1(n_1347),
.B2(n_1344),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1277),
.A2(n_1345),
.B1(n_1347),
.B2(n_1328),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1286),
.B(n_1263),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1272),
.B(n_1320),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1272),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1276),
.B(n_1278),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1303),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1271),
.A2(n_1333),
.B(n_1311),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1331),
.A2(n_1335),
.B(n_1359),
.Y(n_1405)
);

AND2x2_ASAP7_75t_SL g1406 ( 
.A(n_1305),
.B(n_1311),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1337),
.Y(n_1407)
);

AND2x6_ASAP7_75t_L g1408 ( 
.A(n_1311),
.B(n_1294),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1294),
.B(n_1366),
.Y(n_1409)
);

OAI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1272),
.A2(n_1306),
.B1(n_1321),
.B2(n_1351),
.C(n_1339),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1268),
.A2(n_1314),
.B(n_1317),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_1316),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1268),
.A2(n_1364),
.B1(n_1266),
.B2(n_1275),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1299),
.B(n_1318),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1318),
.B(n_1299),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1275),
.A2(n_1349),
.B1(n_1292),
.B2(n_1340),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1315),
.B(n_1296),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1296),
.B(n_1298),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1298),
.B(n_1319),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1334),
.A2(n_1354),
.B(n_1338),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1322),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1308),
.A2(n_1317),
.B(n_1287),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1350),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1312),
.B(n_1313),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1284),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1282),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1326),
.A2(n_1356),
.B1(n_1327),
.B2(n_1357),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1326),
.A2(n_1356),
.B1(n_1327),
.B2(n_1357),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1324),
.B(n_1325),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1270),
.A2(n_984),
.B(n_785),
.Y(n_1431)
);

AOI21xp33_ASAP7_75t_L g1432 ( 
.A1(n_1360),
.A2(n_984),
.B(n_1264),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1326),
.A2(n_1356),
.B1(n_1327),
.B2(n_1357),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1324),
.B(n_1325),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1326),
.A2(n_1356),
.B1(n_1327),
.B2(n_1357),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1367),
.B(n_1374),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1403),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1422),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1394),
.B(n_1393),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1416),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1381),
.B(n_1369),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1399),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1390),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1372),
.B(n_1428),
.Y(n_1444)
);

CKINVDCx8_ASAP7_75t_R g1445 ( 
.A(n_1408),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1381),
.B(n_1369),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1373),
.B(n_1375),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1418),
.B(n_1367),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1370),
.A2(n_1385),
.B(n_1433),
.Y(n_1449)
);

CKINVDCx16_ASAP7_75t_R g1450 ( 
.A(n_1384),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1419),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1425),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1374),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1420),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1391),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1414),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1383),
.B(n_1429),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1391),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1391),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1408),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1392),
.B(n_1426),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1427),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1435),
.B(n_1377),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1432),
.A2(n_1378),
.B1(n_1387),
.B2(n_1389),
.C(n_1386),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1415),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1411),
.A2(n_1404),
.B(n_1387),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1395),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1409),
.Y(n_1468)
);

NAND2x1_ASAP7_75t_L g1469 ( 
.A(n_1441),
.B(n_1431),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1443),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_1455),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1462),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1443),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1368),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1462),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1454),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1462),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1454),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_SL g1479 ( 
.A(n_1441),
.B(n_1413),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1456),
.B(n_1368),
.Y(n_1480)
);

INVx5_ASAP7_75t_SL g1481 ( 
.A(n_1441),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1438),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1442),
.B(n_1380),
.Y(n_1483)
);

AND2x2_ASAP7_75t_SL g1484 ( 
.A(n_1441),
.B(n_1406),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1460),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1451),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1444),
.B(n_1371),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1437),
.Y(n_1488)
);

NOR4xp25_ASAP7_75t_SL g1489 ( 
.A(n_1464),
.B(n_1410),
.C(n_1449),
.D(n_1407),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1448),
.B(n_1405),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1448),
.B(n_1405),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1444),
.A2(n_1371),
.B1(n_1379),
.B2(n_1398),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1452),
.B(n_1421),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1487),
.B(n_1450),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1487),
.A2(n_1464),
.B1(n_1457),
.B2(n_1463),
.C(n_1439),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1472),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1492),
.A2(n_1457),
.B1(n_1463),
.B2(n_1439),
.C(n_1456),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1492),
.A2(n_1441),
.B1(n_1446),
.B2(n_1445),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1486),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1472),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1483),
.B(n_1468),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1471),
.A2(n_1459),
.B(n_1455),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1485),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1484),
.A2(n_1446),
.B1(n_1441),
.B2(n_1466),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1482),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1469),
.A2(n_1441),
.B1(n_1446),
.B2(n_1447),
.C(n_1400),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1484),
.A2(n_1446),
.B1(n_1388),
.B2(n_1466),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1482),
.Y(n_1510)
);

AND3x1_ASAP7_75t_L g1511 ( 
.A(n_1489),
.B(n_1450),
.C(n_1402),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1440),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1470),
.Y(n_1513)
);

AOI21xp33_ASAP7_75t_L g1514 ( 
.A1(n_1474),
.A2(n_1446),
.B(n_1461),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1489),
.B(n_1446),
.C(n_1376),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1475),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1483),
.B(n_1465),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1477),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1470),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1484),
.A2(n_1466),
.B1(n_1481),
.B2(n_1436),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1488),
.Y(n_1521)
);

OAI211xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1480),
.A2(n_1382),
.B(n_1434),
.C(n_1430),
.Y(n_1522)
);

NOR4xp25_ASAP7_75t_SL g1523 ( 
.A(n_1471),
.B(n_1453),
.C(n_1467),
.D(n_1407),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1490),
.B(n_1436),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1478),
.B(n_1452),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1507),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1506),
.B(n_1484),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1521),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1505),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1507),
.B(n_1478),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1505),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1498),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1502),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1501),
.B(n_1486),
.Y(n_1537)
);

BUFx8_ASAP7_75t_L g1538 ( 
.A(n_1507),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1504),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1504),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1501),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1513),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1494),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1473),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1501),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1516),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1519),
.A2(n_1493),
.B(n_1458),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1518),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1518),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1538),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1548),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1545),
.B(n_1525),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1526),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1537),
.B(n_1524),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1545),
.B(n_1524),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1526),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1479),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_R g1560 ( 
.A(n_1530),
.B(n_1384),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1496),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1529),
.B(n_1479),
.Y(n_1562)
);

NAND5xp2_ASAP7_75t_SL g1563 ( 
.A(n_1538),
.B(n_1508),
.C(n_1499),
.D(n_1520),
.E(n_1509),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1528),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1548),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1526),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1537),
.B(n_1501),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1533),
.B(n_1479),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1550),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1537),
.B(n_1512),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1551),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1533),
.B(n_1503),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1538),
.B(n_1511),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1551),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1527),
.B(n_1417),
.C(n_1515),
.Y(n_1576)
);

AOI211x1_ASAP7_75t_SL g1577 ( 
.A1(n_1527),
.A2(n_1515),
.B(n_1500),
.C(n_1495),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1538),
.A2(n_1510),
.B1(n_1466),
.B2(n_1522),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1532),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1532),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1535),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1535),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1541),
.B(n_1517),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1531),
.B(n_1512),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1536),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1576),
.A2(n_1511),
.B1(n_1538),
.B2(n_1530),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1561),
.B(n_1526),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1561),
.B(n_1510),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1552),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1564),
.Y(n_1591)
);

INVx3_ASAP7_75t_SL g1592 ( 
.A(n_1558),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1552),
.B(n_1531),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1573),
.B(n_1541),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1576),
.A2(n_1510),
.B1(n_1523),
.B2(n_1484),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1564),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1558),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1573),
.B(n_1546),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1584),
.B(n_1539),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_SL g1602 ( 
.A(n_1577),
.B(n_1543),
.C(n_1539),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1569),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1558),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1558),
.B(n_1547),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1546),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1579),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1579),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1555),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1566),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1556),
.B(n_1539),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1543),
.Y(n_1613)
);

NAND4xp25_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1514),
.C(n_1397),
.D(n_1543),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1580),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1556),
.B(n_1547),
.Y(n_1616)
);

AO32x1_ASAP7_75t_L g1617 ( 
.A1(n_1563),
.A2(n_1540),
.A3(n_1542),
.B1(n_1534),
.B2(n_1544),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1581),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1557),
.B(n_1491),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1560),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1581),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1396),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1587),
.A2(n_1578),
.B1(n_1574),
.B2(n_1563),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1609),
.B(n_1554),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1600),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1593),
.B(n_1559),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1559),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1610),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1592),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1610),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1589),
.B(n_1422),
.Y(n_1633)
);

AOI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1596),
.A2(n_1578),
.B1(n_1562),
.B2(n_1568),
.C1(n_1565),
.C2(n_1572),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1594),
.B(n_1601),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1622),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1592),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1594),
.B(n_1562),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1588),
.Y(n_1639)
);

INVx3_ASAP7_75t_SL g1640 ( 
.A(n_1598),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1622),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1591),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1607),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1611),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1604),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1611),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1396),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1601),
.B(n_1568),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1624),
.A2(n_1623),
.B1(n_1647),
.B2(n_1621),
.Y(n_1649)
);

AOI211xp5_ASAP7_75t_L g1650 ( 
.A1(n_1637),
.A2(n_1590),
.B(n_1617),
.C(n_1614),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1623),
.A2(n_1617),
.B1(n_1424),
.B2(n_1597),
.Y(n_1651)
);

OAI311xp33_ASAP7_75t_L g1652 ( 
.A1(n_1634),
.A2(n_1617),
.A3(n_1603),
.B1(n_1606),
.C1(n_1599),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1631),
.B(n_1612),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1626),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1647),
.A2(n_1617),
.B(n_1615),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1631),
.B(n_1612),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1639),
.A2(n_1595),
.B1(n_1613),
.B2(n_1618),
.C(n_1608),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1630),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1625),
.A2(n_1554),
.B1(n_1620),
.B2(n_1485),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1635),
.A2(n_1613),
.B1(n_1616),
.B2(n_1605),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1645),
.B(n_1557),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1625),
.B(n_1583),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1664)
);

AOI222xp33_ASAP7_75t_L g1665 ( 
.A1(n_1642),
.A2(n_1565),
.B1(n_1570),
.B2(n_1553),
.C1(n_1572),
.C2(n_1575),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1632),
.B(n_1611),
.Y(n_1666)
);

OAI322xp33_ASAP7_75t_L g1667 ( 
.A1(n_1629),
.A2(n_1553),
.A3(n_1575),
.B1(n_1570),
.B2(n_1542),
.C1(n_1540),
.C2(n_1534),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1633),
.B(n_1605),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1632),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1654),
.B(n_1632),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1657),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1653),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1650),
.B(n_1629),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1666),
.B(n_1640),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1655),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1661),
.B(n_1627),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1664),
.B(n_1640),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1627),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1662),
.B(n_1628),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1640),
.Y(n_1680)
);

NAND4xp25_ASAP7_75t_L g1681 ( 
.A(n_1680),
.B(n_1658),
.C(n_1656),
.D(n_1665),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1673),
.A2(n_1652),
.B(n_1651),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1669),
.B(n_1656),
.C(n_1626),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1671),
.B(n_1663),
.C(n_1642),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1671),
.B(n_1628),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1678),
.B(n_1644),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1670),
.A2(n_1677),
.B(n_1674),
.C(n_1675),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_L g1688 ( 
.A1(n_1676),
.A2(n_1646),
.B(n_1644),
.C(n_1643),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1679),
.A2(n_1667),
.B(n_1660),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1672),
.Y(n_1690)
);

AOI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1673),
.A2(n_1643),
.B1(n_1641),
.B2(n_1636),
.C1(n_1646),
.C2(n_1644),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1673),
.A2(n_1648),
.B1(n_1638),
.B2(n_1646),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1684),
.A2(n_1641),
.B(n_1636),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1685),
.Y(n_1694)
);

NOR2x1p5_ASAP7_75t_L g1695 ( 
.A(n_1686),
.B(n_1681),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1682),
.B(n_1638),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_R g1697 ( 
.A(n_1690),
.B(n_1424),
.Y(n_1697)
);

OAI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1683),
.A2(n_1648),
.B1(n_1547),
.B2(n_1585),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1688),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1694),
.Y(n_1700)
);

INVxp67_ASAP7_75t_SL g1701 ( 
.A(n_1693),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1697),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1699),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1696),
.B(n_1691),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1695),
.B(n_1692),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1698),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1700),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_R g1708 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1703),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1702),
.B(n_1689),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1705),
.B(n_1605),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1711),
.B(n_1704),
.C(n_1706),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1710),
.A2(n_1705),
.B1(n_1701),
.B2(n_1616),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1707),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1713),
.Y(n_1715)
);

AOI22x1_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1709),
.B1(n_1714),
.B2(n_1708),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1716),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1716),
.A2(n_1712),
.B1(n_1567),
.B2(n_1571),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1717),
.A2(n_1412),
.B1(n_1401),
.B2(n_1567),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1718),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1720),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1719),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1721),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1724),
.B(n_1722),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1725),
.A2(n_1567),
.B(n_1582),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1586),
.B1(n_1582),
.B2(n_1567),
.C(n_1585),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1727),
.A2(n_1423),
.B(n_1586),
.C(n_1542),
.Y(n_1728)
);


endmodule