module fake_jpeg_7193_n_109 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

OR2x4_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_23),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_17),
.C(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_21),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_17),
.B(n_24),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_48),
.B(n_31),
.C(n_12),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_24),
.B1(n_23),
.B2(n_15),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_46),
.B1(n_16),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_15),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_43),
.B1(n_40),
.B2(n_27),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_16),
.B1(n_1),
.B2(n_0),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_71),
.B(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_71)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_52),
.B(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_68),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_61),
.B(n_27),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_63),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_27),
.B(n_34),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_33),
.B(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22x1_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_69),
.B1(n_65),
.B2(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_89),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_90),
.B(n_92),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_68),
.C(n_69),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_69),
.C(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_62),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_87),
.B(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_65),
.B1(n_74),
.B2(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_37),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_100),
.C(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_93),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_35),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_104),
.B(n_103),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_97),
.C(n_5),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.C(n_11),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_6),
.CI(n_7),
.CON(n_106),
.SN(n_106)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_6),
.B(n_7),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_8),
.Y(n_109)
);


endmodule