module fake_jpeg_28058_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_74),
.Y(n_90)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_0),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_61),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_63),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_66),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_56),
.B(n_69),
.C(n_59),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_65),
.B1(n_68),
.B2(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_66),
.B1(n_62),
.B2(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_65),
.B1(n_55),
.B2(n_57),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_68),
.B1(n_67),
.B2(n_50),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_51),
.B1(n_52),
.B2(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_54),
.B1(n_58),
.B2(n_57),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_104),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_105),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_78),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_53),
.C(n_62),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_58),
.B1(n_57),
.B2(n_61),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_109),
.B1(n_80),
.B2(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_1),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_110),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_80),
.B(n_85),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_109),
.B1(n_100),
.B2(n_94),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_21),
.B(n_27),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_116),
.B(n_31),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_106),
.B(n_98),
.C(n_95),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_96),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_124),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_96),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_133),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_15),
.B(n_46),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_118),
.C(n_116),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_101),
.C(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_144),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_17),
.B(n_13),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_1),
.CI(n_2),
.CON(n_140),
.SN(n_140)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_16),
.B1(n_45),
.B2(n_44),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_48),
.C(n_42),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_40),
.C(n_38),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_143),
.B1(n_7),
.B2(n_8),
.Y(n_158)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_28),
.B(n_24),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_156),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_139),
.B1(n_134),
.B2(n_140),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_135),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_149),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_135),
.C(n_159),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_148),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_160),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_151),
.C(n_162),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_6),
.B(n_8),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_9),
.B(n_10),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_159),
.Y(n_173)
);


endmodule