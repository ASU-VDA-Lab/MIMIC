module real_jpeg_30788_n_13 (n_123, n_8, n_116, n_0, n_2, n_114, n_10, n_9, n_12, n_6, n_121, n_11, n_120, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_113, n_13);

input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_114;
input n_10;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_120;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_113;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI221x1_ASAP7_75t_L g37 ( 
.A1(n_0),
.A2(n_7),
.B1(n_38),
.B2(n_45),
.C(n_48),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_38),
.C(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_2),
.B(n_103),
.CON(n_102),
.SN(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_5),
.B(n_95),
.Y(n_107)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_76),
.A3(n_78),
.B1(n_82),
.B2(n_106),
.C1(n_108),
.C2(n_123),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B1(n_16),
.B2(n_22),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_23),
.Y(n_13)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI31xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_70),
.A3(n_93),
.B(n_100),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_61),
.C(n_62),
.Y(n_26)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_52),
.B(n_60),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_34),
.B(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_115),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_81),
.C(n_90),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_101),
.B(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_90),
.C(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_119),
.Y(n_78)
);

OA21x2_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_113),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_114),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_116),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_117),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_118),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_120),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_121),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_122),
.Y(n_96)
);


endmodule