module real_aes_18066_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_1280;
wire n_729;
wire n_394;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g1040 ( .A(n_0), .Y(n_1040) );
AOI221x1_ASAP7_75t_SL g1052 ( .A1(n_0), .A2(n_2), .B1(n_1053), .B2(n_1054), .C(n_1055), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_1), .A2(n_6), .B1(n_1283), .B2(n_1286), .Y(n_1296) );
XOR2xp5_ASAP7_75t_L g1486 ( .A(n_1), .B(n_1487), .Y(n_1486) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_1), .A2(n_1533), .B1(n_1538), .B2(n_1579), .Y(n_1532) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_2), .A2(n_22), .B1(n_554), .B2(n_576), .Y(n_1047) );
INVx1_ASAP7_75t_L g1547 ( .A(n_3), .Y(n_1547) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_4), .A2(n_410), .B(n_420), .C(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g470 ( .A(n_4), .Y(n_470) );
INVx1_ASAP7_75t_L g619 ( .A(n_5), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g665 ( .A1(n_5), .A2(n_666), .B(n_668), .C(n_677), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_7), .A2(n_44), .B1(n_1053), .B2(n_1497), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_7), .A2(n_223), .B1(n_580), .B2(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g868 ( .A(n_8), .Y(n_868) );
INVx1_ASAP7_75t_L g571 ( .A(n_9), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_9), .A2(n_115), .B1(n_607), .B2(n_609), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_10), .A2(n_216), .B1(n_967), .B2(n_970), .C(n_971), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_10), .A2(n_216), .B1(n_991), .B2(n_992), .Y(n_990) );
INVxp67_ASAP7_75t_SL g934 ( .A(n_11), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_11), .A2(n_28), .B1(n_552), .B2(n_676), .Y(n_944) );
INVx1_ASAP7_75t_L g965 ( .A(n_12), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_12), .A2(n_269), .B1(n_505), .B2(n_985), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_13), .A2(n_263), .B1(n_672), .B2(n_911), .C(n_960), .Y(n_959) );
AOI222xp33_ASAP7_75t_L g999 ( .A1(n_13), .A2(n_70), .B1(n_151), .B2(n_393), .C1(n_603), .C2(n_1000), .Y(n_999) );
AOI21xp33_ASAP7_75t_L g1046 ( .A1(n_14), .A2(n_573), .B(n_574), .Y(n_1046) );
INVx1_ASAP7_75t_L g1062 ( .A(n_14), .Y(n_1062) );
INVx1_ASAP7_75t_L g294 ( .A(n_15), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_15), .B(n_304), .Y(n_318) );
AND2x2_ASAP7_75t_L g502 ( .A(n_15), .B(n_449), .Y(n_502) );
AND2x2_ASAP7_75t_L g569 ( .A(n_15), .B(n_237), .Y(n_569) );
INVx1_ASAP7_75t_L g1074 ( .A(n_16), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1109 ( .A1(n_16), .A2(n_635), .B(n_880), .C(n_1110), .Y(n_1109) );
OAI211xp5_ASAP7_75t_L g831 ( .A1(n_17), .A2(n_832), .B(n_833), .C(n_838), .Y(n_831) );
INVx1_ASAP7_75t_L g844 ( .A(n_17), .Y(n_844) );
INVx1_ASAP7_75t_L g1126 ( .A(n_18), .Y(n_1126) );
INVx1_ASAP7_75t_L g1139 ( .A(n_19), .Y(n_1139) );
INVx2_ASAP7_75t_L g1279 ( .A(n_20), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_20), .B(n_112), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_20), .B(n_1285), .Y(n_1287) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_21), .A2(n_164), .B1(n_823), .B2(n_825), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_21), .A2(n_164), .B1(n_846), .B2(n_847), .Y(n_845) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_22), .A2(n_180), .B1(n_1054), .B2(n_1058), .C(n_1060), .Y(n_1057) );
INVx1_ASAP7_75t_L g1202 ( .A(n_23), .Y(n_1202) );
INVx1_ASAP7_75t_L g784 ( .A(n_24), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g1312 ( .A1(n_25), .A2(n_244), .B1(n_1283), .B2(n_1286), .Y(n_1312) );
OAI21xp5_ASAP7_75t_L g1522 ( .A1(n_26), .A2(n_1523), .B(n_1524), .Y(n_1522) );
OAI22xp33_ASAP7_75t_L g829 ( .A1(n_27), .A2(n_42), .B1(n_296), .B2(n_830), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_27), .A2(n_42), .B1(n_758), .B2(n_841), .Y(n_840) );
INVxp67_ASAP7_75t_SL g927 ( .A(n_28), .Y(n_927) );
INVx1_ASAP7_75t_L g1204 ( .A(n_29), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_30), .A2(n_198), .B1(n_398), .B2(n_1245), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_30), .A2(n_129), .B1(n_962), .B2(n_1255), .Y(n_1265) );
INVx1_ASAP7_75t_L g1520 ( .A(n_31), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_32), .A2(n_129), .B1(n_398), .B2(n_1245), .Y(n_1244) );
AOI22xp33_ASAP7_75t_SL g1258 ( .A1(n_32), .A2(n_198), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1506 ( .A(n_33), .Y(n_1506) );
INVx1_ASAP7_75t_L g912 ( .A(n_34), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_35), .A2(n_186), .B1(n_415), .B2(n_416), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_35), .A2(n_186), .B1(n_296), .B2(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g486 ( .A(n_36), .Y(n_486) );
INVx1_ASAP7_75t_L g1094 ( .A(n_37), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g1301 ( .A1(n_38), .A2(n_272), .B1(n_1276), .B2(n_1302), .Y(n_1301) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_39), .A2(n_245), .B1(n_654), .B2(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g669 ( .A(n_39), .Y(n_669) );
INVx1_ASAP7_75t_L g867 ( .A(n_40), .Y(n_867) );
INVx1_ASAP7_75t_L g347 ( .A(n_41), .Y(n_347) );
INVx1_ASAP7_75t_L g1073 ( .A(n_43), .Y(n_1073) );
AOI221xp5_ASAP7_75t_L g1510 ( .A1(n_44), .A2(n_124), .B1(n_547), .B2(n_680), .C(n_975), .Y(n_1510) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_45), .A2(n_166), .B1(n_830), .B2(n_916), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_45), .A2(n_166), .B1(n_1106), .B2(n_1108), .Y(n_1105) );
INVx1_ASAP7_75t_L g750 ( .A(n_46), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_47), .A2(n_254), .B1(n_1283), .B2(n_1286), .Y(n_1305) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_48), .A2(n_119), .B1(n_643), .B2(n_645), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_48), .A2(n_245), .B1(n_675), .B2(n_676), .Y(n_681) );
AO22x1_ASAP7_75t_L g1309 ( .A1(n_49), .A2(n_65), .B1(n_1276), .B2(n_1291), .Y(n_1309) );
INVx1_ASAP7_75t_L g929 ( .A(n_50), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_50), .A2(n_136), .B1(n_940), .B2(n_942), .Y(n_939) );
OAI22xp5_ASAP7_75t_SL g1029 ( .A1(n_51), .A2(n_182), .B1(n_537), .B2(n_541), .Y(n_1029) );
INVx1_ASAP7_75t_L g1033 ( .A(n_51), .Y(n_1033) );
OAI211xp5_ASAP7_75t_L g1565 ( .A1(n_52), .A2(n_420), .B(n_1566), .C(n_1568), .Y(n_1565) );
INVx1_ASAP7_75t_L g1575 ( .A(n_52), .Y(n_1575) );
AOI22xp33_ASAP7_75t_SL g1499 ( .A1(n_53), .A2(n_116), .B1(n_644), .B2(n_1251), .Y(n_1499) );
AOI221xp5_ASAP7_75t_L g1514 ( .A1(n_53), .A2(n_83), .B1(n_672), .B2(n_976), .C(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g863 ( .A(n_54), .Y(n_863) );
INVx1_ASAP7_75t_L g377 ( .A(n_55), .Y(n_377) );
INVx1_ASAP7_75t_L g383 ( .A(n_55), .Y(n_383) );
INVx1_ASAP7_75t_L g323 ( .A(n_56), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_57), .A2(n_484), .B1(n_612), .B2(n_613), .Y(n_483) );
INVxp67_ASAP7_75t_L g613 ( .A(n_57), .Y(n_613) );
INVx1_ASAP7_75t_L g652 ( .A(n_58), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_58), .A2(n_251), .B1(n_675), .B2(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g707 ( .A(n_59), .Y(n_707) );
INVxp67_ASAP7_75t_SL g973 ( .A(n_60), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_60), .A2(n_263), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
INVx1_ASAP7_75t_L g786 ( .A(n_61), .Y(n_786) );
INVx1_ASAP7_75t_L g1163 ( .A(n_62), .Y(n_1163) );
INVx1_ASAP7_75t_L g1519 ( .A(n_63), .Y(n_1519) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_64), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_65), .A2(n_615), .B1(n_616), .B2(n_696), .Y(n_614) );
INVxp67_ASAP7_75t_L g696 ( .A(n_65), .Y(n_696) );
INVx1_ASAP7_75t_L g287 ( .A(n_66), .Y(n_287) );
INVx1_ASAP7_75t_L g1552 ( .A(n_67), .Y(n_1552) );
INVx2_ASAP7_75t_L g369 ( .A(n_68), .Y(n_369) );
INVx1_ASAP7_75t_L g1208 ( .A(n_69), .Y(n_1208) );
AOI22xp33_ASAP7_75t_SL g961 ( .A1(n_70), .A2(n_163), .B1(n_940), .B2(n_962), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_71), .A2(n_162), .B1(n_830), .B2(n_916), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_71), .A2(n_162), .B1(n_416), .B2(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g910 ( .A(n_72), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_73), .A2(n_278), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g591 ( .A(n_73), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g1306 ( .A1(n_74), .A2(n_188), .B1(n_1276), .B2(n_1291), .Y(n_1306) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_75), .A2(n_79), .B1(n_296), .B2(n_446), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_75), .A2(n_79), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g874 ( .A(n_76), .Y(n_874) );
AO221x2_ASAP7_75t_L g1348 ( .A1(n_77), .A2(n_230), .B1(n_1283), .B2(n_1286), .C(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1549 ( .A(n_78), .Y(n_1549) );
INVx1_ASAP7_75t_L g1124 ( .A(n_80), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_81), .A2(n_271), .B1(n_823), .B2(n_827), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_81), .A2(n_111), .B1(n_841), .B2(n_846), .Y(n_1190) );
OAI211xp5_ASAP7_75t_L g1071 ( .A1(n_82), .A2(n_747), .B(n_938), .C(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1111 ( .A(n_82), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_83), .A2(n_238), .B1(n_609), .B2(n_1495), .Y(n_1494) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_84), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_84), .A2(n_219), .B1(n_684), .B2(n_685), .C(n_688), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_85), .A2(n_115), .B1(n_552), .B2(n_554), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_85), .A2(n_197), .B1(n_593), .B2(n_596), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g804 ( .A1(n_86), .A2(n_746), .B(n_747), .C(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g816 ( .A(n_86), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_87), .A2(n_183), .B1(n_472), .B2(n_474), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g817 ( .A1(n_87), .A2(n_183), .B1(n_436), .B2(n_765), .Y(n_817) );
INVx1_ASAP7_75t_L g837 ( .A(n_88), .Y(n_837) );
OAI211xp5_ASAP7_75t_L g842 ( .A1(n_88), .A2(n_410), .B(n_635), .C(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g1128 ( .A(n_89), .Y(n_1128) );
XOR2x2_ASAP7_75t_L g818 ( .A(n_90), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g432 ( .A(n_91), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_91), .A2(n_453), .B(n_455), .C(n_461), .Y(n_452) );
INVx1_ASAP7_75t_L g1011 ( .A(n_92), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_93), .A2(n_101), .B1(n_841), .B2(n_1160), .Y(n_1159) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_93), .A2(n_117), .B1(n_296), .B2(n_1169), .Y(n_1168) );
INVx1_ASAP7_75t_L g705 ( .A(n_94), .Y(n_705) );
OAI221xp5_ASAP7_75t_SL g521 ( .A1(n_95), .A2(n_99), .B1(n_522), .B2(n_528), .C(n_534), .Y(n_521) );
INVx1_ASAP7_75t_L g564 ( .A(n_95), .Y(n_564) );
INVx1_ASAP7_75t_L g353 ( .A(n_96), .Y(n_353) );
INVx1_ASAP7_75t_L g1044 ( .A(n_97), .Y(n_1044) );
INVx1_ASAP7_75t_L g352 ( .A(n_98), .Y(n_352) );
INVx1_ASAP7_75t_L g582 ( .A(n_99), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_100), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_101), .A2(n_174), .B1(n_823), .B2(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1228 ( .A(n_102), .Y(n_1228) );
XNOR2xp5_ASAP7_75t_L g1180 ( .A(n_103), .B(n_1181), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_104), .A2(n_1068), .B1(n_1069), .B2(n_1114), .Y(n_1067) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_104), .Y(n_1114) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_105), .Y(n_289) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_105), .B(n_287), .Y(n_1277) );
OAI211xp5_ASAP7_75t_SL g955 ( .A1(n_106), .A2(n_956), .B(n_958), .C(n_963), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_106), .A2(n_217), .B1(n_488), .B2(n_982), .Y(n_981) );
XNOR2xp5_ASAP7_75t_L g953 ( .A(n_107), .B(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g1232 ( .A(n_108), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_108), .A2(n_265), .B1(n_1237), .B2(n_1238), .Y(n_1236) );
INVx1_ASAP7_75t_L g714 ( .A(n_109), .Y(n_714) );
INVx1_ASAP7_75t_L g1140 ( .A(n_110), .Y(n_1140) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_111), .A2(n_173), .B1(n_296), .B2(n_446), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_112), .B(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1285 ( .A(n_112), .Y(n_1285) );
INVx1_ASAP7_75t_L g1233 ( .A(n_113), .Y(n_1233) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_114), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_116), .A2(n_238), .B1(n_577), .B2(n_1034), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_117), .A2(n_174), .B1(n_847), .B2(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g512 ( .A(n_118), .Y(n_512) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_119), .A2(n_574), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g718 ( .A(n_120), .Y(n_718) );
INVx2_ASAP7_75t_L g368 ( .A(n_121), .Y(n_368) );
INVx1_ASAP7_75t_L g408 ( .A(n_121), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_121), .B(n_369), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_122), .A2(n_249), .B1(n_434), .B2(n_436), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_122), .A2(n_249), .B1(n_472), .B2(n_474), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_123), .A2(n_225), .B1(n_1276), .B2(n_1291), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_124), .A2(n_223), .B1(n_1053), .B2(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1225 ( .A(n_125), .Y(n_1225) );
INVx1_ASAP7_75t_L g1082 ( .A(n_126), .Y(n_1082) );
AOI22xp33_ASAP7_75t_SL g1243 ( .A1(n_127), .A2(n_153), .B1(n_998), .B2(n_1000), .Y(n_1243) );
AOI22xp33_ASAP7_75t_SL g1262 ( .A1(n_127), .A2(n_229), .B1(n_1259), .B2(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g807 ( .A(n_128), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g1564 ( .A1(n_130), .A2(n_187), .B1(n_841), .B2(n_1160), .Y(n_1564) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_130), .A2(n_258), .B1(n_472), .B2(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g913 ( .A(n_131), .Y(n_913) );
INVx1_ASAP7_75t_L g1206 ( .A(n_132), .Y(n_1206) );
INVx1_ASAP7_75t_L g774 ( .A(n_133), .Y(n_774) );
INVx1_ASAP7_75t_L g1186 ( .A(n_134), .Y(n_1186) );
OAI211xp5_ASAP7_75t_L g1191 ( .A1(n_134), .A2(n_420), .B(n_725), .C(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1569 ( .A(n_135), .Y(n_1569) );
INVxp67_ASAP7_75t_SL g921 ( .A(n_136), .Y(n_921) );
XOR2xp5_ASAP7_75t_L g1539 ( .A(n_137), .B(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g633 ( .A(n_138), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_138), .A2(n_171), .B1(n_662), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g1090 ( .A(n_139), .Y(n_1090) );
OAI211xp5_ASAP7_75t_L g1183 ( .A1(n_140), .A2(n_832), .B(n_838), .C(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1193 ( .A(n_140), .Y(n_1193) );
INVx1_ASAP7_75t_L g1019 ( .A(n_141), .Y(n_1019) );
INVx1_ASAP7_75t_L g775 ( .A(n_142), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g745 ( .A1(n_143), .A2(n_746), .B(n_747), .C(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g763 ( .A(n_143), .Y(n_763) );
INVx1_ASAP7_75t_L g782 ( .A(n_144), .Y(n_782) );
INVx1_ASAP7_75t_L g1211 ( .A(n_145), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_146), .Y(n_650) );
INVx1_ASAP7_75t_L g330 ( .A(n_147), .Y(n_330) );
INVx1_ASAP7_75t_L g336 ( .A(n_148), .Y(n_336) );
INVx1_ASAP7_75t_L g640 ( .A(n_149), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_149), .A2(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g873 ( .A(n_150), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_151), .A2(n_228), .B1(n_975), .B2(n_976), .C(n_977), .Y(n_974) );
INVx1_ASAP7_75t_L g1135 ( .A(n_152), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_153), .A2(n_276), .B1(n_1255), .B2(n_1256), .Y(n_1254) );
CKINVDCx5p33_ASAP7_75t_R g1490 ( .A(n_154), .Y(n_1490) );
INVx1_ASAP7_75t_L g1555 ( .A(n_155), .Y(n_1555) );
OAI22xp33_ASAP7_75t_L g803 ( .A1(n_156), .A2(n_256), .B1(n_296), .B2(n_446), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_156), .A2(n_256), .B1(n_757), .B2(n_813), .Y(n_812) );
AO22x1_ASAP7_75t_L g1310 ( .A1(n_157), .A2(n_242), .B1(n_1283), .B2(n_1286), .Y(n_1310) );
INVx1_ASAP7_75t_L g1550 ( .A(n_158), .Y(n_1550) );
BUFx3_ASAP7_75t_L g375 ( .A(n_159), .Y(n_375) );
INVx1_ASAP7_75t_L g1093 ( .A(n_160), .Y(n_1093) );
INVx1_ASAP7_75t_L g1556 ( .A(n_161), .Y(n_1556) );
INVx1_ASAP7_75t_L g1006 ( .A(n_163), .Y(n_1006) );
INVx1_ASAP7_75t_L g922 ( .A(n_165), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_167), .A2(n_179), .B1(n_1283), .B2(n_1286), .Y(n_1292) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_168), .Y(n_301) );
INVx1_ASAP7_75t_L g496 ( .A(n_169), .Y(n_496) );
INVx1_ASAP7_75t_L g1201 ( .A(n_170), .Y(n_1201) );
INVx1_ASAP7_75t_L g631 ( .A(n_171), .Y(n_631) );
INVx1_ASAP7_75t_L g727 ( .A(n_172), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_173), .A2(n_271), .B1(n_847), .B2(n_1166), .Y(n_1194) );
INVx1_ASAP7_75t_L g716 ( .A(n_175), .Y(n_716) );
INVx1_ASAP7_75t_L g933 ( .A(n_176), .Y(n_933) );
OAI211xp5_ASAP7_75t_L g1161 ( .A1(n_177), .A2(n_420), .B(n_725), .C(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1174 ( .A(n_177), .Y(n_1174) );
INVx1_ASAP7_75t_L g853 ( .A(n_178), .Y(n_853) );
AOI21xp33_ASAP7_75t_L g1041 ( .A1(n_180), .A2(n_549), .B(n_975), .Y(n_1041) );
INVx1_ASAP7_75t_L g904 ( .A(n_181), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g1038 ( .A(n_182), .Y(n_1038) );
INVx1_ASAP7_75t_L g906 ( .A(n_184), .Y(n_906) );
INVx1_ASAP7_75t_L g1504 ( .A(n_185), .Y(n_1504) );
OAI22xp33_ASAP7_75t_L g1578 ( .A1(n_187), .A2(n_270), .B1(n_296), .B2(n_1169), .Y(n_1578) );
INVx1_ASAP7_75t_L g835 ( .A(n_189), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_190), .A2(n_255), .B1(n_1276), .B2(n_1291), .Y(n_1313) );
INVx1_ASAP7_75t_L g711 ( .A(n_191), .Y(n_711) );
INVx1_ASAP7_75t_L g320 ( .A(n_192), .Y(n_320) );
INVx1_ASAP7_75t_L g753 ( .A(n_193), .Y(n_753) );
OAI211xp5_ASAP7_75t_SL g759 ( .A1(n_193), .A2(n_420), .B(n_760), .C(n_761), .Y(n_759) );
OAI222xp33_ASAP7_75t_L g1021 ( .A1(n_194), .A2(n_240), .B1(n_253), .B2(n_488), .C1(n_1022), .C2(n_1023), .Y(n_1021) );
XOR2x2_ASAP7_75t_L g309 ( .A(n_195), .B(n_310), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_196), .A2(n_279), .B1(n_554), .B2(n_576), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_196), .Y(n_1061) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_197), .A2(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g429 ( .A(n_199), .Y(n_429) );
INVx1_ASAP7_75t_L g930 ( .A(n_200), .Y(n_930) );
INVx1_ASAP7_75t_L g857 ( .A(n_201), .Y(n_857) );
INVx1_ASAP7_75t_L g808 ( .A(n_202), .Y(n_808) );
OAI211xp5_ASAP7_75t_L g814 ( .A1(n_202), .A2(n_635), .B(n_760), .C(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g1088 ( .A(n_203), .Y(n_1088) );
INVx1_ASAP7_75t_L g1132 ( .A(n_204), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_205), .A2(n_250), .B1(n_1276), .B2(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1570 ( .A(n_206), .Y(n_1570) );
OAI211xp5_ASAP7_75t_SL g1573 ( .A1(n_206), .A2(n_746), .B(n_838), .C(n_1574), .Y(n_1573) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
INVx1_ASAP7_75t_L g1084 ( .A(n_208), .Y(n_1084) );
INVx1_ASAP7_75t_L g1097 ( .A(n_209), .Y(n_1097) );
INVx1_ASAP7_75t_L g724 ( .A(n_210), .Y(n_724) );
INVx1_ASAP7_75t_L g790 ( .A(n_211), .Y(n_790) );
INVx1_ASAP7_75t_L g1553 ( .A(n_212), .Y(n_1553) );
INVx1_ASAP7_75t_L g626 ( .A(n_213), .Y(n_626) );
INVx1_ASAP7_75t_L g925 ( .A(n_214), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_215), .A2(n_231), .B1(n_545), .B2(n_547), .C(n_549), .Y(n_544) );
INVx1_ASAP7_75t_L g590 ( .A(n_215), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_218), .A2(n_241), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_218), .A2(n_241), .B1(n_847), .B2(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g623 ( .A(n_219), .Y(n_623) );
INVx1_ASAP7_75t_L g1136 ( .A(n_220), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_221), .Y(n_1027) );
XNOR2xp5_ASAP7_75t_L g1219 ( .A(n_222), .B(n_1220), .Y(n_1219) );
AO22x1_ASAP7_75t_L g1275 ( .A1(n_222), .A2(n_243), .B1(n_1276), .B2(n_1280), .Y(n_1275) );
CKINVDCx16_ASAP7_75t_R g1350 ( .A(n_224), .Y(n_1350) );
INVx1_ASAP7_75t_L g1198 ( .A(n_226), .Y(n_1198) );
INVx1_ASAP7_75t_L g343 ( .A(n_227), .Y(n_343) );
INVxp67_ASAP7_75t_SL g1005 ( .A(n_228), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g1249 ( .A1(n_229), .A2(n_276), .B1(n_1008), .B2(n_1250), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_231), .A2(n_278), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g1224 ( .A(n_232), .Y(n_1224) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_233), .A2(n_261), .B1(n_1283), .B2(n_1286), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_234), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_235), .A2(n_259), .B1(n_472), .B2(n_474), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_235), .A2(n_259), .B1(n_765), .B2(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g779 ( .A(n_236), .Y(n_779) );
BUFx3_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
INVx1_ASAP7_75t_L g449 ( .A(n_237), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_239), .Y(n_952) );
INVx1_ASAP7_75t_L g865 ( .A(n_246), .Y(n_865) );
INVx1_ASAP7_75t_L g1164 ( .A(n_247), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1172 ( .A1(n_247), .A2(n_746), .B(n_747), .C(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1096 ( .A(n_248), .Y(n_1096) );
INVx1_ASAP7_75t_L g641 ( .A(n_251), .Y(n_641) );
INVx2_ASAP7_75t_L g317 ( .A(n_252), .Y(n_317) );
INVx1_ASAP7_75t_L g363 ( .A(n_252), .Y(n_363) );
INVx1_ASAP7_75t_L g407 ( .A(n_252), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_253), .A2(n_262), .B1(n_664), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1489 ( .A(n_257), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1571 ( .A1(n_258), .A2(n_270), .B1(n_416), .B2(n_847), .Y(n_1571) );
AO22x1_ASAP7_75t_L g1282 ( .A1(n_260), .A2(n_274), .B1(n_1283), .B2(n_1286), .Y(n_1282) );
INVx1_ASAP7_75t_L g1028 ( .A(n_262), .Y(n_1028) );
INVx1_ASAP7_75t_L g1199 ( .A(n_264), .Y(n_1199) );
INVx1_ASAP7_75t_L g1230 ( .A(n_265), .Y(n_1230) );
XNOR2xp5_ASAP7_75t_L g700 ( .A(n_266), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g789 ( .A(n_267), .Y(n_789) );
INVx1_ASAP7_75t_L g1185 ( .A(n_268), .Y(n_1185) );
INVx1_ASAP7_75t_L g964 ( .A(n_269), .Y(n_964) );
INVx1_ASAP7_75t_L g1227 ( .A(n_273), .Y(n_1227) );
INVx1_ASAP7_75t_L g1546 ( .A(n_275), .Y(n_1546) );
XOR2x2_ASAP7_75t_L g1119 ( .A(n_277), .B(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1056 ( .A(n_279), .Y(n_1056) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_280), .B(n_770), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_305), .B(n_1268), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g1531 ( .A(n_284), .B(n_293), .Y(n_1531) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g1537 ( .A(n_286), .B(n_289), .Y(n_1537) );
INVx1_ASAP7_75t_L g1583 ( .A(n_286), .Y(n_1583) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_289), .B(n_1583), .Y(n_1585) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g478 ( .A(n_293), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g358 ( .A(n_294), .B(n_304), .Y(n_358) );
AND2x4_ASAP7_75t_L g550 ( .A(n_294), .B(n_303), .Y(n_550) );
INVx1_ASAP7_75t_L g916 ( .A(n_295), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_295), .A2(n_447), .B1(n_1227), .B2(n_1228), .Y(n_1226) );
AND2x4_ASAP7_75t_SL g1530 ( .A(n_295), .B(n_1531), .Y(n_1530) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_302), .Y(n_296) );
INVxp67_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
OR2x6_ASAP7_75t_L g473 ( .A(n_297), .B(n_448), .Y(n_473) );
INVx1_ASAP7_75t_L g1157 ( .A(n_297), .Y(n_1157) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
BUFx4f_ASAP7_75t_L g733 ( .A(n_298), .Y(n_733) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
INVx2_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
NAND2x1_ASAP7_75t_L g339 ( .A(n_300), .B(n_301), .Y(n_339) );
AND2x2_ASAP7_75t_L g450 ( .A(n_300), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g460 ( .A(n_300), .B(n_301), .Y(n_460) );
INVx1_ASAP7_75t_L g469 ( .A(n_300), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_301), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g334 ( .A(n_301), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g451 ( .A(n_301), .Y(n_451) );
BUFx2_ASAP7_75t_L g464 ( .A(n_301), .Y(n_464) );
INVx1_ASAP7_75t_L g504 ( .A(n_301), .Y(n_504) );
AND2x2_ASAP7_75t_L g555 ( .A(n_301), .B(n_328), .Y(n_555) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g457 ( .A(n_303), .Y(n_457) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g463 ( .A(n_304), .Y(n_463) );
AND2x4_ASAP7_75t_L g467 ( .A(n_304), .B(n_468), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_1116), .B1(n_1117), .B2(n_1267), .Y(n_305) );
INVx1_ASAP7_75t_L g1267 ( .A(n_306), .Y(n_1267) );
XNOR2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_895), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_698), .B1(n_893), .B2(n_894), .Y(n_307) );
INVx1_ASAP7_75t_L g894 ( .A(n_308), .Y(n_894) );
AO22x2_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_481), .B1(n_482), .B2(n_697), .Y(n_308) );
INVx1_ASAP7_75t_L g697 ( .A(n_309), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_413), .C(n_444), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_364), .Y(n_311) );
OAI33xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .A3(n_329), .B1(n_340), .B2(n_348), .B3(n_356), .Y(n_312) );
OAI33xp33_ASAP7_75t_L g728 ( .A1(n_313), .A2(n_729), .A3(n_735), .B1(n_739), .B2(n_741), .B3(n_742), .Y(n_728) );
OAI33xp33_ASAP7_75t_L g792 ( .A1(n_313), .A2(n_741), .A3(n_793), .B1(n_797), .B2(n_798), .B3(n_800), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_313), .A2(n_356), .B1(n_936), .B2(n_943), .Y(n_935) );
INVx1_ASAP7_75t_L g1253 ( .A(n_313), .Y(n_1253) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g851 ( .A(n_315), .Y(n_851) );
INVx1_ASAP7_75t_L g1099 ( .A(n_315), .Y(n_1099) );
INVx2_ASAP7_75t_L g1142 ( .A(n_315), .Y(n_1142) );
INVx4_ASAP7_75t_L g1544 ( .A(n_315), .Y(n_1544) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g586 ( .A(n_316), .Y(n_586) );
OR2x6_ASAP7_75t_L g1501 ( .A(n_316), .B(n_1502), .Y(n_1501) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g695 ( .A(n_317), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B1(n_323), .B2(n_324), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_320), .A2(n_343), .B1(n_371), .B2(n_378), .Y(n_370) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_323), .A2(n_347), .B1(n_371), .B2(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g1146 ( .A(n_324), .Y(n_1146) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
INVx1_ASAP7_75t_L g796 ( .A(n_325), .Y(n_796) );
INVx4_ASAP7_75t_L g860 ( .A(n_325), .Y(n_860) );
INVx1_ASAP7_75t_L g1210 ( .A(n_325), .Y(n_1210) );
INVx8_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g476 ( .A(n_326), .B(n_463), .Y(n_476) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_336), .B2(n_337), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_330), .A2(n_352), .B1(n_386), .B2(n_392), .Y(n_385) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g799 ( .A(n_332), .Y(n_799) );
INVx2_ASAP7_75t_L g1148 ( .A(n_332), .Y(n_1148) );
INVx4_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g342 ( .A(n_334), .Y(n_342) );
INVx2_ASAP7_75t_L g738 ( .A(n_334), .Y(n_738) );
BUFx3_ASAP7_75t_L g1152 ( .A(n_334), .Y(n_1152) );
AND2x2_ASAP7_75t_L g503 ( .A(n_335), .B(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_335), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_336), .A2(n_353), .B1(n_397), .B2(n_400), .Y(n_396) );
BUFx4f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx4_ASAP7_75t_L g454 ( .A(n_338), .Y(n_454) );
BUFx4f_ASAP7_75t_L g864 ( .A(n_338), .Y(n_864) );
BUFx4f_ASAP7_75t_L g938 ( .A(n_338), .Y(n_938) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g346 ( .A(n_339), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_344), .B2(n_347), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI211xp5_ASAP7_75t_L g570 ( .A1(n_344), .A2(n_571), .B(n_572), .C(n_575), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_344), .A2(n_711), .B1(n_716), .B2(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_344), .A2(n_736), .B1(n_779), .B2(n_784), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_344), .A2(n_862), .B1(n_867), .B2(n_868), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1551 ( .A1(n_344), .A2(n_1150), .B1(n_1552), .B2(n_1553), .Y(n_1551) );
INVx5_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g670 ( .A(n_346), .Y(n_670) );
BUFx2_ASAP7_75t_SL g740 ( .A(n_346), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B1(n_353), .B2(n_354), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g971 ( .A1(n_349), .A2(n_858), .B1(n_972), .B2(n_973), .C(n_974), .Y(n_971) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g856 ( .A(n_351), .Y(n_856) );
INVx5_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx6_ASAP7_75t_L g734 ( .A(n_355), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g741 ( .A(n_357), .Y(n_741) );
AOI33xp33_ASAP7_75t_L g1252 ( .A1(n_357), .A2(n_1253), .A3(n_1254), .B1(n_1258), .B2(n_1262), .B3(n_1265), .Y(n_1252) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx4_ASAP7_75t_L g574 ( .A(n_358), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_358), .B(n_359), .Y(n_871) );
INVx1_ASAP7_75t_SL g960 ( .A(n_358), .Y(n_960) );
INVx4_ASAP7_75t_L g1515 ( .A(n_358), .Y(n_1515) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g366 ( .A(n_361), .B(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_361), .Y(n_443) );
OR2x2_ASAP7_75t_L g510 ( .A(n_361), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g480 ( .A(n_362), .Y(n_480) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI33xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_370), .A3(n_385), .B1(n_396), .B2(n_404), .B3(n_409), .Y(n_364) );
OAI33xp33_ASAP7_75t_L g772 ( .A1(n_365), .A2(n_720), .A3(n_773), .B1(n_778), .B2(n_783), .B3(n_788), .Y(n_772) );
BUFx8_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_366), .Y(n_597) );
BUFx4f_ASAP7_75t_L g647 ( .A(n_366), .Y(n_647) );
BUFx2_ASAP7_75t_L g995 ( .A(n_366), .Y(n_995) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_369), .Y(n_367) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_368), .Y(n_441) );
INVx1_ASAP7_75t_L g493 ( .A(n_368), .Y(n_493) );
AND3x4_ASAP7_75t_L g1065 ( .A(n_368), .B(n_427), .C(n_695), .Y(n_1065) );
INVx3_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
BUFx3_ASAP7_75t_L g427 ( .A(n_369), .Y(n_427) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x4_ASAP7_75t_L g415 ( .A(n_374), .B(n_405), .Y(n_415) );
OR2x4_ASAP7_75t_L g435 ( .A(n_374), .B(n_418), .Y(n_435) );
INVx2_ASAP7_75t_L g507 ( .A(n_374), .Y(n_507) );
BUFx3_ASAP7_75t_L g706 ( .A(n_374), .Y(n_706) );
BUFx4f_ASAP7_75t_L g879 ( .A(n_374), .Y(n_879) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_375), .Y(n_384) );
INVx2_ASAP7_75t_L g391 ( .A(n_375), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_375), .B(n_383), .Y(n_395) );
AND2x4_ASAP7_75t_L g422 ( .A(n_375), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g491 ( .A(n_376), .Y(n_491) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g390 ( .A(n_377), .Y(n_390) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_SL g1567 ( .A(n_379), .Y(n_1567) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
BUFx3_ASAP7_75t_L g777 ( .A(n_381), .Y(n_777) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
BUFx2_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
BUFx2_ASAP7_75t_L g428 ( .A(n_384), .Y(n_428) );
INVx2_ASAP7_75t_L g527 ( .A(n_384), .Y(n_527) );
AND2x4_ASAP7_75t_L g605 ( .A(n_384), .B(n_533), .Y(n_605) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g515 ( .A(n_387), .B(n_509), .Y(n_515) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g603 ( .A(n_388), .Y(n_603) );
BUFx2_ASAP7_75t_L g649 ( .A(n_388), .Y(n_649) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_389), .Y(n_399) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_389), .Y(n_713) );
BUFx8_ASAP7_75t_L g988 ( .A(n_389), .Y(n_988) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x4_ASAP7_75t_L g490 ( .A(n_391), .B(n_491), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_392), .A2(n_639), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_392), .A2(n_711), .B1(n_712), .B2(n_714), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_392), .A2(n_779), .B1(n_780), .B2(n_782), .Y(n_778) );
CKINVDCx8_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g651 ( .A(n_393), .Y(n_651) );
INVx3_ASAP7_75t_L g719 ( .A(n_393), .Y(n_719) );
INVx3_ASAP7_75t_L g883 ( .A(n_393), .Y(n_883) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g538 ( .A(n_394), .Y(n_538) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g403 ( .A(n_395), .Y(n_403) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g417 ( .A(n_399), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g589 ( .A(n_399), .Y(n_589) );
INVx1_ASAP7_75t_L g717 ( .A(n_399), .Y(n_717) );
INVx2_ASAP7_75t_L g926 ( .A(n_399), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_400), .A2(n_589), .B1(n_590), .B2(n_591), .C(n_592), .Y(n_588) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g1133 ( .A(n_402), .Y(n_1133) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x6_ASAP7_75t_L g438 ( .A(n_403), .B(n_405), .Y(n_438) );
BUFx3_ASAP7_75t_L g787 ( .A(n_403), .Y(n_787) );
INVx3_ASAP7_75t_L g611 ( .A(n_404), .Y(n_611) );
INVx3_ASAP7_75t_L g1003 ( .A(n_404), .Y(n_1003) );
NAND3x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .C(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g418 ( .A(n_405), .Y(n_418) );
AND2x4_ASAP7_75t_L g421 ( .A(n_405), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g492 ( .A(n_405), .B(n_493), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g1502 ( .A(n_405), .B(n_408), .Y(n_1502) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g525 ( .A(n_407), .Y(n_525) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g760 ( .A(n_411), .Y(n_760) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g541 ( .A(n_412), .B(n_510), .Y(n_541) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_412), .Y(n_709) );
INVx3_ASAP7_75t_L g726 ( .A(n_412), .Y(n_726) );
OAI31xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_419), .A3(n_433), .B(n_439), .Y(n_413) );
INVx2_ASAP7_75t_SL g632 ( .A(n_415), .Y(n_632) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_415), .Y(n_757) );
INVx1_ASAP7_75t_L g951 ( .A(n_415), .Y(n_951) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_415), .Y(n_1107) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_417), .A2(n_619), .B1(n_620), .B2(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g758 ( .A(n_417), .Y(n_758) );
INVx1_ASAP7_75t_L g813 ( .A(n_417), .Y(n_813) );
INVx2_ASAP7_75t_L g1108 ( .A(n_417), .Y(n_1108) );
INVx1_ASAP7_75t_L g1166 ( .A(n_417), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_417), .A2(n_632), .B1(n_1227), .B2(n_1228), .Y(n_1241) );
CKINVDCx8_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
CKINVDCx8_ASAP7_75t_R g635 ( .A(n_421), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g1235 ( .A1(n_421), .A2(n_645), .B(n_1233), .C(n_1236), .Y(n_1235) );
BUFx2_ASAP7_75t_L g596 ( .A(n_422), .Y(n_596) );
BUFx2_ASAP7_75t_L g600 ( .A(n_422), .Y(n_600) );
INVx2_ASAP7_75t_L g610 ( .A(n_422), .Y(n_610) );
BUFx2_ASAP7_75t_L g629 ( .A(n_422), .Y(n_629) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_422), .Y(n_1000) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_422), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_422), .Y(n_1251) );
INVx1_ASAP7_75t_L g533 ( .A(n_423), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_429), .B1(n_430), .B2(n_432), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_425), .A2(n_430), .B1(n_1163), .B2(n_1164), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_425), .A2(n_430), .B1(n_1185), .B2(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1237 ( .A(n_425), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1568 ( .A1(n_425), .A2(n_430), .B1(n_1569), .B2(n_1570), .Y(n_1568) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
AND2x4_ASAP7_75t_L g430 ( .A(n_426), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g625 ( .A(n_426), .B(n_428), .Y(n_625) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_429), .A2(n_462), .B1(n_465), .B2(n_470), .Y(n_461) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_430), .Y(n_627) );
INVx1_ASAP7_75t_L g1238 ( .A(n_430), .Y(n_1238) );
INVx1_ASAP7_75t_L g1240 ( .A(n_434), .Y(n_1240) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g634 ( .A(n_435), .Y(n_634) );
BUFx2_ASAP7_75t_L g765 ( .A(n_435), .Y(n_765) );
BUFx2_ASAP7_75t_L g846 ( .A(n_435), .Y(n_846) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g621 ( .A(n_438), .Y(n_621) );
INVx1_ASAP7_75t_L g767 ( .A(n_438), .Y(n_767) );
BUFx3_ASAP7_75t_L g847 ( .A(n_438), .Y(n_847) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_442), .Y(n_439) );
AND2x4_ASAP7_75t_L g636 ( .A(n_440), .B(n_442), .Y(n_636) );
AND2x2_ASAP7_75t_SL g768 ( .A(n_440), .B(n_442), .Y(n_768) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_452), .A3(n_471), .B(n_477), .Y(n_444) );
INVx4_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_SL g830 ( .A(n_447), .Y(n_830) );
CKINVDCx16_ASAP7_75t_R g1169 ( .A(n_447), .Y(n_1169) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_450), .Y(n_519) );
INVx2_ASAP7_75t_L g673 ( .A(n_450), .Y(n_673) );
BUFx3_ASAP7_75t_L g975 ( .A(n_450), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g1035 ( .A(n_453), .B(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g832 ( .A(n_454), .Y(n_832) );
INVx2_ASAP7_75t_L g1045 ( .A(n_454), .Y(n_1045) );
INVx2_ASAP7_75t_L g1205 ( .A(n_454), .Y(n_1205) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AND2x2_ASAP7_75t_L g748 ( .A(n_457), .B(n_548), .Y(n_748) );
INVx1_ASAP7_75t_L g1264 ( .A(n_458), .Y(n_1264) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g566 ( .A(n_459), .Y(n_566) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_460), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_462), .A2(n_750), .B1(n_751), .B2(n_753), .Y(n_749) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AND2x4_ASAP7_75t_L g806 ( .A(n_463), .B(n_464), .Y(n_806) );
AND2x2_ASAP7_75t_L g905 ( .A(n_463), .B(n_675), .Y(n_905) );
INVx1_ASAP7_75t_L g563 ( .A(n_464), .Y(n_563) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_464), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_465), .A2(n_834), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g752 ( .A(n_467), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_467), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
BUFx3_ASAP7_75t_L g836 ( .A(n_467), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_468), .B(n_569), .Y(n_690) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g824 ( .A(n_473), .Y(n_824) );
HB1xp67_ASAP7_75t_L g1077 ( .A(n_473), .Y(n_1077) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g1078 ( .A(n_475), .Y(n_1078) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g828 ( .A(n_476), .Y(n_828) );
BUFx2_ASAP7_75t_L g908 ( .A(n_476), .Y(n_908) );
OAI31xp33_ASAP7_75t_L g743 ( .A1(n_477), .A2(n_744), .A3(n_745), .B(n_754), .Y(n_743) );
OAI31xp33_ASAP7_75t_L g1182 ( .A1(n_477), .A2(n_1183), .A3(n_1187), .B(n_1188), .Y(n_1182) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_SL g810 ( .A(n_478), .Y(n_810) );
INVx1_ASAP7_75t_L g820 ( .A(n_478), .Y(n_820) );
BUFx2_ASAP7_75t_L g917 ( .A(n_478), .Y(n_917) );
OAI31xp33_ASAP7_75t_L g1070 ( .A1(n_478), .A2(n_1071), .A3(n_1075), .B(n_1076), .Y(n_1070) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_478), .A2(n_636), .B1(n_1222), .B2(n_1234), .Y(n_1221) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g494 ( .A(n_480), .Y(n_494) );
INVx1_ASAP7_75t_L g500 ( .A(n_480), .Y(n_500) );
OR2x2_ASAP7_75t_L g983 ( .A(n_480), .B(n_690), .Y(n_983) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
XOR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_614), .Y(n_482) );
INVx1_ASAP7_75t_L g612 ( .A(n_484), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .C(n_520), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_486), .A2(n_579), .B1(n_582), .B2(n_583), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g1488 ( .A1(n_487), .A2(n_1012), .B1(n_1489), .B2(n_1490), .C(n_1491), .Y(n_1488) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
BUFx3_ASAP7_75t_L g595 ( .A(n_490), .Y(n_595) );
INVx8_ASAP7_75t_L g608 ( .A(n_490), .Y(n_608) );
BUFx3_ASAP7_75t_L g644 ( .A(n_490), .Y(n_644) );
HB1xp67_ASAP7_75t_L g1495 ( .A(n_490), .Y(n_1495) );
AND2x4_ASAP7_75t_L g524 ( .A(n_492), .B(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_512), .B2(n_513), .Y(n_495) );
INVxp67_ASAP7_75t_L g1022 ( .A(n_497), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AND2x4_ASAP7_75t_L g517 ( .A(n_500), .B(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_501), .Y(n_663) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x2_ASAP7_75t_L g518 ( .A(n_502), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g579 ( .A(n_502), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_SL g584 ( .A(n_502), .B(n_548), .Y(n_584) );
AND2x4_ASAP7_75t_L g667 ( .A(n_502), .B(n_519), .Y(n_667) );
AND2x4_ASAP7_75t_L g957 ( .A(n_502), .B(n_676), .Y(n_957) );
INVx3_ASAP7_75t_L g553 ( .A(n_503), .Y(n_553) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_503), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_503), .B(n_569), .Y(n_684) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx2_ASAP7_75t_SL g889 ( .A(n_506), .Y(n_889) );
OAI22xp33_ASAP7_75t_L g1213 ( .A1(n_506), .A2(n_880), .B1(n_1198), .B2(n_1204), .Y(n_1213) );
OAI22xp33_ASAP7_75t_L g1558 ( .A1(n_506), .A2(n_890), .B1(n_1546), .B2(n_1552), .Y(n_1558) );
OAI22xp33_ASAP7_75t_L g1562 ( .A1(n_506), .A2(n_725), .B1(n_1547), .B2(n_1553), .Y(n_1562) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g723 ( .A(n_507), .Y(n_723) );
INVxp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g537 ( .A(n_510), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g987 ( .A(n_510), .Y(n_987) );
INVx1_ASAP7_75t_L g1023 ( .A(n_513), .Y(n_1023) );
NAND2x1_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_515), .A2(n_1519), .B1(n_1520), .B2(n_1525), .Y(n_1524) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_519), .Y(n_573) );
NOR3xp33_ASAP7_75t_SL g520 ( .A(n_521), .B(n_542), .C(n_587), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_SL g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AND2x4_ASAP7_75t_SL g529 ( .A(n_524), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g599 ( .A(n_524), .B(n_600), .Y(n_599) );
NAND2x1_ASAP7_75t_L g991 ( .A(n_524), .B(n_526), .Y(n_991) );
AND2x4_ASAP7_75t_L g993 ( .A(n_524), .B(n_530), .Y(n_993) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_524), .B(n_526), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_525), .B(n_684), .Y(n_1014) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_539), .B2(n_540), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_535), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_537), .B(n_1014), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_539), .A2(n_560), .B1(n_562), .B2(n_564), .C(n_565), .Y(n_559) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g982 ( .A(n_541), .B(n_983), .Y(n_982) );
AND2x4_ASAP7_75t_L g1523 ( .A(n_541), .B(n_983), .Y(n_1523) );
AOI31xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_570), .A3(n_578), .B(n_585), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_551), .B(n_556), .Y(n_543) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x6_ASAP7_75t_L g691 ( .A(n_548), .B(n_569), .Y(n_691) );
BUFx3_ASAP7_75t_L g911 ( .A(n_548), .Y(n_911) );
BUFx3_ASAP7_75t_L g976 ( .A(n_548), .Y(n_976) );
BUFx3_ASAP7_75t_L g1231 ( .A(n_548), .Y(n_1231) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g680 ( .A(n_550), .Y(n_680) );
INVx1_ASAP7_75t_L g977 ( .A(n_550), .Y(n_977) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g558 ( .A(n_553), .Y(n_558) );
INVx1_ASAP7_75t_L g576 ( .A(n_553), .Y(n_576) );
INVx1_ASAP7_75t_L g1255 ( .A(n_553), .Y(n_1255) );
INVx1_ASAP7_75t_SL g1257 ( .A(n_554), .Y(n_1257) );
BUFx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx3_ASAP7_75t_L g577 ( .A(n_555), .Y(n_577) );
INVx2_ASAP7_75t_L g581 ( .A(n_555), .Y(n_581) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_555), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B(n_567), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_560), .A2(n_1027), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_563), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g1261 ( .A(n_565), .Y(n_1261) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_568), .A2(n_1033), .B(n_1034), .C(n_1035), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g687 ( .A(n_569), .Y(n_687) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_569), .B(n_1037), .Y(n_1512) );
BUFx3_ASAP7_75t_L g1259 ( .A(n_573), .Y(n_1259) );
INVx2_ASAP7_75t_L g664 ( .A(n_579), .Y(n_664) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI211xp5_ASAP7_75t_SL g682 ( .A1(n_583), .A2(n_626), .B(n_683), .C(n_691), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g1509 ( .A1(n_583), .A2(n_1504), .B1(n_1506), .B2(n_1510), .C1(n_1511), .C2(n_1512), .Y(n_1509) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g969 ( .A(n_584), .Y(n_969) );
INVx1_ASAP7_75t_L g978 ( .A(n_585), .Y(n_978) );
BUFx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI211xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_597), .B(n_598), .C(n_601), .Y(n_587) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g998 ( .A(n_595), .Y(n_998) );
OAI33xp33_ASAP7_75t_L g703 ( .A1(n_597), .A2(n_704), .A3(n_710), .B1(n_715), .B2(n_720), .B3(n_721), .Y(n_703) );
OAI33xp33_ASAP7_75t_L g875 ( .A1(n_597), .A2(n_658), .A3(n_876), .B1(n_882), .B2(n_884), .B3(n_887), .Y(n_875) );
OAI33xp33_ASAP7_75t_L g1212 ( .A1(n_597), .A2(n_658), .A3(n_1213), .B1(n_1214), .B2(n_1216), .B3(n_1217), .Y(n_1212) );
OAI33xp33_ASAP7_75t_L g1557 ( .A1(n_597), .A2(n_1558), .A3(n_1559), .B1(n_1560), .B2(n_1561), .B3(n_1562), .Y(n_1557) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_599), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_599), .A2(n_611), .B1(n_1052), .B2(n_1057), .C(n_1064), .Y(n_1051) );
INVx3_ASAP7_75t_L g1492 ( .A(n_599), .Y(n_1492) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_606), .C(n_611), .Y(n_601) );
INVx1_ASAP7_75t_L g639 ( .A(n_603), .Y(n_639) );
INVx1_ASAP7_75t_L g785 ( .A(n_603), .Y(n_785) );
BUFx12f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_605), .Y(n_1054) );
INVx5_ASAP7_75t_L g1246 ( .A(n_605), .Y(n_1246) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx8_ASAP7_75t_L g1008 ( .A(n_608), .Y(n_1008) );
INVx2_ASAP7_75t_L g1526 ( .A(n_608), .Y(n_1526) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g645 ( .A(n_610), .Y(n_645) );
INVx2_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_611), .Y(n_720) );
INVx2_ASAP7_75t_L g1561 ( .A(n_611), .Y(n_1561) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_636), .B(n_637), .C(n_659), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .C(n_630), .D(n_635), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_621), .A2(n_634), .B1(n_904), .B2(n_906), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_621), .A2(n_1224), .B1(n_1225), .B2(n_1240), .Y(n_1239) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_626), .B2(n_627), .C1(n_628), .C2(n_629), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_624), .A2(n_627), .B1(n_807), .B2(n_816), .Y(n_815) );
AOI222xp33_ASAP7_75t_L g947 ( .A1(n_624), .A2(n_627), .B1(n_656), .B2(n_910), .C1(n_912), .C2(n_913), .Y(n_947) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx3_ASAP7_75t_L g762 ( .A(n_625), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_627), .A2(n_750), .B1(n_762), .B2(n_763), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_627), .A2(n_762), .B1(n_835), .B2(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_627), .A2(n_762), .B1(n_1073), .B2(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_628), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g657 ( .A(n_629), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
INVx2_ASAP7_75t_L g841 ( .A(n_632), .Y(n_841) );
INVx1_ASAP7_75t_L g1113 ( .A(n_634), .Y(n_1113) );
INVx2_ASAP7_75t_L g1160 ( .A(n_634), .Y(n_1160) );
NAND3xp33_ASAP7_75t_L g946 ( .A(n_635), .B(n_947), .C(n_948), .Y(n_946) );
CKINVDCx14_ASAP7_75t_R g848 ( .A(n_636), .Y(n_848) );
OAI31xp33_ASAP7_75t_L g1563 ( .A1(n_636), .A2(n_1564), .A3(n_1565), .B(n_1571), .Y(n_1563) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_646), .B1(n_648), .B2(n_658), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_639), .A2(n_863), .B1(n_873), .B2(n_883), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_639), .A2(n_1085), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g655 ( .A(n_644), .Y(n_655) );
OAI33xp33_ASAP7_75t_L g919 ( .A1(n_646), .A2(n_720), .A3(n_920), .B1(n_924), .B2(n_928), .B3(n_932), .Y(n_919) );
OAI33xp33_ASAP7_75t_L g1080 ( .A1(n_646), .A2(n_1001), .A3(n_1081), .B1(n_1087), .B2(n_1091), .B3(n_1095), .Y(n_1080) );
OAI33xp33_ASAP7_75t_L g1122 ( .A1(n_646), .A2(n_658), .A3(n_1123), .B1(n_1127), .B2(n_1134), .B3(n_1137), .Y(n_1122) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_651), .B2(n_652), .C(n_653), .Y(n_648) );
OAI211xp5_ASAP7_75t_SL g677 ( .A1(n_650), .A2(n_670), .B(n_678), .C(n_681), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_651), .A2(n_865), .B1(n_874), .B2(n_885), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_651), .A2(n_1092), .B1(n_1202), .B2(n_1211), .Y(n_1216) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_682), .B(n_692), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_663), .A2(n_667), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_663), .A2(n_667), .B1(n_1519), .B2(n_1520), .Y(n_1518) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_671), .C(n_674), .Y(n_668) );
BUFx2_ASAP7_75t_L g746 ( .A(n_670), .Y(n_746) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g679 ( .A(n_673), .Y(n_679) );
INVx3_ASAP7_75t_L g941 ( .A(n_675), .Y(n_941) );
BUFx6f_ASAP7_75t_L g1034 ( .A(n_675), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_676), .Y(n_942) );
BUFx2_ASAP7_75t_L g962 ( .A(n_676), .Y(n_962) );
BUFx2_ASAP7_75t_L g970 ( .A(n_685), .Y(n_970) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_691), .A2(n_959), .B(n_961), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_691), .A2(n_957), .B1(n_1489), .B2(n_1514), .C(n_1516), .Y(n_1513) );
INVx1_ASAP7_75t_L g1521 ( .A(n_692), .Y(n_1521) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_693), .Y(n_1050) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g893 ( .A(n_698), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_818), .B1(n_891), .B2(n_892), .Y(n_698) );
INVx1_ASAP7_75t_L g891 ( .A(n_699), .Y(n_891) );
XOR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_769), .Y(n_699) );
AND3x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_743), .C(n_755), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_728), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_705), .A2(n_724), .B1(n_730), .B2(n_734), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_706), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_706), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
OAI22xp33_ASAP7_75t_L g920 ( .A1(n_706), .A2(n_921), .B1(n_922), .B2(n_923), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_706), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_707), .A2(n_727), .B1(n_736), .B2(n_740), .Y(n_739) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_709), .Y(n_931) );
INVx1_ASAP7_75t_L g1086 ( .A(n_709), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1559 ( .A1(n_712), .A2(n_787), .B1(n_1549), .B2(n_1555), .Y(n_1559) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx5_ASAP7_75t_L g781 ( .A(n_713), .Y(n_781) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_713), .Y(n_886) );
INVx3_ASAP7_75t_L g1131 ( .A(n_713), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_714), .A2(n_718), .B1(n_732), .B2(n_734), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_717), .A2(n_719), .B1(n_933), .B2(n_934), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_719), .A2(n_1138), .B1(n_1139), .B2(n_1140), .Y(n_1137) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_724), .B1(n_725), .B2(n_727), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_722), .A2(n_760), .B1(n_1044), .B2(n_1056), .Y(n_1055) );
BUFx4f_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g1063 ( .A(n_726), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_730), .A2(n_858), .B1(n_1082), .B2(n_1096), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_730), .A2(n_858), .B1(n_1090), .B2(n_1094), .Y(n_1103) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_733), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_734), .A2(n_782), .B1(n_786), .B2(n_801), .Y(n_800) );
INVx4_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g862 ( .A(n_738), .Y(n_862) );
INVx2_ASAP7_75t_L g937 ( .A(n_738), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_740), .A2(n_775), .B1(n_790), .B2(n_799), .Y(n_798) );
OAI33xp33_ASAP7_75t_L g1141 ( .A1(n_741), .A2(n_1142), .A3(n_1143), .B1(n_1147), .B2(n_1149), .B3(n_1153), .Y(n_1141) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx3_ASAP7_75t_L g838 ( .A(n_748), .Y(n_838) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g914 ( .A(n_752), .Y(n_914) );
OAI31xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .A3(n_764), .B(n_768), .Y(n_755) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI31xp33_ASAP7_75t_L g811 ( .A1(n_768), .A2(n_812), .A3(n_814), .B(n_817), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g945 ( .A1(n_768), .A2(n_946), .B(n_949), .Y(n_945) );
OAI31xp33_ASAP7_75t_L g1104 ( .A1(n_768), .A2(n_1105), .A3(n_1109), .B(n_1112), .Y(n_1104) );
OAI31xp33_ASAP7_75t_SL g1158 ( .A1(n_768), .A2(n_1159), .A3(n_1161), .B(n_1165), .Y(n_1158) );
OAI31xp33_ASAP7_75t_SL g1189 ( .A1(n_768), .A2(n_1190), .A3(n_1191), .B(n_1194), .Y(n_1189) );
AND3x1_ASAP7_75t_L g770 ( .A(n_771), .B(n_802), .C(n_811), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_792), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_774), .A2(n_789), .B1(n_794), .B2(n_796), .Y(n_793) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_777), .Y(n_791) );
INVx2_ASAP7_75t_L g881 ( .A(n_777), .Y(n_881) );
BUFx6f_ASAP7_75t_L g890 ( .A(n_777), .Y(n_890) );
BUFx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx8_ASAP7_75t_L g1053 ( .A(n_781), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_786), .B2(n_787), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g1004 ( .A1(n_785), .A2(n_883), .B1(n_1005), .B2(n_1006), .C(n_1007), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_787), .A2(n_925), .B1(n_926), .B2(n_927), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_787), .A2(n_1201), .B1(n_1208), .B2(n_1215), .Y(n_1214) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g801 ( .A(n_795), .Y(n_801) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_795), .Y(n_1144) );
OAI31xp33_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_804), .A3(n_809), .B(n_810), .Y(n_802) );
BUFx3_ASAP7_75t_L g834 ( .A(n_806), .Y(n_834) );
AOI222xp33_ASAP7_75t_L g1229 ( .A1(n_806), .A2(n_914), .B1(n_1230), .B2(n_1231), .C1(n_1232), .C2(n_1233), .Y(n_1229) );
OAI31xp33_ASAP7_75t_L g1167 ( .A1(n_810), .A2(n_1168), .A3(n_1170), .B(n_1172), .Y(n_1167) );
OAI31xp33_ASAP7_75t_L g1572 ( .A1(n_810), .A2(n_1573), .A3(n_1576), .B(n_1578), .Y(n_1572) );
INVx1_ASAP7_75t_L g892 ( .A(n_818), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_821), .B1(n_839), .B2(n_848), .C(n_849), .Y(n_819) );
NOR3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_829), .C(n_831), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_828), .A2(n_905), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_832), .A2(n_1040), .B(n_1041), .C(n_1042), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g1153 ( .A1(n_832), .A2(n_1132), .B1(n_1136), .B2(n_1154), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_833) );
AOI222xp33_ASAP7_75t_L g909 ( .A1(n_834), .A2(n_910), .B1(n_911), .B2(n_912), .C1(n_913), .C2(n_914), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_834), .A2(n_836), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_834), .A2(n_836), .B1(n_1163), .B2(n_1174), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_834), .A2(n_836), .B1(n_1569), .B2(n_1575), .Y(n_1574) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_838), .B(n_903), .C(n_909), .Y(n_902) );
NAND4xp25_ASAP7_75t_L g1222 ( .A(n_838), .B(n_1223), .C(n_1226), .D(n_1229), .Y(n_1222) );
NOR3xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_842), .C(n_845), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_875), .Y(n_849) );
OAI33xp33_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .A3(n_861), .B1(n_866), .B2(n_869), .B3(n_872), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_854), .B1(n_857), .B2(n_858), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_853), .A2(n_867), .B1(n_877), .B2(n_880), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_854), .A2(n_858), .B1(n_873), .B2(n_874), .Y(n_872) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g887 ( .A1(n_857), .A2(n_868), .B1(n_888), .B2(n_890), .Y(n_887) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_862), .A2(n_864), .B1(n_1088), .B2(n_1093), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_862), .A2(n_864), .B1(n_1084), .B2(n_1097), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_864), .A2(n_1148), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
OAI33xp33_ASAP7_75t_L g1098 ( .A1(n_869), .A2(n_1099), .A3(n_1100), .B1(n_1101), .B2(n_1102), .B3(n_1103), .Y(n_1098) );
OAI33xp33_ASAP7_75t_L g1196 ( .A1(n_869), .A2(n_1099), .A3(n_1197), .B1(n_1200), .B2(n_1203), .B3(n_1207), .Y(n_1196) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
OAI33xp33_ASAP7_75t_L g1543 ( .A1(n_871), .A2(n_1544), .A3(n_1545), .B1(n_1548), .B2(n_1551), .B3(n_1554), .Y(n_1543) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_879), .A2(n_1061), .B1(n_1062), .B2(n_1063), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_879), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_879), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_880), .A2(n_1083), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g923 ( .A(n_881), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_883), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_883), .A2(n_1092), .B1(n_1093), .B2(n_1094), .Y(n_1091) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g1083 ( .A(n_889), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g1123 ( .A1(n_890), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1123) );
OAI22xp33_ASAP7_75t_L g1217 ( .A1(n_890), .A2(n_1125), .B1(n_1199), .B2(n_1206), .Y(n_1217) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
OA22x2_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_898), .B1(n_1016), .B2(n_1017), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
XNOR2x1_ASAP7_75t_L g898 ( .A(n_899), .B(n_953), .Y(n_898) );
XOR2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_952), .Y(n_899) );
NAND3x1_ASAP7_75t_L g900 ( .A(n_901), .B(n_918), .C(n_945), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_915), .B(n_917), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_905), .B1(n_906), .B2(n_907), .Y(n_903) );
INVx1_ASAP7_75t_L g1171 ( .A(n_907), .Y(n_1171) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
HB1xp67_ASAP7_75t_L g1577 ( .A(n_908), .Y(n_1577) );
NOR2x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_935), .Y(n_918) );
OAI221xp5_ASAP7_75t_SL g943 ( .A1(n_922), .A2(n_930), .B1(n_937), .B2(n_938), .C(n_944), .Y(n_943) );
OAI221xp5_ASAP7_75t_SL g936 ( .A1(n_925), .A2(n_933), .B1(n_937), .B2(n_938), .C(n_939), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_938), .A2(n_1128), .B1(n_1135), .B2(n_1148), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1548 ( .A1(n_938), .A2(n_1148), .B1(n_1549), .B2(n_1550), .Y(n_1548) );
INVx2_ASAP7_75t_SL g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g1517 ( .A(n_941), .Y(n_1517) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OAI22xp5_ASAP7_75t_SL g1349 ( .A1(n_952), .A2(n_1350), .B1(n_1351), .B2(n_1352), .Y(n_1349) );
O2A1O1Ixp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_966), .B(n_978), .C(n_979), .Y(n_954) );
INVx3_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g1049 ( .A(n_968), .Y(n_1049) );
INVx4_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
OAI21xp5_ASAP7_75t_L g996 ( .A1(n_972), .A2(n_997), .B(n_999), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_989), .C(n_1010), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_981), .B(n_984), .Y(n_980) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
AND2x4_ASAP7_75t_L g1525 ( .A(n_987), .B(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_988), .Y(n_1059) );
INVx3_ASAP7_75t_L g1092 ( .A(n_988), .Y(n_1092) );
INVx3_ASAP7_75t_L g1215 ( .A(n_988), .Y(n_1215) );
NOR2xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_994), .Y(n_989) );
INVx2_ASAP7_75t_L g1026 ( .A(n_991), .Y(n_1026) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_993), .A2(n_1026), .B1(n_1027), .B2(n_1028), .C(n_1029), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_993), .A2(n_1504), .B1(n_1505), .B2(n_1506), .Y(n_1503) );
OAI22xp5_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_996), .B1(n_1001), .B2(n_1004), .Y(n_994) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_1003), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1012), .B(n_1015), .Y(n_1010) );
INVx8_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
AO22x2_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1066), .B1(n_1067), .B2(n_1115), .Y(n_1017) );
INVx1_ASAP7_75t_SL g1115 ( .A(n_1018), .Y(n_1115) );
XNOR2x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
NOR2x1_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1024), .Y(n_1020) );
NAND3xp33_ASAP7_75t_SL g1024 ( .A(n_1025), .B(n_1030), .C(n_1051), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1048), .B(n_1050), .Y(n_1030) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1039), .C(n_1043), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B(n_1046), .C(n_1047), .Y(n_1043) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1053), .Y(n_1089) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
AOI33xp33_ASAP7_75t_L g1242 ( .A1(n_1064), .A2(n_1243), .A3(n_1244), .B1(n_1247), .B2(n_1248), .B3(n_1249), .Y(n_1242) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
AOI33xp33_ASAP7_75t_L g1493 ( .A1(n_1065), .A2(n_1494), .A3(n_1496), .B1(n_1498), .B2(n_1499), .B3(n_1500), .Y(n_1493) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
NAND3xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1079), .C(n_1104), .Y(n_1069) );
NOR2xp33_ASAP7_75t_SL g1079 ( .A(n_1080), .B(n_1098), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1081) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_1086), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1560 ( .A1(n_1089), .A2(n_1133), .B1(n_1550), .B2(n_1556), .Y(n_1560) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_1118), .A2(n_1119), .B1(n_1175), .B2(n_1176), .Y(n_1117) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1119), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1158), .C(n_1167), .Y(n_1120) );
NOR2xp33_ASAP7_75t_SL g1121 ( .A(n_1122), .B(n_1141), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_1124), .A2(n_1139), .B1(n_1144), .B2(n_1145), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_1126), .A2(n_1140), .B1(n_1145), .B2(n_1150), .Y(n_1149) );
OAI22xp33_ASAP7_75t_SL g1127 ( .A1(n_1128), .A2(n_1129), .B1(n_1132), .B2(n_1133), .Y(n_1127) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_1144), .A2(n_1145), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_1144), .A2(n_1208), .B1(n_1209), .B2(n_1211), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1545 ( .A1(n_1144), .A2(n_1145), .B1(n_1546), .B2(n_1547), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g1554 ( .A1(n_1144), .A2(n_1209), .B1(n_1555), .B2(n_1556), .Y(n_1554) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_1150), .A2(n_1204), .B1(n_1205), .B2(n_1206), .Y(n_1203) );
INVx3_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1178), .B1(n_1218), .B2(n_1266), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
BUFx3_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
NAND3xp33_ASAP7_75t_SL g1181 ( .A(n_1182), .B(n_1189), .C(n_1195), .Y(n_1181) );
NOR2xp33_ASAP7_75t_SL g1195 ( .A(n_1196), .B(n_1212), .Y(n_1195) );
BUFx3_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_SL g1266 ( .A(n_1218), .Y(n_1266) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NAND3x1_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1242), .C(n_1252), .Y(n_1220) );
NAND3xp33_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1239), .C(n_1241), .Y(n_1234) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx2_ASAP7_75t_R g1497 ( .A(n_1246), .Y(n_1497) );
HB1xp67_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_SL g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_1269), .A2(n_1481), .B1(n_1484), .B2(n_1527), .C(n_1532), .Y(n_1268) );
NOR3xp33_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1418), .C(n_1457), .Y(n_1269) );
NAND3xp33_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1353), .C(n_1385), .Y(n_1270) );
AOI211xp5_ASAP7_75t_L g1271 ( .A1(n_1272), .A2(n_1297), .B(n_1314), .C(n_1333), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1272), .B(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1272), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1288), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1273), .B(n_1294), .Y(n_1401) );
NAND3xp33_ASAP7_75t_L g1405 ( .A(n_1273), .B(n_1391), .C(n_1406), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1273), .B(n_1323), .Y(n_1411) );
OR2x2_ASAP7_75t_L g1429 ( .A(n_1273), .B(n_1294), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1273), .B(n_1386), .Y(n_1443) );
CKINVDCx6p67_ASAP7_75t_R g1273 ( .A(n_1274), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1274), .B(n_1294), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1392 ( .A(n_1274), .B(n_1393), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1274), .B(n_1323), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1274), .B(n_1294), .Y(n_1422) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_1274), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_1274), .B(n_1348), .Y(n_1450) );
OR2x6_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1282), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1434 ( .A(n_1275), .B(n_1282), .Y(n_1434) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1276), .Y(n_1351) );
AND2x6_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1277), .B(n_1281), .Y(n_1280) );
AND2x4_ASAP7_75t_L g1283 ( .A(n_1277), .B(n_1284), .Y(n_1283) );
AND2x6_ASAP7_75t_L g1286 ( .A(n_1277), .B(n_1287), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1277), .B(n_1281), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1277), .B(n_1281), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1279), .B(n_1285), .Y(n_1284) );
INVx2_ASAP7_75t_L g1483 ( .A(n_1286), .Y(n_1483) );
HB1xp67_ASAP7_75t_L g1582 ( .A(n_1287), .Y(n_1582) );
AOI21xp33_ASAP7_75t_L g1370 ( .A1(n_1288), .A2(n_1347), .B(n_1371), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1288), .B(n_1318), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1293), .Y(n_1288) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1289), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1289), .B(n_1294), .Y(n_1335) );
OR2x2_ASAP7_75t_L g1384 ( .A(n_1289), .B(n_1294), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_1289), .B(n_1304), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1292), .Y(n_1289) );
INVxp67_ASAP7_75t_L g1352 ( .A(n_1291), .Y(n_1352) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
OAI221xp5_ASAP7_75t_L g1314 ( .A1(n_1294), .A2(n_1315), .B1(n_1319), .B2(n_1325), .C(n_1331), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1294), .B(n_1324), .Y(n_1346) );
A2O1A1Ixp33_ASAP7_75t_L g1353 ( .A1(n_1294), .A2(n_1354), .B(n_1368), .C(n_1369), .Y(n_1353) );
INVx3_ASAP7_75t_L g1414 ( .A(n_1294), .Y(n_1414) );
O2A1O1Ixp33_ASAP7_75t_L g1458 ( .A1(n_1294), .A2(n_1459), .B(n_1460), .C(n_1461), .Y(n_1458) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1294), .B(n_1304), .Y(n_1472) );
AND2x4_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1296), .Y(n_1294) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
AOI21xp5_ASAP7_75t_L g1461 ( .A1(n_1298), .A2(n_1384), .B(n_1462), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1303), .Y(n_1298) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1299), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1299), .B(n_1328), .Y(n_1332) );
BUFx2_ASAP7_75t_L g1359 ( .A(n_1299), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1299), .B(n_1307), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1299), .B(n_1373), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1301), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1307), .Y(n_1303) );
INVx2_ASAP7_75t_L g1318 ( .A(n_1304), .Y(n_1318) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1304), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1304), .B(n_1359), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1304), .B(n_1377), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1304), .B(n_1427), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1304), .B(n_1328), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1307), .B(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1307), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1307), .B(n_1448), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1307), .B(n_1366), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1311), .Y(n_1307) );
INVx2_ASAP7_75t_L g1329 ( .A(n_1308), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1308), .B(n_1330), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1308), .B(n_1359), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1310), .Y(n_1308) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1311), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1311), .B(n_1316), .Y(n_1339) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1311), .B(n_1359), .Y(n_1358) );
AND3x1_ASAP7_75t_L g1362 ( .A(n_1311), .B(n_1316), .C(n_1329), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1311), .B(n_1359), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1311), .B(n_1329), .Y(n_1391) );
OAI21xp33_ASAP7_75t_L g1423 ( .A1(n_1311), .A2(n_1424), .B(n_1425), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1317), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1316), .B(n_1326), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1316), .B(n_1328), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1316), .B(n_1373), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1316), .B(n_1329), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1316), .B(n_1318), .Y(n_1448) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1318), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1318), .B(n_1373), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1318), .B(n_1380), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1318), .B(n_1377), .Y(n_1399) );
O2A1O1Ixp33_ASAP7_75t_L g1408 ( .A1(n_1318), .A2(n_1342), .B(n_1409), .C(n_1410), .Y(n_1408) );
NOR2xp33_ASAP7_75t_L g1417 ( .A(n_1318), .B(n_1358), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1318), .B(n_1323), .Y(n_1432) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1322), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
OAI21xp33_ASAP7_75t_L g1402 ( .A1(n_1321), .A2(n_1403), .B(n_1405), .Y(n_1402) );
OAI222xp33_ASAP7_75t_L g1451 ( .A1(n_1321), .A2(n_1410), .B1(n_1452), .B2(n_1453), .C1(n_1454), .C2(n_1456), .Y(n_1451) );
OAI211xp5_ASAP7_75t_L g1354 ( .A1(n_1322), .A2(n_1355), .B(n_1360), .C(n_1363), .Y(n_1354) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1322), .Y(n_1416) );
O2A1O1Ixp33_ASAP7_75t_L g1437 ( .A1(n_1322), .A2(n_1378), .B(n_1404), .C(n_1438), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1322), .B(n_1480), .Y(n_1479) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1323), .B(n_1364), .Y(n_1363) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
OAI211xp5_ASAP7_75t_SL g1428 ( .A1(n_1325), .A2(n_1386), .B(n_1429), .C(n_1430), .Y(n_1428) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1326), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1328), .Y(n_1326) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1327), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1327), .B(n_1383), .Y(n_1382) );
NAND2xp5_ASAP7_75t_SL g1424 ( .A(n_1327), .B(n_1335), .Y(n_1424) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1328), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1328), .B(n_1382), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1328), .B(n_1448), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1330), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_1329), .B(n_1359), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1329), .B(n_1359), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1332), .Y(n_1456) );
O2A1O1Ixp33_ASAP7_75t_SL g1333 ( .A1(n_1334), .A2(n_1336), .B(n_1340), .C(n_1347), .Y(n_1333) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
OAI21xp5_ASAP7_75t_SL g1439 ( .A1(n_1335), .A2(n_1440), .B(n_1441), .Y(n_1439) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1338), .B(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
AOI21xp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1344), .B(n_1345), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
AOI221xp5_ASAP7_75t_L g1430 ( .A1(n_1344), .A2(n_1366), .B1(n_1391), .B2(n_1431), .C(n_1433), .Y(n_1430) );
AOI21xp33_ASAP7_75t_L g1438 ( .A1(n_1344), .A2(n_1345), .B(n_1409), .Y(n_1438) );
OAI21xp5_ASAP7_75t_L g1374 ( .A1(n_1346), .A2(n_1375), .B(n_1378), .Y(n_1374) );
CKINVDCx6p67_ASAP7_75t_R g1393 ( .A(n_1346), .Y(n_1393) );
INVx3_ASAP7_75t_L g1368 ( .A(n_1347), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1347), .B(n_1414), .Y(n_1413) );
INVx2_ASAP7_75t_SL g1347 ( .A(n_1348), .Y(n_1347) );
INVx2_ASAP7_75t_SL g1386 ( .A(n_1348), .Y(n_1386) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
NOR2xp33_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1357), .B(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1357), .Y(n_1397) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
A2O1A1Ixp33_ASAP7_75t_L g1470 ( .A1(n_1361), .A2(n_1414), .B(n_1449), .C(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_SL g1478 ( .A(n_1362), .B(n_1383), .Y(n_1478) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1363), .Y(n_1459) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1367), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1366), .B(n_1373), .Y(n_1440) );
O2A1O1Ixp33_ASAP7_75t_L g1446 ( .A1(n_1368), .A2(n_1383), .B(n_1447), .C(n_1449), .Y(n_1446) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1374), .C(n_1381), .Y(n_1369) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
OAI211xp5_ASAP7_75t_L g1436 ( .A1(n_1376), .A2(n_1393), .B(n_1437), .C(n_1439), .Y(n_1436) );
AOI211xp5_ASAP7_75t_L g1400 ( .A1(n_1378), .A2(n_1401), .B(n_1402), .C(n_1408), .Y(n_1400) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1380), .Y(n_1476) );
OAI21xp5_ASAP7_75t_L g1394 ( .A1(n_1383), .A2(n_1395), .B(n_1399), .Y(n_1394) );
INVx2_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
AOI22xp5_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1387), .B1(n_1412), .B2(n_1415), .Y(n_1385) );
NAND3xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1394), .C(n_1400), .Y(n_1387) );
INVxp67_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1392), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
AOI211xp5_ASAP7_75t_L g1464 ( .A1(n_1395), .A2(n_1414), .B(n_1465), .C(n_1467), .Y(n_1464) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1398), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1398), .B(n_1431), .Y(n_1466) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1398), .Y(n_1475) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVxp33_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1417), .Y(n_1415) );
AOI21xp5_ASAP7_75t_L g1477 ( .A1(n_1416), .A2(n_1460), .B(n_1478), .Y(n_1477) );
AOI221xp5_ASAP7_75t_SL g1418 ( .A1(n_1419), .A2(n_1434), .B1(n_1435), .B2(n_1442), .C(n_1444), .Y(n_1418) );
O2A1O1Ixp33_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1422), .B(n_1423), .C(n_1428), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVxp67_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
AOI211xp5_ASAP7_75t_L g1444 ( .A1(n_1436), .A2(n_1445), .B(n_1446), .C(n_1451), .Y(n_1444) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1440), .Y(n_1452) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
A2O1A1Ixp33_ASAP7_75t_L g1457 ( .A1(n_1445), .A2(n_1458), .B(n_1464), .C(n_1470), .Y(n_1457) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
CKINVDCx14_ASAP7_75t_R g1454 ( .A(n_1455), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1455), .B(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVxp67_ASAP7_75t_SL g1467 ( .A(n_1468), .Y(n_1467) );
OAI211xp5_ASAP7_75t_SL g1471 ( .A1(n_1472), .A2(n_1473), .B(n_1477), .C(n_1479), .Y(n_1471) );
INVxp67_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
NAND2xp5_ASAP7_75t_SL g1474 ( .A(n_1475), .B(n_1476), .Y(n_1474) );
CKINVDCx20_ASAP7_75t_R g1481 ( .A(n_1482), .Y(n_1481) );
CKINVDCx20_ASAP7_75t_R g1482 ( .A(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
HB1xp67_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1507), .Y(n_1487) );
NAND3xp33_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .C(n_1503), .Y(n_1491) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
AOI21xp5_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1521), .B(n_1522), .Y(n_1507) );
NAND3xp33_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1513), .C(n_1518), .Y(n_1508) );
CKINVDCx20_ASAP7_75t_R g1527 ( .A(n_1528), .Y(n_1527) );
CKINVDCx20_ASAP7_75t_R g1528 ( .A(n_1529), .Y(n_1528) );
INVx3_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
HB1xp67_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
BUFx3_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVxp33_ASAP7_75t_SL g1538 ( .A(n_1539), .Y(n_1538) );
HB1xp67_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
NAND3xp33_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1563), .C(n_1572), .Y(n_1541) );
NOR2xp33_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1557), .Y(n_1542) );
HB1xp67_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx2_ASAP7_75t_SL g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
OAI21xp5_ASAP7_75t_L g1581 ( .A1(n_1582), .A2(n_1583), .B(n_1584), .Y(n_1581) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
endmodule