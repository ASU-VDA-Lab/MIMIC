module real_aes_1586_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_666;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_749;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_0), .A2(n_138), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_1), .A2(n_44), .B1(n_428), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_2), .A2(n_93), .B1(n_543), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_3), .A2(n_7), .B1(n_560), .B2(n_772), .Y(n_771) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_4), .A2(n_199), .B1(n_288), .B2(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g746 ( .A(n_4), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_5), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_6), .A2(n_17), .B1(n_378), .B2(n_599), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_8), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_9), .A2(n_180), .B1(n_377), .B2(n_378), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_10), .A2(n_71), .B1(n_339), .B2(n_491), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_11), .A2(n_46), .B1(n_720), .B2(n_722), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_12), .A2(n_122), .B1(n_319), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_13), .A2(n_255), .B1(n_457), .B2(n_607), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_14), .A2(n_147), .B1(n_310), .B2(n_429), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_15), .A2(n_246), .B1(n_533), .B2(n_619), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_16), .B(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_18), .A2(n_238), .B1(n_537), .B2(n_538), .Y(n_691) );
AOI22x1_ASAP7_75t_L g694 ( .A1(n_19), .A2(n_119), .B1(n_425), .B2(n_545), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_20), .A2(n_115), .B1(n_387), .B2(n_388), .Y(n_386) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_21), .A2(n_66), .B1(n_288), .B2(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_21), .B(n_745), .Y(n_744) );
AO222x2_ASAP7_75t_L g615 ( .A1(n_22), .A2(n_65), .B1(n_222), .B2(n_407), .C1(n_530), .C2(n_533), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_23), .A2(n_123), .B1(n_341), .B2(n_490), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_24), .A2(n_223), .B1(n_537), .B2(n_538), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_25), .A2(n_148), .B1(n_332), .B2(n_445), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_26), .A2(n_141), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_27), .A2(n_190), .B1(n_319), .B2(n_377), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_28), .A2(n_263), .B1(n_447), .B2(n_448), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_29), .A2(n_226), .B1(n_310), .B2(n_381), .Y(n_380) );
XNOR2xp5_ASAP7_75t_L g678 ( .A(n_30), .B(n_679), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_30), .B(n_679), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_31), .A2(n_35), .B1(n_545), .B2(n_546), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_32), .A2(n_45), .B1(n_310), .B2(n_385), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_33), .A2(n_221), .B1(n_313), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_34), .A2(n_233), .B1(n_412), .B2(n_413), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_36), .A2(n_218), .B1(n_424), .B2(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_37), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_38), .A2(n_118), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_39), .A2(n_217), .B1(n_559), .B2(n_560), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_40), .A2(n_250), .B1(n_532), .B2(n_533), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_41), .B(n_369), .Y(n_368) );
OA22x2_ASAP7_75t_L g467 ( .A1(n_42), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_42), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_43), .A2(n_165), .B1(n_237), .B2(n_354), .C1(n_445), .C2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_47), .A2(n_104), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_48), .A2(n_171), .B1(n_317), .B2(n_455), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_49), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_50), .A2(n_161), .B1(n_372), .B2(n_643), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_51), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_52), .A2(n_265), .B1(n_484), .B2(n_486), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_53), .A2(n_264), .B1(n_364), .B2(n_559), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_54), .A2(n_146), .B1(n_484), .B2(n_486), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_55), .A2(n_254), .B1(n_445), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_56), .A2(n_186), .B1(n_442), .B2(n_444), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_57), .A2(n_638), .B1(n_639), .B2(n_653), .Y(n_637) );
INVxp67_ASAP7_75t_L g653 ( .A(n_57), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_58), .A2(n_214), .B1(n_410), .B2(n_413), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_59), .A2(n_149), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_60), .A2(n_259), .B1(n_724), .B2(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_61), .B(n_438), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_62), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_63), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_64), .A2(n_169), .B1(n_317), .B2(n_319), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_67), .A2(n_97), .B1(n_530), .B2(n_618), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_68), .A2(n_132), .B1(n_608), .B2(n_648), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_69), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_70), .A2(n_134), .B1(n_323), .B2(n_327), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_72), .A2(n_257), .B1(n_332), .B2(n_334), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_73), .A2(n_172), .B1(n_545), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_74), .A2(n_241), .B1(n_543), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_75), .A2(n_236), .B1(n_537), .B2(n_538), .Y(n_673) );
AO21x1_ASAP7_75t_L g749 ( .A1(n_76), .A2(n_750), .B(n_757), .Y(n_749) );
INVx3_ASAP7_75t_L g288 ( .A(n_77), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_78), .A2(n_153), .B1(n_542), .B2(n_546), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_79), .A2(n_162), .B1(n_341), .B2(n_372), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_80), .A2(n_191), .B1(n_384), .B2(n_385), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_81), .A2(n_200), .B1(n_606), .B2(n_608), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_82), .A2(n_121), .B1(n_542), .B2(n_543), .Y(n_541) );
AO21x2_ASAP7_75t_L g713 ( .A1(n_83), .A2(n_714), .B(n_733), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_83), .B(n_716), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_84), .A2(n_85), .B1(n_478), .B2(n_480), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_86), .A2(n_253), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_87), .A2(n_133), .B1(n_341), .B2(n_417), .Y(n_804) );
AO222x2_ASAP7_75t_L g665 ( .A1(n_88), .A2(n_145), .B1(n_173), .B2(n_407), .C1(n_412), .C2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_89), .A2(n_203), .B1(n_381), .B2(n_721), .Y(n_776) );
INVx1_ASAP7_75t_L g711 ( .A(n_90), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_91), .A2(n_150), .B1(n_618), .B2(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_92), .Y(n_495) );
INVx1_ASAP7_75t_SL g293 ( .A(n_94), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_94), .B(n_129), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_95), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_96), .Y(n_683) );
INVx2_ASAP7_75t_L g754 ( .A(n_98), .Y(n_754) );
OA22x2_ASAP7_75t_L g277 ( .A1(n_99), .A2(n_278), .B1(n_279), .B2(n_280), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_99), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_100), .A2(n_140), .B1(n_384), .B2(n_385), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_101), .A2(n_243), .B1(n_417), .B2(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_102), .A2(n_234), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_103), .A2(n_247), .B1(n_542), .B2(n_543), .Y(n_676) );
OA22x2_ASAP7_75t_L g357 ( .A1(n_105), .A2(n_358), .B1(n_390), .B2(n_391), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_105), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_106), .A2(n_114), .B1(n_347), .B2(n_364), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_107), .A2(n_266), .B1(n_323), .B2(n_501), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_108), .A2(n_174), .B1(n_429), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_109), .A2(n_194), .B1(n_317), .B2(n_422), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_110), .A2(n_144), .B1(n_478), .B2(n_480), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_111), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_112), .A2(n_197), .B1(n_384), .B2(n_432), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_113), .A2(n_125), .B1(n_457), .B2(n_607), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_116), .A2(n_224), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_117), .A2(n_166), .B1(n_329), .B2(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_120), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_124), .A2(n_139), .B1(n_505), .B2(n_799), .Y(n_798) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_126), .A2(n_790), .B(n_806), .Y(n_789) );
INVx1_ASAP7_75t_L g808 ( .A(n_126), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_127), .A2(n_245), .B1(n_339), .B2(n_341), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_128), .A2(n_242), .B1(n_347), .B2(n_349), .Y(n_346) );
AO22x2_ASAP7_75t_L g287 ( .A1(n_129), .A2(n_210), .B1(n_288), .B2(n_289), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_130), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_131), .A2(n_229), .B1(n_431), .B2(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_135), .A2(n_155), .B1(n_349), .B2(n_559), .Y(n_594) );
AND2x2_ASAP7_75t_L g793 ( .A(n_136), .B(n_438), .Y(n_793) );
OA22x2_ASAP7_75t_L g433 ( .A1(n_137), .A2(n_434), .B1(n_435), .B2(n_461), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_137), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_142), .A2(n_167), .B1(n_381), .B2(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_143), .A2(n_160), .B1(n_364), .B2(n_365), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_151), .A2(n_220), .B1(n_372), .B2(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g294 ( .A(n_152), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_154), .B(n_354), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_156), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_157), .A2(n_159), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_158), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_163), .A2(n_178), .B1(n_625), .B2(n_628), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_164), .A2(n_212), .B1(n_417), .B2(n_418), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_168), .A2(n_209), .B1(n_317), .B2(n_455), .Y(n_704) );
INVx1_ASAP7_75t_L g402 ( .A(n_170), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_175), .A2(n_239), .B1(n_489), .B2(n_491), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_176), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_177), .A2(n_202), .B1(n_428), .B2(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_179), .A2(n_189), .B1(n_283), .B2(n_302), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_181), .A2(n_251), .B1(n_310), .B2(n_313), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_182), .A2(n_256), .B1(n_372), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_183), .A2(n_198), .B1(n_422), .B2(n_454), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_184), .A2(n_232), .B1(n_425), .B2(n_431), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_185), .A2(n_206), .B1(n_332), .B2(n_362), .Y(n_361) );
AO22x1_ASAP7_75t_L g794 ( .A1(n_187), .A2(n_248), .B1(n_442), .B2(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_188), .B(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_192), .A2(n_216), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_193), .A2(n_267), .B1(n_424), .B2(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_195), .B(n_369), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_196), .A2(n_215), .B1(n_347), .B2(n_349), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_201), .A2(n_759), .B1(n_760), .B2(n_784), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_201), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_204), .A2(n_231), .B1(n_431), .B2(n_781), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_205), .A2(n_225), .B1(n_546), .B2(n_625), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_207), .A2(n_268), .B1(n_313), .B2(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_208), .A2(n_612), .B1(n_613), .B2(n_630), .Y(n_611) );
INVx1_ASAP7_75t_L g630 ( .A(n_208), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_211), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_213), .A2(n_261), .B1(n_412), .B2(n_413), .Y(n_526) );
INVx1_ASAP7_75t_L g741 ( .A(n_219), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_219), .B(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_227), .A2(n_260), .B1(n_489), .B2(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g742 ( .A(n_228), .Y(n_742) );
AND2x2_ASAP7_75t_R g786 ( .A(n_228), .B(n_741), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_230), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_235), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_240), .A2(n_258), .B1(n_332), .B2(n_445), .Y(n_592) );
INVxp67_ASAP7_75t_L g756 ( .A(n_244), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_249), .A2(n_269), .B1(n_543), .B2(n_573), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_252), .B(n_556), .Y(n_729) );
XNOR2x1_ASAP7_75t_L g586 ( .A(n_262), .B(n_587), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_748), .B(n_749), .Y(n_270) );
AOI21xp33_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_579), .B(n_738), .Y(n_271) );
OR2x2_ASAP7_75t_L g748 ( .A(n_272), .B(n_579), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_395), .B2(n_396), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_357), .B1(n_393), .B2(n_394), .Y(n_276) );
INVx1_ASAP7_75t_L g393 ( .A(n_277), .Y(n_393) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2x1_ASAP7_75t_L g280 ( .A(n_281), .B(n_330), .Y(n_280) );
NAND4xp25_ASAP7_75t_L g281 ( .A(n_282), .B(n_309), .C(n_316), .D(n_322), .Y(n_281) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g387 ( .A(n_284), .Y(n_387) );
INVx3_ASAP7_75t_L g428 ( .A(n_284), .Y(n_428) );
INVx2_ASAP7_75t_SL g601 ( .A(n_284), .Y(n_601) );
INVx2_ASAP7_75t_L g648 ( .A(n_284), .Y(n_648) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g721 ( .A(n_285), .Y(n_721) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_295), .Y(n_285) );
AND2x2_ASAP7_75t_L g318 ( .A(n_286), .B(n_307), .Y(n_318) );
AND2x4_ASAP7_75t_L g340 ( .A(n_286), .B(n_315), .Y(n_340) );
AND2x2_ASAP7_75t_L g532 ( .A(n_286), .B(n_315), .Y(n_532) );
AND2x2_ASAP7_75t_SL g537 ( .A(n_286), .B(n_307), .Y(n_537) );
AND2x6_ASAP7_75t_L g545 ( .A(n_286), .B(n_295), .Y(n_545) );
AND2x2_ASAP7_75t_L g619 ( .A(n_286), .B(n_315), .Y(n_619) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
BUFx2_ASAP7_75t_L g320 ( .A(n_287), .Y(n_320) );
AND2x2_ASAP7_75t_L g345 ( .A(n_287), .B(n_291), .Y(n_345) );
INVx1_ASAP7_75t_L g289 ( .A(n_288), .Y(n_289) );
OAI22x1_ASAP7_75t_L g291 ( .A1(n_288), .A2(n_292), .B1(n_293), .B2(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_288), .Y(n_292) );
INVx2_ASAP7_75t_L g298 ( .A(n_288), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_288), .Y(n_301) );
AND2x4_ASAP7_75t_L g305 ( .A(n_290), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g326 ( .A(n_291), .B(n_306), .Y(n_326) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
AND2x4_ASAP7_75t_L g312 ( .A(n_295), .B(n_305), .Y(n_312) );
AND2x4_ASAP7_75t_L g325 ( .A(n_295), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g356 ( .A(n_295), .B(n_345), .Y(n_356) );
AND2x4_ASAP7_75t_L g407 ( .A(n_295), .B(n_345), .Y(n_407) );
AND2x2_ASAP7_75t_L g542 ( .A(n_295), .B(n_326), .Y(n_542) );
AND2x2_ASAP7_75t_L g573 ( .A(n_295), .B(n_326), .Y(n_573) );
AND2x2_ASAP7_75t_L g625 ( .A(n_295), .B(n_305), .Y(n_625) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g308 ( .A(n_297), .Y(n_308) );
AND2x4_ASAP7_75t_L g315 ( .A(n_297), .B(n_299), .Y(n_315) );
AND2x2_ASAP7_75t_L g321 ( .A(n_297), .B(n_300), .Y(n_321) );
INVxp67_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g307 ( .A(n_300), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g381 ( .A(n_303), .Y(n_381) );
INVx2_ASAP7_75t_L g429 ( .A(n_303), .Y(n_429) );
INVx2_ASAP7_75t_L g508 ( .A(n_303), .Y(n_508) );
INVx2_ASAP7_75t_SL g567 ( .A(n_303), .Y(n_567) );
INVx2_ASAP7_75t_SL g602 ( .A(n_303), .Y(n_602) );
INVx2_ASAP7_75t_L g722 ( .A(n_303), .Y(n_722) );
INVx2_ASAP7_75t_L g799 ( .A(n_303), .Y(n_799) );
INVx8_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AND2x4_ASAP7_75t_L g314 ( .A(n_305), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g329 ( .A(n_305), .B(n_321), .Y(n_329) );
AND2x4_ASAP7_75t_L g543 ( .A(n_305), .B(n_321), .Y(n_543) );
AND2x6_ASAP7_75t_L g546 ( .A(n_305), .B(n_307), .Y(n_546) );
AND2x2_ASAP7_75t_L g628 ( .A(n_305), .B(n_315), .Y(n_628) );
AND2x2_ASAP7_75t_L g348 ( .A(n_307), .B(n_326), .Y(n_348) );
AND2x4_ASAP7_75t_L g618 ( .A(n_307), .B(n_326), .Y(n_618) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx3_ASAP7_75t_SL g431 ( .A(n_311), .Y(n_431) );
INVx2_ASAP7_75t_SL g452 ( .A(n_311), .Y(n_452) );
INVx2_ASAP7_75t_L g571 ( .A(n_311), .Y(n_571) );
INVx4_ASAP7_75t_L g607 ( .A(n_311), .Y(n_607) );
INVx8_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_313), .Y(n_781) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g389 ( .A(n_314), .Y(n_389) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_314), .Y(n_425) );
BUFx3_ASAP7_75t_L g608 ( .A(n_314), .Y(n_608) );
AND2x2_ASAP7_75t_L g333 ( .A(n_315), .B(n_326), .Y(n_333) );
AND2x4_ASAP7_75t_L g412 ( .A(n_315), .B(n_326), .Y(n_412) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g377 ( .A(n_318), .Y(n_377) );
INVx2_ASAP7_75t_L g515 ( .A(n_318), .Y(n_515) );
INVx5_ASAP7_75t_SL g379 ( .A(n_319), .Y(n_379) );
BUFx2_ASAP7_75t_L g422 ( .A(n_319), .Y(n_422) );
BUFx3_ASAP7_75t_L g778 ( .A(n_319), .Y(n_778) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x4_ASAP7_75t_L g538 ( .A(n_320), .B(n_321), .Y(n_538) );
AND2x2_ASAP7_75t_L g336 ( .A(n_321), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_321), .B(n_337), .Y(n_413) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_321), .B(n_337), .Y(n_666) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_324), .A2(n_458), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx3_ASAP7_75t_L g783 ( .A(n_324), .Y(n_783) );
INVx6_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g424 ( .A(n_325), .Y(n_424) );
BUFx3_ASAP7_75t_L g651 ( .A(n_325), .Y(n_651) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_SL g460 ( .A(n_328), .Y(n_460) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx3_ASAP7_75t_L g385 ( .A(n_329), .Y(n_385) );
BUFx3_ASAP7_75t_L g432 ( .A(n_329), .Y(n_432) );
BUFx2_ASAP7_75t_SL g501 ( .A(n_329), .Y(n_501) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_329), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g330 ( .A(n_331), .B(n_338), .C(n_346), .D(n_353), .Y(n_330) );
BUFx5_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g443 ( .A(n_333), .Y(n_443) );
BUFx3_ASAP7_75t_L g481 ( .A(n_333), .Y(n_481) );
INVx2_ASAP7_75t_L g554 ( .A(n_333), .Y(n_554) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
INVx3_ASAP7_75t_L g479 ( .A(n_335), .Y(n_479) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx12f_ASAP7_75t_L g445 ( .A(n_336), .Y(n_445) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
BUFx2_ASAP7_75t_L g417 ( .A(n_340), .Y(n_417) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_340), .Y(n_490) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g373 ( .A(n_342), .Y(n_373) );
INVx2_ASAP7_75t_L g418 ( .A(n_342), .Y(n_418) );
INVx1_ASAP7_75t_L g440 ( .A(n_342), .Y(n_440) );
INVx2_ASAP7_75t_L g491 ( .A(n_342), .Y(n_491) );
INVx2_ASAP7_75t_L g563 ( .A(n_342), .Y(n_563) );
INVx2_ASAP7_75t_L g643 ( .A(n_342), .Y(n_643) );
INVx6_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g533 ( .A(n_344), .B(n_345), .Y(n_533) );
AND2x4_ASAP7_75t_L g350 ( .A(n_345), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g530 ( .A(n_345), .B(n_351), .Y(n_530) );
AND2x2_ASAP7_75t_L g670 ( .A(n_345), .B(n_351), .Y(n_670) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_347), .Y(n_447) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g366 ( .A(n_348), .Y(n_366) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_348), .Y(n_559) );
BUFx4f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_SL g364 ( .A(n_350), .Y(n_364) );
BUFx3_ASAP7_75t_L g487 ( .A(n_350), .Y(n_487) );
INVx2_ASAP7_75t_L g561 ( .A(n_350), .Y(n_561) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g590 ( .A(n_354), .Y(n_590) );
INVx4_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g369 ( .A(n_355), .Y(n_369) );
INVx3_ASAP7_75t_SL g475 ( .A(n_355), .Y(n_475) );
INVx4_ASAP7_75t_SL g525 ( .A(n_355), .Y(n_525) );
INVx3_ASAP7_75t_L g556 ( .A(n_355), .Y(n_556) );
INVx6_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
INVx1_ASAP7_75t_L g656 ( .A(n_357), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_374), .Y(n_358) );
NOR3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_367), .C(n_370), .Y(n_359) );
NOR4xp25_ASAP7_75t_L g391 ( .A(n_360), .B(n_375), .C(n_382), .D(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_364), .Y(n_448) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g485 ( .A(n_366), .Y(n_485) );
INVx4_ASAP7_75t_L g529 ( .A(n_366), .Y(n_529) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_368), .B(n_371), .Y(n_392) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_369), .Y(n_438) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_382), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
BUFx2_ASAP7_75t_L g454 ( .A(n_377), .Y(n_454) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g455 ( .A(n_379), .Y(n_455) );
OAI22xp33_ASAP7_75t_SL g510 ( .A1(n_379), .A2(n_511), .B1(n_516), .B2(n_517), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .Y(n_382) );
BUFx2_ASAP7_75t_L g505 ( .A(n_387), .Y(n_505) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_463), .B(n_578), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_397), .B(n_465), .Y(n_578) );
AO22x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_433), .B2(n_462), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
XNOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
NAND2x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_419), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_405), .B(n_414), .Y(n_404) );
OAI21xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_408), .B(n_409), .Y(n_405) );
OAI222xp33_ASAP7_75t_L g681 ( .A1(n_406), .A2(n_411), .B1(n_682), .B2(n_683), .C1(n_684), .C2(n_685), .Y(n_681) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g685 ( .A(n_413), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g458 ( .A(n_425), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g462 ( .A(n_433), .Y(n_462) );
INVx1_ASAP7_75t_L g461 ( .A(n_435), .Y(n_461) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_449), .Y(n_435) );
NAND4xp25_ASAP7_75t_SL g436 ( .A(n_437), .B(n_439), .C(n_441), .D(n_446), .Y(n_436) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g768 ( .A(n_444), .Y(n_768) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g796 ( .A(n_445), .Y(n_796) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .C(n_456), .D(n_459), .Y(n_449) );
INVx1_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OAI22x1_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_518), .B1(n_519), .B2(n_577), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g577 ( .A(n_467), .Y(n_577) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND3x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_492), .C(n_502), .Y(n_470) );
NOR2xp67_ASAP7_75t_SL g471 ( .A(n_472), .B(n_482), .Y(n_471) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_476), .B(n_477), .Y(n_472) );
OAI222xp33_ASAP7_75t_L g763 ( .A1(n_473), .A2(n_764), .B1(n_766), .B2(n_767), .C1(n_768), .C2(n_769), .Y(n_763) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_483), .B(n_488), .Y(n_482) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
OAI22xp33_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B1(n_507), .B2(n_509), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g599 ( .A(n_513), .Y(n_599) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g725 ( .A(n_515), .Y(n_725) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AO22x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_548), .B1(n_575), .B2(n_576), .Y(n_519) );
INVx1_ASAP7_75t_SL g576 ( .A(n_520), .Y(n_576) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_547), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_522), .B(n_534), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .Y(n_540) );
INVx2_ASAP7_75t_L g575 ( .A(n_548), .Y(n_575) );
XOR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_574), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_550), .B(n_564), .Y(n_549) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_553), .Y(n_765) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g710 ( .A(n_554), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
BUFx6f_ASAP7_75t_SL g772 ( .A(n_559), .Y(n_772) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
XNOR2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_635), .Y(n_579) );
AOI22xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_609), .B1(n_631), .B2(n_632), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g634 ( .A(n_585), .Y(n_634) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_596), .Y(n_587) );
NOR2xp67_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_610), .Y(n_631) );
BUFx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_621), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_654), .B1(n_736), .B2(n_737), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_SL g737 ( .A(n_637), .Y(n_737) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_640), .B(n_646), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .C(n_644), .D(n_645), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .C(n_650), .D(n_652), .Y(n_646) );
INVx1_ASAP7_75t_L g736 ( .A(n_654), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B1(n_658), .B2(n_735), .Y(n_654) );
INVx1_ASAP7_75t_SL g735 ( .A(n_655), .Y(n_735) );
BUFx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22x1_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_712), .B1(n_713), .B2(n_734), .Y(n_658) );
INVx2_ASAP7_75t_L g734 ( .A(n_659), .Y(n_734) );
XNOR2x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_698), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_678), .B(n_696), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_661), .B(n_697), .Y(n_696) );
XNOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_671), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_680), .B(n_689), .Y(n_679) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_686), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
XOR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_711), .Y(n_698) );
NAND4xp75_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .C(n_706), .D(n_709), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_728), .Y(n_716) );
NAND4xp25_ASAP7_75t_SL g717 ( .A(n_718), .B(n_719), .C(n_723), .D(n_726), .Y(n_717) );
BUFx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND4xp25_ASAP7_75t_SL g728 ( .A(n_729), .B(n_730), .C(n_731), .D(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_740), .B(n_744), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g751 ( .A(n_742), .Y(n_751) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
NOR2x1_ASAP7_75t_R g750 ( .A(n_751), .B(n_752), .Y(n_750) );
OR2x2_ASAP7_75t_L g812 ( .A(n_751), .B(n_753), .Y(n_812) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
OAI222xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_785), .B1(n_787), .B2(n_808), .C1(n_809), .C2(n_812), .Y(n_757) );
CKINVDCx16_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_762), .B(n_774), .Y(n_761) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_770), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_779), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_790), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_803), .Y(n_791) );
NOR3xp33_ASAP7_75t_SL g792 ( .A(n_793), .B(n_794), .C(n_797), .Y(n_792) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND4xp25_ASAP7_75t_L g797 ( .A(n_798), .B(n_800), .C(n_801), .D(n_802), .Y(n_797) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
CKINVDCx6p67_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
endmodule