module fake_jpeg_2277_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_38),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_35),
.C(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_50),
.B1(n_5),
.B2(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_48),
.B1(n_46),
.B2(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_67),
.B1(n_73),
.B2(n_9),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_51),
.B1(n_46),
.B2(n_52),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_55),
.C(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_8),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_7),
.B(n_8),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_10),
.C(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_70),
.B1(n_65),
.B2(n_11),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_9),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_84),
.B(n_12),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_10),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_84),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_99),
.B(n_92),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_17),
.C(n_23),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_94),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_87),
.B1(n_95),
.B2(n_91),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_99),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_97),
.B(n_91),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_89),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_93),
.B1(n_24),
.B2(n_25),
.Y(n_108)
);


endmodule