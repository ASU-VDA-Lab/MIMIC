module fake_jpeg_14245_n_567 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_567);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_567;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_77),
.Y(n_137)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_79),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_18),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_35),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_90),
.Y(n_152)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_25),
.B(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_93),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_96),
.B(n_102),
.Y(n_171)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_30),
.B(n_16),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_44),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_46),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_126),
.B(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_44),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_26),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_141),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_49),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_105),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_26),
.C(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_46),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_146),
.B(n_156),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_76),
.B(n_39),
.Y(n_156)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_56),
.Y(n_159)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_90),
.B(n_28),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_51),
.Y(n_208)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_103),
.B(n_28),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_50),
.Y(n_192)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_112),
.B(n_55),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_101),
.C(n_154),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_182),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_75),
.B1(n_88),
.B2(n_94),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_181),
.A2(n_145),
.B1(n_118),
.B2(n_148),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_111),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_183),
.A2(n_194),
.B(n_208),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_184),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_21),
.B1(n_22),
.B2(n_49),
.Y(n_185)
);

OAI22x1_ASAP7_75t_L g291 ( 
.A1(n_185),
.A2(n_197),
.B1(n_204),
.B2(n_211),
.Y(n_291)
);

BUFx16f_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_92),
.B1(n_57),
.B2(n_100),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g275 ( 
.A1(n_188),
.A2(n_140),
.A3(n_53),
.B1(n_52),
.B2(n_41),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_111),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_189),
.B(n_192),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_193),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_67),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

CKINVDCx12_ASAP7_75t_R g196 ( 
.A(n_110),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_196),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_125),
.A2(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_43),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_206),
.Y(n_252)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_80),
.B1(n_98),
.B2(n_59),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_202),
.A2(n_36),
.B1(n_42),
.B2(n_33),
.Y(n_287)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_139),
.A2(n_22),
.B1(n_34),
.B2(n_37),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_223),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_131),
.B(n_47),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_136),
.Y(n_207)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_37),
.B1(n_34),
.B2(n_43),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_128),
.A2(n_47),
.B1(n_51),
.B2(n_48),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_212),
.A2(n_219),
.B1(n_122),
.B2(n_147),
.Y(n_253)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_137),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_214),
.B(n_222),
.Y(n_289)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_160),
.A2(n_48),
.B1(n_33),
.B2(n_42),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_121),
.A2(n_89),
.B1(n_48),
.B2(n_52),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_220),
.A2(n_235),
.B1(n_162),
.B2(n_158),
.Y(n_264)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_157),
.B(n_50),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_110),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_226),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_33),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_171),
.B(n_1),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_231),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_130),
.B(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_130),
.B(n_3),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_115),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

CKINVDCx12_ASAP7_75t_R g234 ( 
.A(n_168),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_154),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_235)
);

NAND2x1_ASAP7_75t_SL g236 ( 
.A(n_137),
.B(n_102),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_70),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_245),
.C(n_247),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_176),
.B(n_164),
.C(n_64),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_206),
.A2(n_147),
.B1(n_122),
.B2(n_124),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_250),
.A2(n_284),
.B(n_256),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_164),
.C(n_64),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_194),
.C(n_178),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_208),
.A2(n_101),
.B(n_120),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_256),
.A2(n_183),
.B(n_177),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_188),
.A2(n_145),
.B1(n_159),
.B2(n_118),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_261),
.A2(n_270),
.B1(n_287),
.B2(n_229),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_228),
.A2(n_142),
.B1(n_147),
.B2(n_122),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_262),
.A2(n_177),
.B1(n_187),
.B2(n_200),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_264),
.A2(n_265),
.B1(n_275),
.B2(n_283),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_186),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_188),
.A2(n_162),
.B1(n_158),
.B2(n_148),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_274),
.B(n_3),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_42),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_232),
.B(n_42),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_198),
.B(n_191),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_178),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_188),
.A2(n_58),
.B(n_54),
.C(n_129),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_200),
.B1(n_179),
.B2(n_194),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_220),
.A2(n_95),
.B1(n_52),
.B2(n_54),
.Y(n_283)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_194),
.A2(n_58),
.A3(n_95),
.B1(n_42),
.B2(n_33),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_227),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_288),
.Y(n_310)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_294),
.B(n_329),
.C(n_4),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_313),
.C(n_245),
.Y(n_351)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_174),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_297),
.B(n_306),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_235),
.B1(n_230),
.B2(n_175),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_298),
.A2(n_311),
.B1(n_316),
.B2(n_320),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_247),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_300),
.A2(n_302),
.B(n_273),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_304),
.Y(n_342)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_305),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_244),
.B(n_186),
.Y(n_306)
);

INVx5_ASAP7_75t_SL g307 ( 
.A(n_258),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_307),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_291),
.A2(n_187),
.B1(n_217),
.B2(n_224),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_250),
.B(n_291),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_175),
.B1(n_221),
.B2(n_213),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_318),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_241),
.B(n_183),
.C(n_180),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_190),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_314),
.B(n_317),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_269),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_333),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_201),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_252),
.B(n_195),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_239),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_319),
.B(n_326),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_282),
.A2(n_207),
.B1(n_215),
.B2(n_184),
.Y(n_320)
);

BUFx12f_ASAP7_75t_SL g321 ( 
.A(n_271),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_321),
.B(n_328),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_252),
.B(n_199),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_327),
.Y(n_352)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_209),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_215),
.Y(n_327)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_237),
.Y(n_332)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_272),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_336),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_264),
.A2(n_193),
.B1(n_36),
.B2(n_33),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_243),
.B1(n_242),
.B2(n_267),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_272),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_339),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_290),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_238),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_343),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_293),
.B(n_263),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_345),
.B(n_351),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_346),
.A2(n_383),
.B1(n_311),
.B2(n_340),
.Y(n_393)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_255),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_348),
.A2(n_368),
.B(n_373),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_279),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_364),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_293),
.B(n_277),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_251),
.C(n_238),
.Y(n_364)
);

OAI32xp33_ASAP7_75t_L g366 ( 
.A1(n_308),
.A2(n_327),
.A3(n_312),
.B1(n_318),
.B2(n_323),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_376),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_260),
.B1(n_283),
.B2(n_242),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_377),
.B1(n_335),
.B2(n_300),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_274),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_302),
.A2(n_290),
.B(n_239),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_372),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_338),
.A2(n_243),
.B(n_254),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_308),
.B(n_288),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_267),
.B1(n_254),
.B2(n_249),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g378 ( 
.A(n_295),
.B(n_249),
.C(n_257),
.Y(n_378)
);

NOR4xp25_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g385 ( 
.A1(n_381),
.A2(n_307),
.B(n_5),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_248),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_6),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_322),
.A2(n_257),
.B1(n_248),
.B2(n_240),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_418),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_334),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_386),
.B(n_406),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_390),
.B1(n_395),
.B2(n_396),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_338),
.B1(n_299),
.B2(n_300),
.Y(n_390)
);

NAND2x1_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_292),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_392),
.A2(n_348),
.B(n_359),
.Y(n_449)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_393),
.Y(n_426)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_344),
.A2(n_310),
.B1(n_332),
.B2(n_325),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_344),
.A2(n_310),
.B1(n_325),
.B2(n_337),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_331),
.B1(n_324),
.B2(n_303),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_398),
.A2(n_399),
.B1(n_401),
.B2(n_380),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_368),
.B1(n_376),
.B2(n_350),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_330),
.B1(n_296),
.B2(n_333),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_400),
.A2(n_405),
.B1(n_420),
.B2(n_342),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_352),
.A2(n_336),
.B1(n_339),
.B2(n_240),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_345),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_411),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_305),
.B1(n_304),
.B2(n_223),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_223),
.Y(n_406)
);

XOR2x1_ASAP7_75t_L g453 ( 
.A(n_407),
.B(n_364),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_343),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_408)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_341),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_409),
.B(n_416),
.Y(n_428)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_347),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_415),
.Y(n_445)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_413),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_361),
.B(n_7),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_7),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g418 ( 
.A(n_361),
.Y(n_418)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_346),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_350),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_422),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_401),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_424),
.A2(n_429),
.B1(n_434),
.B2(n_439),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_360),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_414),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_389),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_412),
.B(n_388),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_430),
.B(n_359),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_351),
.C(n_378),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_392),
.C(n_404),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_402),
.A2(n_372),
.B(n_368),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_419),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_403),
.A2(n_365),
.B1(n_380),
.B2(n_374),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_435),
.A2(n_446),
.B1(n_447),
.B2(n_453),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_392),
.A2(n_348),
.B(n_365),
.Y(n_437)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_437),
.A2(n_432),
.B(n_440),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_391),
.A2(n_366),
.B1(n_361),
.B2(n_356),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_438),
.A2(n_450),
.B1(n_384),
.B2(n_393),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_405),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_443),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_389),
.A2(n_353),
.B(n_371),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_391),
.A2(n_356),
.B1(n_369),
.B2(n_374),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_389),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_449),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_384),
.A2(n_369),
.B1(n_371),
.B2(n_375),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_390),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_456),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_399),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_457),
.B(n_458),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_414),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_394),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_461),
.C(n_462),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_460),
.A2(n_480),
.B1(n_442),
.B2(n_439),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_410),
.C(n_403),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_433),
.B(n_395),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_463),
.B(n_468),
.Y(n_486)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_417),
.C(n_413),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_471),
.C(n_473),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_453),
.B(n_407),
.Y(n_468)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_396),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_398),
.C(n_357),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_355),
.C(n_357),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_432),
.C(n_452),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_423),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_428),
.Y(n_502)
);

FAx1_ASAP7_75t_SL g477 ( 
.A(n_436),
.B(n_437),
.CI(n_445),
.CON(n_477),
.SN(n_477)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_443),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_481),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_445),
.A2(n_400),
.B1(n_415),
.B2(n_420),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_411),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_465),
.A2(n_425),
.B1(n_442),
.B2(n_436),
.Y(n_482)
);

AOI322xp5_ASAP7_75t_L g517 ( 
.A1(n_482),
.A2(n_477),
.A3(n_375),
.B1(n_10),
.B2(n_12),
.C1(n_8),
.C2(n_14),
.Y(n_517)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_466),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_463),
.Y(n_508)
);

OAI22x1_ASAP7_75t_L g485 ( 
.A1(n_477),
.A2(n_447),
.B1(n_426),
.B2(n_444),
.Y(n_485)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_485),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_444),
.B(n_426),
.Y(n_487)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_487),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_489),
.B(n_9),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_461),
.A2(n_421),
.B(n_451),
.Y(n_490)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_490),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_443),
.C(n_450),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_496),
.C(n_497),
.Y(n_505)
);

NOR2x1_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_455),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_9),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_494),
.A2(n_502),
.B1(n_504),
.B2(n_472),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_454),
.B(n_424),
.C(n_451),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_456),
.B(n_452),
.C(n_355),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_478),
.B(n_434),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_459),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_458),
.C(n_473),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_514),
.C(n_516),
.Y(n_523)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_508),
.Y(n_525)
);

INVx13_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_489),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_512),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_469),
.B1(n_481),
.B2(n_471),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_522),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_455),
.C(n_475),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_492),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_467),
.C(n_468),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_517),
.A2(n_521),
.B1(n_500),
.B2(n_498),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_8),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_518),
.A2(n_519),
.B(n_498),
.Y(n_530)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_483),
.C(n_491),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_528),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_527),
.A2(n_535),
.B(n_520),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_483),
.C(n_501),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_530),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_518),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_533),
.B(n_537),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_495),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_536),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_511),
.A2(n_496),
.B(n_486),
.Y(n_535)
);

FAx1_ASAP7_75t_SL g536 ( 
.A(n_516),
.B(n_486),
.CI(n_497),
.CON(n_536),
.SN(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_501),
.C(n_495),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_534),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_539),
.B(n_548),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_540),
.A2(n_545),
.B(n_536),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_532),
.A2(n_520),
.B1(n_507),
.B2(n_511),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_541),
.A2(n_507),
.B1(n_531),
.B2(n_525),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_523),
.B(n_510),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_546),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_523),
.A2(n_526),
.B(n_531),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_508),
.C(n_512),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_524),
.B(n_519),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_537),
.C(n_524),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_552),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_542),
.A2(n_535),
.B(n_530),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_555),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_554),
.A2(n_547),
.B(n_544),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_546),
.B(n_522),
.C(n_536),
.Y(n_555)
);

INVx13_ASAP7_75t_L g556 ( 
.A(n_551),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_556),
.B(n_550),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_559),
.A2(n_551),
.B(n_509),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_560),
.B(n_561),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_562),
.B(n_557),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_563),
.B(n_558),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_521),
.B(n_12),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_10),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_567)
);


endmodule