module real_aes_9760_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_719;
wire n_465;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g829 ( .A(n_0), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_0), .A2(n_176), .B1(n_295), .B2(n_405), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g1488 ( .A1(n_1), .A2(n_48), .B1(n_806), .B2(n_923), .C(n_1489), .Y(n_1488) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_1), .A2(n_278), .B1(n_1500), .B2(n_1503), .Y(n_1499) );
AO221x1_ASAP7_75t_L g1213 ( .A1(n_2), .A2(n_170), .B1(n_1214), .B2(n_1220), .C(n_1223), .Y(n_1213) );
INVx1_ASAP7_75t_L g606 ( .A(n_3), .Y(n_606) );
INVx1_ASAP7_75t_L g959 ( .A(n_4), .Y(n_959) );
INVxp33_ASAP7_75t_L g599 ( .A(n_5), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_5), .A2(n_568), .B(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_6), .A2(n_188), .B1(n_368), .B2(n_376), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_6), .A2(n_188), .B1(n_453), .B2(n_454), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_7), .A2(n_119), .B1(n_433), .B2(n_434), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_7), .A2(n_119), .B1(n_453), .B2(n_1197), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_8), .Y(n_294) );
INVx1_ASAP7_75t_L g446 ( .A(n_8), .Y(n_446) );
AND2x2_ASAP7_75t_L g615 ( .A(n_8), .B(n_372), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_8), .B(n_209), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_9), .A2(n_101), .B1(n_585), .B2(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_9), .A2(n_101), .B1(n_1111), .B2(n_1113), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1251 ( .A1(n_10), .A2(n_127), .B1(n_1214), .B2(n_1222), .Y(n_1251) );
OAI21xp33_ASAP7_75t_SL g1527 ( .A1(n_11), .A2(n_818), .B(n_1528), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_11), .A2(n_135), .B1(n_434), .B2(n_1553), .Y(n_1552) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_12), .A2(n_39), .B1(n_438), .B2(n_1155), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_12), .A2(n_39), .B1(n_714), .B2(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g608 ( .A(n_13), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_13), .A2(n_279), .B1(n_623), .B2(n_630), .C(n_632), .Y(n_622) );
AOI221xp5_ASAP7_75t_SL g912 ( .A1(n_14), .A2(n_34), .B1(n_913), .B2(n_914), .C(n_915), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_14), .A2(n_34), .B1(n_454), .B2(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g1128 ( .A(n_15), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_16), .A2(n_217), .B1(n_422), .B2(n_426), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_16), .A2(n_217), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_17), .A2(n_268), .B1(n_455), .B2(n_757), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_17), .A2(n_268), .B1(n_368), .B2(n_376), .Y(n_809) );
INVx1_ASAP7_75t_L g1530 ( .A(n_18), .Y(n_1530) );
OAI222xp33_ASAP7_75t_L g1538 ( .A1(n_18), .A2(n_25), .B1(n_267), .B2(n_639), .C1(n_700), .C2(n_1539), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_19), .A2(n_212), .B1(n_353), .B2(n_775), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g920 ( .A1(n_19), .A2(n_212), .B1(n_722), .B2(n_921), .C(n_924), .Y(n_920) );
AO221x2_ASAP7_75t_L g1304 ( .A1(n_20), .A2(n_184), .B1(n_1220), .B2(n_1305), .C(n_1307), .Y(n_1304) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_21), .A2(n_89), .B1(n_552), .B2(n_553), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_21), .A2(n_89), .B1(n_577), .B2(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g325 ( .A(n_22), .Y(n_325) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_22), .B(n_1440), .Y(n_1502) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_23), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_23), .A2(n_264), .B1(n_664), .B2(n_680), .Y(n_679) );
INVxp33_ASAP7_75t_L g702 ( .A(n_24), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_24), .A2(n_243), .B1(n_743), .B2(n_760), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g1561 ( .A1(n_25), .A2(n_186), .B1(n_1558), .B2(n_1562), .Y(n_1561) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_26), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_27), .A2(n_242), .B1(n_473), .B2(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_27), .Y(n_516) );
INVx1_ASAP7_75t_L g1079 ( .A(n_28), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_28), .A2(n_123), .B1(n_664), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_29), .A2(n_205), .B1(n_494), .B2(n_496), .Y(n_493) );
OAI211xp5_ASAP7_75t_SL g500 ( .A1(n_29), .A2(n_388), .B(n_501), .C(n_504), .Y(n_500) );
BUFx2_ASAP7_75t_L g365 ( .A(n_30), .Y(n_365) );
BUFx2_ASAP7_75t_L g408 ( .A(n_30), .Y(n_408) );
INVx1_ASAP7_75t_L g444 ( .A(n_30), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_31), .A2(n_50), .B1(n_833), .B2(n_835), .Y(n_832) );
OAI211xp5_ASAP7_75t_L g870 ( .A1(n_31), .A2(n_388), .B(n_871), .C(n_874), .Y(n_870) );
INVx1_ASAP7_75t_L g1019 ( .A(n_32), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_32), .A2(n_229), .B1(n_437), .B2(n_806), .Y(n_1035) );
INVx1_ASAP7_75t_L g1072 ( .A(n_33), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_33), .A2(n_105), .B1(n_779), .B2(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1088 ( .A(n_35), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_35), .A2(n_49), .B1(n_585), .B2(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1131 ( .A(n_36), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_36), .A2(n_104), .B1(n_426), .B2(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1532 ( .A(n_37), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_37), .A2(n_186), .B1(n_295), .B2(n_405), .Y(n_1537) );
INVxp33_ASAP7_75t_L g601 ( .A(n_38), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_38), .A2(n_102), .B1(n_412), .B2(n_434), .C(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g1133 ( .A(n_40), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_40), .A2(n_159), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_41), .A2(n_192), .B1(n_426), .B2(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_41), .A2(n_192), .B1(n_484), .B2(n_485), .Y(n_483) );
INVxp33_ASAP7_75t_L g1183 ( .A(n_42), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_42), .A2(n_168), .B1(n_412), .B2(n_620), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_43), .A2(n_53), .B1(n_433), .B2(n_1153), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_43), .A2(n_53), .B1(n_492), .B2(n_1161), .Y(n_1160) );
INVxp33_ASAP7_75t_SL g525 ( .A(n_44), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_44), .A2(n_51), .B1(n_589), .B2(n_590), .Y(n_588) );
AO22x2_ASAP7_75t_L g1060 ( .A1(n_45), .A2(n_1061), .B1(n_1062), .B2(n_1115), .Y(n_1060) );
INVx1_ASAP7_75t_L g1115 ( .A(n_45), .Y(n_1115) );
INVx1_ASAP7_75t_L g547 ( .A(n_46), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_46), .A2(n_187), .B1(n_558), .B2(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g712 ( .A(n_47), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_47), .A2(n_155), .B1(n_729), .B2(n_739), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_48), .A2(n_64), .B1(n_1505), .B2(n_1507), .Y(n_1504) );
INVx1_ASAP7_75t_L g1081 ( .A(n_49), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_50), .A2(n_114), .B1(n_368), .B2(n_376), .Y(n_877) );
INVxp33_ASAP7_75t_SL g527 ( .A(n_51), .Y(n_527) );
INVx1_ASAP7_75t_L g1229 ( .A(n_52), .Y(n_1229) );
INVx1_ASAP7_75t_L g990 ( .A(n_54), .Y(n_990) );
OAI211xp5_ASAP7_75t_L g994 ( .A1(n_54), .A2(n_348), .B(n_818), .C(n_995), .Y(n_994) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_55), .B(n_310), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_56), .A2(n_156), .B1(n_426), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_56), .A2(n_156), .B1(n_496), .B2(n_743), .Y(n_742) );
INVxp33_ASAP7_75t_SL g534 ( .A(n_57), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_57), .A2(n_60), .B1(n_585), .B2(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g900 ( .A(n_58), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_58), .A2(n_202), .B1(n_940), .B2(n_941), .Y(n_939) );
XOR2xp5_ASAP7_75t_L g1521 ( .A(n_59), .B(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g529 ( .A(n_60), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_61), .Y(n_917) );
INVx1_ASAP7_75t_L g1071 ( .A(n_62), .Y(n_1071) );
AOI22xp33_ASAP7_75t_SL g1103 ( .A1(n_62), .A2(n_83), .B1(n_567), .B2(n_1104), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_63), .Y(n_1012) );
INVx1_ASAP7_75t_L g1485 ( .A(n_64), .Y(n_1485) );
AOI22xp33_ASAP7_75t_SL g1458 ( .A1(n_65), .A2(n_266), .B1(n_492), .B2(n_757), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_65), .A2(n_266), .B1(n_1471), .B2(n_1472), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_66), .A2(n_235), .B1(n_422), .B2(n_426), .Y(n_480) );
INVx1_ASAP7_75t_L g511 ( .A(n_66), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_67), .A2(n_91), .B1(n_353), .B2(n_358), .Y(n_767) );
INVx1_ASAP7_75t_L g788 ( .A(n_67), .Y(n_788) );
INVxp33_ASAP7_75t_L g1177 ( .A(n_68), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_68), .A2(n_100), .B1(n_484), .B2(n_714), .Y(n_1200) );
INVxp33_ASAP7_75t_SL g543 ( .A(n_69), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_69), .A2(n_150), .B1(n_552), .B2(n_562), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_70), .A2(n_258), .B1(n_775), .B2(n_776), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_70), .A2(n_258), .B1(n_722), .B2(n_735), .C(n_787), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_71), .A2(n_200), .B1(n_295), .B2(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_71), .A2(n_196), .B1(n_450), .B2(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g866 ( .A(n_72), .Y(n_866) );
OAI211xp5_ASAP7_75t_SL g881 ( .A1(n_72), .A2(n_609), .B(n_882), .C(n_884), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_73), .A2(n_227), .B1(n_1547), .B2(n_1549), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1555 ( .A1(n_73), .A2(n_237), .B1(n_1556), .B2(n_1558), .Y(n_1555) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_74), .A2(n_947), .B1(n_997), .B2(n_998), .Y(n_946) );
INVx1_ASAP7_75t_L g998 ( .A(n_74), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_75), .A2(n_79), .B1(n_368), .B2(n_376), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_75), .A2(n_79), .B1(n_453), .B2(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g330 ( .A(n_76), .Y(n_330) );
INVx1_ASAP7_75t_L g347 ( .A(n_77), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_77), .A2(n_137), .B1(n_433), .B2(n_434), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_78), .A2(n_251), .B1(n_722), .B2(n_725), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_78), .A2(n_251), .B1(n_746), .B2(n_749), .Y(n_745) );
INVxp67_ASAP7_75t_SL g1143 ( .A(n_80), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_80), .A2(n_160), .B1(n_664), .B2(n_666), .Y(n_1164) );
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_81), .A2(n_274), .B1(n_473), .B2(n_737), .Y(n_1029) );
AOI22xp33_ASAP7_75t_SL g1039 ( .A1(n_81), .A2(n_274), .B1(n_487), .B2(n_491), .Y(n_1039) );
INVx1_ASAP7_75t_L g1174 ( .A(n_82), .Y(n_1174) );
OAI222xp33_ASAP7_75t_L g1065 ( .A1(n_83), .A2(n_171), .B1(n_263), .B2(n_1066), .C1(n_1067), .C2(n_1069), .Y(n_1065) );
INVx1_ASAP7_75t_L g698 ( .A(n_84), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_85), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_86), .Y(n_896) );
AO221x1_ASAP7_75t_L g1258 ( .A1(n_87), .A2(n_133), .B1(n_1214), .B2(n_1222), .C(n_1259), .Y(n_1258) );
AO22x2_ASAP7_75t_L g1166 ( .A1(n_88), .A2(n_1167), .B1(n_1202), .B2(n_1203), .Y(n_1166) );
INVx1_ASAP7_75t_L g1202 ( .A(n_88), .Y(n_1202) );
INVxp33_ASAP7_75t_SL g1126 ( .A(n_90), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_90), .A2(n_178), .B1(n_433), .B2(n_434), .Y(n_1148) );
INVx1_ASAP7_75t_L g808 ( .A(n_91), .Y(n_808) );
AO22x2_ASAP7_75t_L g1004 ( .A1(n_92), .A2(n_1005), .B1(n_1045), .B2(n_1046), .Y(n_1004) );
INVxp67_ASAP7_75t_L g1045 ( .A(n_92), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_93), .A2(n_202), .B1(n_368), .B2(n_376), .Y(n_893) );
INVx1_ASAP7_75t_L g938 ( .A(n_93), .Y(n_938) );
AO221x1_ASAP7_75t_L g1254 ( .A1(n_94), .A2(n_172), .B1(n_1214), .B2(n_1222), .C(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g519 ( .A(n_95), .Y(n_519) );
INVx1_ASAP7_75t_L g363 ( .A(n_96), .Y(n_363) );
INVx1_ASAP7_75t_L g1440 ( .A(n_96), .Y(n_1440) );
INVx1_ASAP7_75t_L g506 ( .A(n_97), .Y(n_506) );
INVx1_ASAP7_75t_L g960 ( .A(n_98), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_99), .A2(n_111), .B1(n_556), .B2(n_558), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_99), .A2(n_111), .B1(n_571), .B2(n_574), .Y(n_570) );
INVx1_ASAP7_75t_L g1173 ( .A(n_100), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_102), .Y(n_604) );
INVx1_ASAP7_75t_L g782 ( .A(n_103), .Y(n_782) );
INVxp33_ASAP7_75t_SL g1125 ( .A(n_104), .Y(n_1125) );
INVx1_ASAP7_75t_L g1075 ( .A(n_105), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_106), .A2(n_152), .B1(n_491), .B2(n_492), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_106), .A2(n_152), .B1(n_368), .B2(n_376), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_107), .A2(n_122), .B1(n_414), .B2(n_419), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_107), .A2(n_122), .B1(n_664), .B2(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g988 ( .A(n_108), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_108), .A2(n_163), .B1(n_353), .B2(n_775), .Y(n_993) );
INVx1_ASAP7_75t_L g1008 ( .A(n_109), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g1044 ( .A1(n_109), .A2(n_245), .B1(n_757), .B2(n_758), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_110), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_112), .A2(n_145), .B1(n_1094), .B2(n_1098), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_112), .A2(n_145), .B1(n_1106), .B2(n_1108), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_113), .A2(n_220), .B1(n_422), .B2(n_1031), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_113), .A2(n_220), .B1(n_449), .B2(n_762), .Y(n_1038) );
INVx1_ASAP7_75t_L g831 ( .A(n_114), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_115), .A2(n_231), .B1(n_1214), .B2(n_1222), .Y(n_1269) );
INVx1_ASAP7_75t_L g530 ( .A(n_116), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_117), .A2(n_165), .B1(n_666), .B2(n_962), .Y(n_961) );
INVxp67_ASAP7_75t_SL g975 ( .A(n_117), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1534 ( .A1(n_118), .A2(n_141), .B1(n_353), .B2(n_775), .Y(n_1534) );
AOI22xp33_ASAP7_75t_SL g1551 ( .A1(n_118), .A2(n_141), .B1(n_552), .B2(n_556), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_120), .Y(n_1453) );
INVx1_ASAP7_75t_L g861 ( .A(n_121), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_121), .A2(n_143), .B1(n_353), .B2(n_775), .Y(n_879) );
INVx1_ASAP7_75t_L g1078 ( .A(n_123), .Y(n_1078) );
INVx1_ASAP7_75t_L g1261 ( .A(n_124), .Y(n_1261) );
INVx1_ASAP7_75t_L g286 ( .A(n_125), .Y(n_286) );
XNOR2xp5_ASAP7_75t_L g811 ( .A(n_126), .B(n_812), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_128), .A2(n_219), .B1(n_779), .B2(n_780), .C(n_781), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_128), .A2(n_219), .B1(n_757), .B2(n_758), .Y(n_797) );
INVx1_ASAP7_75t_L g773 ( .A(n_129), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_130), .A2(n_388), .B(n_951), .C(n_952), .Y(n_950) );
INVx1_ASAP7_75t_L g967 ( .A(n_130), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g1246 ( .A1(n_131), .A2(n_213), .B1(n_1238), .B2(n_1241), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_132), .A2(n_205), .B1(n_295), .B2(n_405), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_132), .A2(n_235), .B1(n_353), .B2(n_358), .Y(n_518) );
INVx1_ASAP7_75t_L g1260 ( .A(n_134), .Y(n_1260) );
INVxp67_ASAP7_75t_SL g1533 ( .A(n_135), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_136), .Y(n_1016) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_137), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_138), .A2(n_177), .B1(n_823), .B2(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g843 ( .A(n_138), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_139), .A2(n_189), .B1(n_1214), .B2(n_1222), .Y(n_1247) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_140), .A2(n_280), .B1(n_1238), .B2(n_1241), .Y(n_1270) );
INVx1_ASAP7_75t_L g689 ( .A(n_142), .Y(n_689) );
INVx1_ASAP7_75t_L g857 ( .A(n_143), .Y(n_857) );
CKINVDCx14_ASAP7_75t_R g764 ( .A(n_144), .Y(n_764) );
INVx1_ASAP7_75t_L g772 ( .A(n_146), .Y(n_772) );
INVx1_ASAP7_75t_L g1308 ( .A(n_147), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_148), .A2(n_237), .B1(n_1106), .B2(n_1108), .Y(n_1550) );
AOI22xp33_ASAP7_75t_SL g1559 ( .A1(n_148), .A2(n_227), .B1(n_578), .B2(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1178 ( .A(n_149), .Y(n_1178) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_150), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_151), .A2(n_158), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_151), .A2(n_158), .B1(n_453), .B2(n_487), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_153), .A2(n_200), .B1(n_353), .B2(n_358), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_153), .A2(n_234), .B1(n_437), .B2(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g531 ( .A(n_154), .Y(n_531) );
INVxp33_ASAP7_75t_L g707 ( .A(n_155), .Y(n_707) );
INVxp33_ASAP7_75t_L g1171 ( .A(n_157), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_157), .A2(n_167), .B1(n_453), .B2(n_492), .Y(n_1201) );
INVx1_ASAP7_75t_L g1132 ( .A(n_159), .Y(n_1132) );
INVxp33_ASAP7_75t_L g1142 ( .A(n_160), .Y(n_1142) );
INVx1_ASAP7_75t_L g1175 ( .A(n_161), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_162), .Y(n_897) );
INVx1_ASAP7_75t_L g981 ( .A(n_163), .Y(n_981) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_164), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_164), .A2(n_215), .B1(n_734), .B2(n_735), .Y(n_733) );
INVxp67_ASAP7_75t_SL g977 ( .A(n_165), .Y(n_977) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_166), .Y(n_916) );
INVxp33_ASAP7_75t_L g1170 ( .A(n_167), .Y(n_1170) );
INVxp33_ASAP7_75t_L g1185 ( .A(n_168), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_169), .A2(n_238), .B1(n_426), .B2(n_1150), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_169), .A2(n_238), .B1(n_485), .B2(n_1042), .Y(n_1195) );
INVx1_ASAP7_75t_L g1085 ( .A(n_171), .Y(n_1085) );
INVx1_ASAP7_75t_L g693 ( .A(n_173), .Y(n_693) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_174), .Y(n_288) );
AND3x2_ASAP7_75t_L g1218 ( .A(n_174), .B(n_286), .C(n_1219), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_174), .B(n_286), .Y(n_1226) );
INVx1_ASAP7_75t_L g1456 ( .A(n_175), .Y(n_1456) );
OAI221xp5_ASAP7_75t_L g1473 ( .A1(n_175), .A2(n_644), .B1(n_1474), .B2(n_1475), .C(n_1479), .Y(n_1473) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_176), .A2(n_244), .B1(n_358), .B2(n_776), .Y(n_880) );
INVx1_ASAP7_75t_L g850 ( .A(n_177), .Y(n_850) );
INVxp33_ASAP7_75t_SL g1129 ( .A(n_178), .Y(n_1129) );
INVx1_ASAP7_75t_L g321 ( .A(n_179), .Y(n_321) );
INVxp33_ASAP7_75t_SL g1145 ( .A(n_180), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_180), .A2(n_247), .B1(n_714), .B2(n_1159), .Y(n_1163) );
INVxp33_ASAP7_75t_L g1186 ( .A(n_181), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_181), .A2(n_185), .B1(n_422), .B2(n_426), .Y(n_1193) );
INVx2_ASAP7_75t_L g299 ( .A(n_182), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_183), .A2(n_522), .B1(n_593), .B2(n_594), .Y(n_521) );
INVxp67_ASAP7_75t_L g593 ( .A(n_183), .Y(n_593) );
INVx1_ASAP7_75t_L g1181 ( .A(n_185), .Y(n_1181) );
INVxp33_ASAP7_75t_SL g540 ( .A(n_187), .Y(n_540) );
INVx1_ASAP7_75t_L g954 ( .A(n_190), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_191), .A2(n_210), .B1(n_412), .B2(n_417), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_191), .A2(n_210), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_193), .A2(n_440), .B(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_193), .Y(n_662) );
INVx1_ASAP7_75t_L g1219 ( .A(n_194), .Y(n_1219) );
INVxp67_ASAP7_75t_SL g694 ( .A(n_195), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_195), .A2(n_233), .B1(n_755), .B2(n_758), .Y(n_754) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_196), .A2(n_383), .B(n_388), .C(n_395), .Y(n_382) );
INVx1_ASAP7_75t_L g648 ( .A(n_197), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_198), .A2(n_201), .B1(n_1460), .B2(n_1466), .Y(n_1459) );
INVx1_ASAP7_75t_L g1494 ( .A(n_198), .Y(n_1494) );
INVx1_ASAP7_75t_L g536 ( .A(n_199), .Y(n_536) );
INVx1_ASAP7_75t_L g1491 ( .A(n_201), .Y(n_1491) );
INVx1_ASAP7_75t_L g1025 ( .A(n_203), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_203), .A2(n_249), .B1(n_433), .B2(n_979), .Y(n_1034) );
INVxp33_ASAP7_75t_SL g1542 ( .A(n_204), .Y(n_1542) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_204), .A2(n_259), .B1(n_577), .B2(n_578), .Y(n_1563) );
INVx1_ASAP7_75t_L g1434 ( .A(n_206), .Y(n_1434) );
INVx1_ASAP7_75t_L g799 ( .A(n_207), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_208), .A2(n_277), .B1(n_295), .B2(n_405), .Y(n_949) );
INVx1_ASAP7_75t_L g965 ( .A(n_208), .Y(n_965) );
INVx1_ASAP7_75t_L g301 ( .A(n_209), .Y(n_301) );
INVx2_ASAP7_75t_L g372 ( .A(n_209), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g768 ( .A1(n_211), .A2(n_348), .B(n_769), .C(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g791 ( .A(n_211), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g1250 ( .A1(n_214), .A2(n_236), .B1(n_1238), .B2(n_1241), .Y(n_1250) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_215), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g595 ( .A(n_216), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g1011 ( .A(n_218), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_218), .A2(n_273), .B1(n_835), .B2(n_1042), .Y(n_1041) );
OAI211xp5_ASAP7_75t_L g1049 ( .A1(n_218), .A2(n_388), .B(n_1050), .C(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1256 ( .A(n_221), .Y(n_1256) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_222), .Y(n_696) );
INVx1_ASAP7_75t_L g646 ( .A(n_223), .Y(n_646) );
INVx1_ASAP7_75t_L g784 ( .A(n_224), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_225), .A2(n_275), .B1(n_491), .B2(n_758), .Y(n_1454) );
INVx1_ASAP7_75t_L g1476 ( .A(n_225), .Y(n_1476) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_226), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_228), .A2(n_348), .B(n_882), .C(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g927 ( .A(n_228), .Y(n_927) );
INVx1_ASAP7_75t_L g1023 ( .A(n_229), .Y(n_1023) );
OAI211xp5_ASAP7_75t_L g1055 ( .A1(n_229), .A2(n_348), .B(n_1056), .C(n_1058), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_230), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_232), .Y(n_898) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_233), .Y(n_704) );
INVx1_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_239), .A2(n_255), .B1(n_358), .B2(n_776), .Y(n_908) );
INVx1_ASAP7_75t_L g925 ( .A(n_239), .Y(n_925) );
INVx1_ASAP7_75t_L g953 ( .A(n_240), .Y(n_953) );
INVx1_ASAP7_75t_L g1450 ( .A(n_241), .Y(n_1450) );
AOI21xp33_ASAP7_75t_L g1481 ( .A1(n_241), .A2(n_841), .B(n_1112), .Y(n_1481) );
INVx1_ASAP7_75t_L g517 ( .A(n_242), .Y(n_517) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_243), .Y(n_697) );
INVx1_ASAP7_75t_L g864 ( .A(n_244), .Y(n_864) );
INVx1_ASAP7_75t_L g1009 ( .A(n_245), .Y(n_1009) );
XOR2x2_ASAP7_75t_L g1121 ( .A(n_246), .B(n_1122), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1137 ( .A(n_247), .Y(n_1137) );
INVx1_ASAP7_75t_L g1217 ( .A(n_248), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_248), .B(n_1228), .Y(n_1232) );
INVx1_ASAP7_75t_L g1020 ( .A(n_249), .Y(n_1020) );
INVx1_ASAP7_75t_L g505 ( .A(n_250), .Y(n_505) );
AO22x2_ASAP7_75t_L g889 ( .A1(n_252), .A2(n_890), .B1(n_891), .B2(n_943), .Y(n_889) );
INVxp67_ASAP7_75t_L g943 ( .A(n_252), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_253), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_254), .Y(n_635) );
INVx1_ASAP7_75t_L g901 ( .A(n_255), .Y(n_901) );
INVx1_ASAP7_75t_L g1457 ( .A(n_256), .Y(n_1457) );
OAI211xp5_ASAP7_75t_SL g1482 ( .A1(n_256), .A2(n_1483), .B(n_1484), .C(n_1490), .Y(n_1482) );
AO22x1_ASAP7_75t_L g1235 ( .A1(n_257), .A2(n_262), .B1(n_1222), .B2(n_1236), .Y(n_1235) );
INVxp33_ASAP7_75t_L g1541 ( .A(n_259), .Y(n_1541) );
INVx2_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
AO22x1_ASAP7_75t_L g1237 ( .A1(n_261), .A2(n_265), .B1(n_1238), .B2(n_1241), .Y(n_1237) );
XNOR2xp5_ASAP7_75t_L g1431 ( .A(n_262), .B(n_1432), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_262), .A2(n_1516), .B1(n_1520), .B2(n_1564), .Y(n_1515) );
INVx1_ASAP7_75t_L g1086 ( .A(n_263), .Y(n_1086) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_264), .Y(n_613) );
INVx1_ASAP7_75t_L g1529 ( .A(n_267), .Y(n_1529) );
BUFx3_ASAP7_75t_L g319 ( .A(n_269), .Y(n_319) );
INVx1_ASAP7_75t_L g346 ( .A(n_269), .Y(n_346) );
BUFx3_ASAP7_75t_L g320 ( .A(n_270), .Y(n_320) );
INVx1_ASAP7_75t_L g339 ( .A(n_270), .Y(n_339) );
INVx1_ASAP7_75t_L g983 ( .A(n_271), .Y(n_983) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_271), .A2(n_277), .B1(n_358), .B2(n_776), .Y(n_996) );
INVx1_ASAP7_75t_L g800 ( .A(n_272), .Y(n_800) );
INVx1_ASAP7_75t_L g1015 ( .A(n_273), .Y(n_1015) );
INVx1_ASAP7_75t_L g1478 ( .A(n_275), .Y(n_1478) );
INVx1_ASAP7_75t_L g603 ( .A(n_276), .Y(n_603) );
INVx1_ASAP7_75t_L g1487 ( .A(n_278), .Y(n_1487) );
INVx1_ASAP7_75t_L g607 ( .A(n_279), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_302), .B(n_1207), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
AND2x4_ASAP7_75t_L g1514 ( .A(n_284), .B(n_290), .Y(n_1514) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_SL g1519 ( .A(n_285), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_285), .B(n_287), .Y(n_1569) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_287), .B(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x6_ASAP7_75t_L g407 ( .A(n_292), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_292), .B(n_408), .Y(n_1543) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g430 ( .A(n_293), .B(n_301), .Y(n_430) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g841 ( .A(n_294), .B(n_371), .Y(n_841) );
INVx8_ASAP7_75t_L g535 ( .A(n_295), .Y(n_535) );
OR2x6_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
OR2x6_ASAP7_75t_L g405 ( .A(n_296), .B(n_370), .Y(n_405) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_296), .A2(n_430), .B(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_296), .Y(n_783) );
INVx2_ASAP7_75t_SL g790 ( .A(n_296), .Y(n_790) );
INVx2_ASAP7_75t_SL g853 ( .A(n_296), .Y(n_853) );
BUFx6f_ASAP7_75t_L g972 ( .A(n_296), .Y(n_972) );
INVx1_ASAP7_75t_L g987 ( .A(n_296), .Y(n_987) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g375 ( .A(n_298), .Y(n_375) );
AND2x4_ASAP7_75t_L g380 ( .A(n_298), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g387 ( .A(n_298), .Y(n_387) );
INVx1_ASAP7_75t_L g394 ( .A(n_298), .Y(n_394) );
AND2x2_ASAP7_75t_L g425 ( .A(n_298), .B(n_299), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_299), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g381 ( .A(n_299), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_299), .Y(n_386) );
INVx1_ASAP7_75t_L g399 ( .A(n_299), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_299), .Y(n_416) );
AND2x4_ASAP7_75t_L g398 ( .A(n_300), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_301), .B(n_402), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1539 ( .A(n_301), .B(n_402), .Y(n_1539) );
XNOR2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_1000), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_886), .B1(n_887), .B2(n_999), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_810), .B2(n_885), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_305), .A2(n_306), .B1(n_810), .B2(n_885), .Y(n_999) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
XOR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_686), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_520), .B1(n_684), .B2(n_685), .Y(n_307) );
INVx2_ASAP7_75t_L g684 ( .A(n_308), .Y(n_684) );
XOR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_468), .Y(n_308) );
NAND3x1_ASAP7_75t_L g310 ( .A(n_311), .B(n_366), .C(n_409), .Y(n_310) );
OAI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_352), .B(n_361), .Y(n_311) );
NAND3xp33_ASAP7_75t_SL g312 ( .A(n_313), .B(n_335), .C(n_348), .Y(n_312) );
AOI222xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_321), .B2(n_322), .C1(n_330), .C2(n_331), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g512 ( .A(n_316), .Y(n_512) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_SL g451 ( .A(n_317), .Y(n_451) );
BUFx3_ASAP7_75t_L g587 ( .A(n_317), .Y(n_587) );
BUFx4f_ASAP7_75t_L g714 ( .A(n_317), .Y(n_714) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_317), .Y(n_762) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g333 ( .A(n_319), .Y(n_333) );
AND2x4_ASAP7_75t_L g338 ( .A(n_319), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g329 ( .A(n_320), .Y(n_329) );
AND2x4_ASAP7_75t_L g345 ( .A(n_320), .B(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_321), .A2(n_330), .B1(n_396), .B2(n_400), .Y(n_395) );
AOI222xp33_ASAP7_75t_L g546 ( .A1(n_322), .A2(n_331), .B1(n_496), .B2(n_530), .C1(n_531), .C2(n_547), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_322), .A2(n_331), .B1(n_587), .B2(n_606), .C1(n_607), .C2(n_608), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g1130 ( .A1(n_322), .A2(n_331), .B1(n_574), .B2(n_1131), .C1(n_1132), .C2(n_1133), .Y(n_1130) );
AOI222xp33_ASAP7_75t_L g1180 ( .A1(n_322), .A2(n_331), .B1(n_574), .B2(n_1174), .C1(n_1175), .C2(n_1181), .Y(n_1180) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_323), .B(n_326), .Y(n_322) );
AND2x4_ASAP7_75t_L g359 ( .A(n_323), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g716 ( .A(n_323), .B(n_326), .Y(n_716) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g334 ( .A(n_325), .Y(n_334) );
INVx1_ASAP7_75t_L g343 ( .A(n_325), .Y(n_343) );
AND2x2_ASAP7_75t_L g459 ( .A(n_325), .B(n_363), .Y(n_459) );
INVx2_ASAP7_75t_L g467 ( .A(n_325), .Y(n_467) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g514 ( .A(n_327), .Y(n_514) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g1464 ( .A(n_328), .Y(n_1464) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g360 ( .A(n_329), .B(n_333), .Y(n_360) );
AOI222xp33_ASAP7_75t_L g510 ( .A1(n_331), .A2(n_505), .B1(n_506), .B2(n_511), .C1(n_512), .C2(n_513), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g711 ( .A1(n_331), .A2(n_696), .B1(n_698), .B2(n_712), .C1(n_713), .C2(n_715), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_331), .A2(n_716), .B1(n_772), .B2(n_773), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_331), .A2(n_716), .B1(n_875), .B2(n_876), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_331), .A2(n_715), .B1(n_896), .B2(n_898), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_331), .A2(n_716), .B1(n_953), .B2(n_954), .Y(n_995) );
AOI222xp33_ASAP7_75t_L g1021 ( .A1(n_331), .A2(n_715), .B1(n_1012), .B2(n_1013), .C1(n_1022), .C2(n_1023), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_331), .A2(n_716), .B1(n_1012), .B2(n_1013), .Y(n_1058) );
INVx3_ASAP7_75t_L g1069 ( .A(n_331), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1528 ( .A1(n_331), .A2(n_513), .B1(n_1529), .B2(n_1530), .Y(n_1528) );
AND2x6_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
BUFx3_ASAP7_75t_L g1468 ( .A(n_332), .Y(n_1468) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g337 ( .A(n_334), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B1(n_341), .B2(n_347), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_336), .A2(n_341), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_336), .A2(n_540), .B1(n_541), .B2(n_543), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_336), .A2(n_599), .B1(n_600), .B2(n_601), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_336), .A2(n_541), .B1(n_707), .B2(n_708), .Y(n_706) );
CKINVDCx6p67_ASAP7_75t_R g775 ( .A(n_336), .Y(n_775) );
AOI22xp5_ASAP7_75t_SL g1018 ( .A1(n_336), .A2(n_600), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_336), .A2(n_600), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_336), .A2(n_541), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_336), .A2(n_600), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
AND2x6_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g350 ( .A(n_337), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_337), .Y(n_354) );
AND2x2_ASAP7_75t_L g770 ( .A(n_337), .B(n_485), .Y(n_770) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_338), .Y(n_453) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_338), .Y(n_491) );
BUFx2_ASAP7_75t_L g577 ( .A(n_338), .Y(n_577) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_338), .Y(n_665) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_338), .Y(n_748) );
BUFx3_ASAP7_75t_L g757 ( .A(n_338), .Y(n_757) );
INVx2_ASAP7_75t_SL g963 ( .A(n_338), .Y(n_963) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_338), .Y(n_1098) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_338), .Y(n_1161) );
INVx1_ASAP7_75t_L g357 ( .A(n_339), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_341), .A2(n_359), .B1(n_536), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_341), .A2(n_359), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_341), .A2(n_359), .B1(n_693), .B2(n_710), .Y(n_709) );
INVx4_ASAP7_75t_L g776 ( .A(n_341), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_341), .A2(n_359), .B1(n_1016), .B2(n_1025), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_341), .A2(n_359), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_341), .A2(n_359), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_341), .A2(n_349), .B1(n_359), .B2(n_1178), .C(n_1183), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_341), .A2(n_359), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
AND2x6_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
AND2x4_ASAP7_75t_L g541 ( .A(n_342), .B(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g600 ( .A(n_342), .B(n_542), .Y(n_600) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g513 ( .A(n_343), .B(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_344), .Y(n_492) );
INVx1_ASAP7_75t_L g681 ( .A(n_344), .Y(n_681) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_344), .Y(n_758) );
INVx2_ASAP7_75t_L g826 ( .A(n_344), .Y(n_826) );
INVx1_ASAP7_75t_L g1198 ( .A(n_344), .Y(n_1198) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_345), .Y(n_455) );
INVx1_ASAP7_75t_L g488 ( .A(n_345), .Y(n_488) );
INVx1_ASAP7_75t_L g579 ( .A(n_345), .Y(n_579) );
INVx2_ASAP7_75t_L g669 ( .A(n_345), .Y(n_669) );
INVx1_ASAP7_75t_L g356 ( .A(n_346), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g509 ( .A(n_348), .B(n_510), .C(n_515), .Y(n_509) );
NAND4xp25_ASAP7_75t_SL g538 ( .A(n_348), .B(n_539), .C(n_544), .D(n_546), .Y(n_538) );
NAND4xp25_ASAP7_75t_L g1123 ( .A(n_348), .B(n_1124), .C(n_1127), .D(n_1130), .Y(n_1123) );
CKINVDCx8_ASAP7_75t_R g348 ( .A(n_349), .Y(n_348) );
INVx5_ASAP7_75t_L g609 ( .A(n_349), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g1064 ( .A(n_349), .B(n_1065), .Y(n_1064) );
NOR2xp33_ASAP7_75t_SL g1526 ( .A(n_349), .B(n_1527), .Y(n_1526) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_351), .Y(n_485) );
INVx2_ASAP7_75t_L g497 ( .A(n_351), .Y(n_497) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_351), .Y(n_575) );
INVx1_ASAP7_75t_L g836 ( .A(n_351), .Y(n_836) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g659 ( .A(n_355), .Y(n_659) );
INVx2_ASAP7_75t_L g675 ( .A(n_355), .Y(n_675) );
BUFx2_ASAP7_75t_L g817 ( .A(n_355), .Y(n_817) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g661 ( .A(n_356), .B(n_357), .Y(n_661) );
INVx4_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g449 ( .A(n_360), .Y(n_449) );
INVx2_ASAP7_75t_L g463 ( .A(n_360), .Y(n_463) );
INVx6_ASAP7_75t_L g495 ( .A(n_360), .Y(n_495) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_360), .B(n_1438), .Y(n_1437) );
OAI21xp5_ASAP7_75t_SL g508 ( .A1(n_361), .A2(n_509), .B(n_518), .Y(n_508) );
OAI31xp33_ASAP7_75t_L g766 ( .A1(n_361), .A2(n_767), .A3(n_768), .B(n_774), .Y(n_766) );
OAI31xp33_ASAP7_75t_SL g992 ( .A1(n_361), .A2(n_993), .A3(n_994), .B(n_996), .Y(n_992) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
AND2x4_ASAP7_75t_L g548 ( .A(n_362), .B(n_364), .Y(n_548) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g466 ( .A(n_363), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g1497 ( .A(n_364), .Y(n_1497) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g429 ( .A(n_365), .Y(n_429) );
OR2x6_ASAP7_75t_L g840 ( .A(n_365), .B(n_841), .Y(n_840) );
OAI31xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_382), .A3(n_404), .B(n_406), .Y(n_366) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g377 ( .A(n_370), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g526 ( .A(n_370), .B(n_414), .Y(n_526) );
AND2x4_ASAP7_75t_L g703 ( .A(n_370), .B(n_378), .Y(n_703) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
BUFx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g846 ( .A(n_374), .Y(n_846) );
INVx1_ASAP7_75t_L g860 ( .A(n_374), .Y(n_860) );
AND2x4_ASAP7_75t_L g414 ( .A(n_375), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g631 ( .A(n_375), .Y(n_631) );
INVx5_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_377), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_377), .A2(n_526), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_377), .A2(n_526), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
INVx1_ASAP7_75t_L g565 ( .A(n_380), .Y(n_565) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_380), .Y(n_737) );
AND2x4_ASAP7_75t_L g393 ( .A(n_381), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g865 ( .A(n_384), .Y(n_865) );
INVx1_ASAP7_75t_L g973 ( .A(n_384), .Y(n_973) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g503 ( .A(n_385), .Y(n_503) );
INVx3_ASAP7_75t_L g639 ( .A(n_385), .Y(n_639) );
INVx2_ASAP7_75t_L g989 ( .A(n_385), .Y(n_989) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_386), .B(n_387), .Y(n_873) );
INVx1_ASAP7_75t_L g402 ( .A(n_387), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g523 ( .A(n_388), .B(n_524), .C(n_528), .D(n_533), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_388), .B(n_692), .C(n_695), .D(n_701), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_388), .B(n_804), .C(n_807), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_388), .B(n_895), .C(n_899), .Y(n_894) );
NAND4xp25_ASAP7_75t_L g1006 ( .A(n_388), .B(n_1007), .C(n_1010), .D(n_1014), .Y(n_1006) );
NAND4xp25_ASAP7_75t_SL g1076 ( .A(n_388), .B(n_1077), .C(n_1080), .D(n_1087), .Y(n_1076) );
NAND4xp25_ASAP7_75t_L g1168 ( .A(n_388), .B(n_1169), .C(n_1172), .D(n_1176), .Y(n_1168) );
CKINVDCx11_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g1135 ( .A1(n_389), .A2(n_1136), .B(n_1137), .C(n_1138), .Y(n_1135) );
NOR3xp33_ASAP7_75t_L g1536 ( .A(n_389), .B(n_1537), .C(n_1538), .Y(n_1536) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g403 ( .A(n_391), .Y(n_403) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_392), .B(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_393), .Y(n_440) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_393), .Y(n_559) );
BUFx3_ASAP7_75t_L g806 ( .A(n_393), .Y(n_806) );
INVx1_ASAP7_75t_L g1032 ( .A(n_393), .Y(n_1032) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_393), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_396), .A2(n_400), .B1(n_953), .B2(n_954), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_396), .A2(n_400), .B1(n_1012), .B2(n_1013), .Y(n_1051) );
AOI222xp33_ASAP7_75t_L g1172 ( .A1(n_396), .A2(n_532), .B1(n_1084), .B2(n_1173), .C1(n_1174), .C2(n_1175), .Y(n_1172) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_398), .A2(n_400), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_398), .A2(n_440), .B1(n_529), .B2(n_530), .C1(n_531), .C2(n_532), .Y(n_528) );
INVx2_ASAP7_75t_L g700 ( .A(n_398), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g804 ( .A1(n_398), .A2(n_400), .B1(n_772), .B2(n_773), .C1(n_800), .C2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_398), .A2(n_400), .B1(n_875), .B2(n_876), .Y(n_874) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_398), .A2(n_400), .B1(n_559), .B2(n_896), .C1(n_897), .C2(n_898), .Y(n_895) );
INVx2_ASAP7_75t_L g1139 ( .A(n_398), .Y(n_1139) );
INVx1_ASAP7_75t_L g625 ( .A(n_399), .Y(n_625) );
HB1xp67_ASAP7_75t_L g1493 ( .A(n_399), .Y(n_1493) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_400), .A2(n_558), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_699), .Y(n_695) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
AND2x4_ASAP7_75t_L g532 ( .A(n_401), .B(n_403), .Y(n_532) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx4_ASAP7_75t_L g537 ( .A(n_405), .Y(n_537) );
INVx5_ASAP7_75t_L g902 ( .A(n_405), .Y(n_902) );
OAI31xp33_ASAP7_75t_SL g498 ( .A1(n_406), .A2(n_499), .A3(n_500), .B(n_507), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_406), .A2(n_523), .B1(n_538), .B2(n_548), .C(n_549), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_406), .A2(n_691), .B1(n_705), .B2(n_717), .C(n_719), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_406), .A2(n_803), .B(n_809), .Y(n_802) );
OAI31xp33_ASAP7_75t_SL g868 ( .A1(n_406), .A2(n_869), .A3(n_870), .B(n_877), .Y(n_868) );
O2A1O1Ixp33_ASAP7_75t_L g892 ( .A1(n_406), .A2(n_893), .B(n_894), .C(n_903), .Y(n_892) );
OAI31xp33_ASAP7_75t_L g948 ( .A1(n_406), .A2(n_949), .A3(n_950), .B(n_955), .Y(n_948) );
AOI221x1_ASAP7_75t_L g1005 ( .A1(n_406), .A2(n_610), .B1(n_1006), .B2(n_1017), .C(n_1026), .Y(n_1005) );
OAI31xp33_ASAP7_75t_L g1047 ( .A1(n_406), .A2(n_1048), .A3(n_1049), .B(n_1052), .Y(n_1047) );
AOI221x1_ASAP7_75t_L g1062 ( .A1(n_406), .A2(n_610), .B1(n_1063), .B2(n_1076), .C(n_1089), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_406), .A2(n_548), .B1(n_1123), .B2(n_1134), .C(n_1146), .Y(n_1122) );
AOI221x1_ASAP7_75t_L g1167 ( .A1(n_406), .A2(n_548), .B1(n_1168), .B2(n_1179), .C(n_1187), .Y(n_1167) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g465 ( .A(n_408), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g592 ( .A(n_408), .B(n_466), .Y(n_592) );
AND2x4_ASAP7_75t_L g1436 ( .A(n_408), .B(n_1437), .Y(n_1436) );
AND4x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_431), .C(n_447), .D(n_460), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_421), .C(n_428), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g552 ( .A(n_413), .Y(n_552) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_414), .Y(n_433) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
AND2x2_ASAP7_75t_L g614 ( .A(n_414), .B(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_414), .Y(n_724) );
BUFx2_ASAP7_75t_L g734 ( .A(n_414), .Y(n_734) );
BUFx2_ASAP7_75t_L g779 ( .A(n_414), .Y(n_779) );
INVx1_ASAP7_75t_L g1107 ( .A(n_414), .Y(n_1107) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g863 ( .A(n_417), .Y(n_863) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g554 ( .A(n_419), .Y(n_554) );
INVx1_ASAP7_75t_L g849 ( .A(n_419), .Y(n_849) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_420), .Y(n_435) );
INVx3_ASAP7_75t_L g727 ( .A(n_420), .Y(n_727) );
INVx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g476 ( .A(n_423), .Y(n_476) );
INVx2_ASAP7_75t_L g1150 ( .A(n_423), .Y(n_1150) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g437 ( .A(n_424), .Y(n_437) );
AND2x4_ASAP7_75t_L g649 ( .A(n_424), .B(n_615), .Y(n_649) );
BUFx6f_ASAP7_75t_L g923 ( .A(n_424), .Y(n_923) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g557 ( .A(n_425), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g1010 ( .A1(n_426), .A2(n_532), .B1(n_699), .B2(n_1011), .C1(n_1012), .C2(n_1013), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_426), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g647 ( .A(n_427), .B(n_618), .Y(n_647) );
INVx1_ASAP7_75t_L g1114 ( .A(n_427), .Y(n_1114) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_428), .B(n_472), .C(n_475), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_428), .B(n_551), .C(n_555), .Y(n_550) );
INVx2_ASAP7_75t_L g731 ( .A(n_428), .Y(n_731) );
BUFx3_ASAP7_75t_L g785 ( .A(n_428), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g1028 ( .A(n_428), .B(n_1029), .C(n_1030), .Y(n_1028) );
AOI33xp33_ASAP7_75t_L g1099 ( .A1(n_428), .A2(n_441), .A3(n_1100), .B1(n_1103), .B2(n_1105), .B3(n_1110), .Y(n_1099) );
NAND3xp33_ASAP7_75t_L g1151 ( .A(n_428), .B(n_1152), .C(n_1154), .Y(n_1151) );
NAND3xp33_ASAP7_75t_L g1188 ( .A(n_428), .B(n_1189), .C(n_1190), .Y(n_1188) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OR2x2_ASAP7_75t_L g457 ( .A(n_429), .B(n_458), .Y(n_457) );
OR2x6_ASAP7_75t_L g581 ( .A(n_429), .B(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g655 ( .A(n_429), .Y(n_655) );
OR2x2_ASAP7_75t_L g793 ( .A(n_429), .B(n_582), .Y(n_793) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_429), .B(n_642), .Y(n_1036) );
INVx2_ASAP7_75t_L g1442 ( .A(n_429), .Y(n_1442) );
AND2x4_ASAP7_75t_L g1545 ( .A(n_429), .B(n_430), .Y(n_1545) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .C(n_441), .Y(n_431) );
INVx1_ASAP7_75t_L g984 ( .A(n_434), .Y(n_984) );
INVx1_ASAP7_75t_L g1477 ( .A(n_434), .Y(n_1477) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx2_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
INVx3_ASAP7_75t_L g979 ( .A(n_435), .Y(n_979) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_440), .Y(n_1104) );
BUFx2_ASAP7_75t_L g1553 ( .A(n_440), .Y(n_1553) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_441), .B(n_561), .C(n_566), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_441), .B(n_733), .C(n_738), .Y(n_732) );
CKINVDCx8_ASAP7_75t_R g867 ( .A(n_441), .Y(n_867) );
NAND3xp33_ASAP7_75t_L g1147 ( .A(n_441), .B(n_1148), .C(n_1149), .Y(n_1147) );
INVx5_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx6_ASAP7_75t_L g481 ( .A(n_442), .Y(n_481) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g1447 ( .A(n_443), .B(n_1438), .Y(n_1447) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_444), .B(n_1502), .Y(n_1501) );
INVx2_ASAP7_75t_L g642 ( .A(n_445), .Y(n_642) );
BUFx2_ASAP7_75t_L g1489 ( .A(n_445), .Y(n_1489) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .C(n_456), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g1092 ( .A(n_451), .Y(n_1092) );
INVx1_ASAP7_75t_L g1558 ( .A(n_451), .Y(n_1558) );
BUFx3_ASAP7_75t_L g589 ( .A(n_453), .Y(n_589) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g590 ( .A(n_455), .Y(n_590) );
INVx1_ASAP7_75t_L g942 ( .A(n_455), .Y(n_942) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_456), .B(n_483), .C(n_486), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g1037 ( .A(n_456), .B(n_1038), .C(n_1039), .Y(n_1037) );
AOI33xp33_ASAP7_75t_L g1090 ( .A1(n_456), .A2(n_683), .A3(n_1091), .B1(n_1093), .B2(n_1095), .B3(n_1097), .Y(n_1090) );
NAND3xp33_ASAP7_75t_L g1157 ( .A(n_456), .B(n_1158), .C(n_1160), .Y(n_1157) );
NAND3xp33_ASAP7_75t_L g1194 ( .A(n_456), .B(n_1195), .C(n_1196), .Y(n_1194) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g582 ( .A(n_459), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .C(n_465), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g484 ( .A(n_463), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_465), .B(n_490), .C(n_493), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g1040 ( .A(n_465), .B(n_1041), .C(n_1044), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_465), .B(n_1163), .C(n_1164), .Y(n_1162) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_465), .B(n_1200), .C(n_1201), .Y(n_1199) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_467), .B(n_1439), .Y(n_1438) );
XOR2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_519), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_498), .C(n_508), .Y(n_469) );
AND4x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_477), .C(n_482), .D(n_489), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .C(n_481), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_481), .A2(n_778), .B1(n_785), .B2(n_786), .C(n_792), .Y(n_777) );
INVx1_ASAP7_75t_L g991 ( .A(n_481), .Y(n_991) );
AOI33xp33_ASAP7_75t_L g1544 ( .A1(n_481), .A2(n_1545), .A3(n_1546), .B1(n_1550), .B2(n_1551), .B3(n_1552), .Y(n_1544) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_485), .Y(n_1022) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_488), .B(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g834 ( .A(n_491), .Y(n_834) );
BUFx3_ASAP7_75t_L g937 ( .A(n_491), .Y(n_937) );
INVx2_ASAP7_75t_L g1557 ( .A(n_491), .Y(n_1557) );
INVx1_ASAP7_75t_L g830 ( .A(n_492), .Y(n_830) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g542 ( .A(n_495), .Y(n_542) );
INVx2_ASAP7_75t_SL g573 ( .A(n_495), .Y(n_573) );
INVx2_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
INVx2_ASAP7_75t_L g744 ( .A(n_495), .Y(n_744) );
BUFx6f_ASAP7_75t_L g1043 ( .A(n_495), .Y(n_1043) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g1096 ( .A(n_497), .Y(n_1096) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x6_ASAP7_75t_L g644 ( .A(n_503), .B(n_627), .Y(n_644) );
INVx2_ASAP7_75t_L g1066 ( .A(n_513), .Y(n_1066) );
OAI22xp33_ASAP7_75t_L g1255 ( .A1(n_519), .A2(n_1224), .B1(n_1231), .B2(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g685 ( .A(n_520), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_595), .Y(n_520) );
INVx1_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_526), .A2(n_537), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_526), .A2(n_703), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_526), .A2(n_703), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1540 ( .A1(n_526), .A2(n_703), .B1(n_1541), .B2(n_1542), .Y(n_1540) );
AOI222xp33_ASAP7_75t_L g1080 ( .A1(n_532), .A2(n_699), .B1(n_1081), .B2(n_1082), .C1(n_1085), .C2(n_1086), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_535), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_535), .A2(n_537), .B1(n_799), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_535), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_535), .A2(n_537), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_535), .A2(n_537), .B1(n_1074), .B2(n_1088), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_535), .A2(n_902), .B1(n_1128), .B2(n_1145), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_535), .A2(n_902), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_548), .Y(n_610) );
INVx1_ASAP7_75t_L g718 ( .A(n_548), .Y(n_718) );
OAI31xp33_ASAP7_75t_SL g878 ( .A1(n_548), .A2(n_879), .A3(n_880), .B(n_881), .Y(n_878) );
OAI21xp5_ASAP7_75t_L g1524 ( .A1(n_548), .A2(n_1525), .B(n_1534), .Y(n_1524) );
NAND4xp25_ASAP7_75t_SL g549 ( .A(n_550), .B(n_560), .C(n_569), .D(n_583), .Y(n_549) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g729 ( .A(n_556), .Y(n_729) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g568 ( .A(n_557), .Y(n_568) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_557), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g740 ( .A(n_559), .Y(n_740) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g1109 ( .A(n_564), .Y(n_1109) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g620 ( .A(n_565), .Y(n_620) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_568), .B(n_652), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_576), .C(n_580), .Y(n_569) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g749 ( .A(n_579), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g671 ( .A(n_581), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_581), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_581), .A2(n_753), .B1(n_815), .B2(n_827), .Y(n_814) );
OAI22xp5_ASAP7_75t_SL g930 ( .A1(n_581), .A2(n_753), .B1(n_931), .B2(n_935), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_581), .A2(n_682), .B1(n_958), .B2(n_964), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .C(n_591), .Y(n_583) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx4f_ASAP7_75t_L g683 ( .A(n_592), .Y(n_683) );
INVx4_ASAP7_75t_L g753 ( .A(n_592), .Y(n_753) );
AOI221x1_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_610), .B1(n_611), .B2(n_653), .C(n_656), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .C(n_605), .D(n_609), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_603), .A2(n_646), .B1(n_647), .B2(n_648), .C1(n_649), .C2(n_650), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_606), .A2(n_639), .B(n_640), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_609), .B(n_706), .C(n_709), .D(n_711), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g1017 ( .A(n_609), .B(n_1018), .C(n_1021), .D(n_1024), .Y(n_1017) );
INVx1_ASAP7_75t_L g910 ( .A(n_610), .Y(n_910) );
OAI31xp33_ASAP7_75t_L g1053 ( .A1(n_610), .A2(n_1054), .A3(n_1055), .B(n_1059), .Y(n_1053) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_621), .C(n_645), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_616), .B2(n_617), .Y(n_612) );
INVx3_ASAP7_75t_L g1471 ( .A(n_614), .Y(n_1471) );
INVx2_ASAP7_75t_L g619 ( .A(n_615), .Y(n_619) );
INVx3_ASAP7_75t_L g1472 ( .A(n_617), .Y(n_1472) );
AND2x4_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g1102 ( .A(n_620), .Y(n_1102) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_637), .C(n_643), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x6_ASAP7_75t_L g630 ( .A(n_627), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g652 ( .A(n_627), .Y(n_652) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
CKINVDCx11_ASAP7_75t_R g1495 ( .A(n_630), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_636), .Y(n_632) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_635), .A2(n_658), .B1(n_660), .B2(n_662), .C(n_663), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_639), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
OAI22xp33_ASAP7_75t_SL g787 ( .A1(n_639), .A2(n_788), .B1(n_789), .B2(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g855 ( .A(n_639), .Y(n_855) );
BUFx2_ASAP7_75t_L g951 ( .A(n_639), .Y(n_951) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g672 ( .A1(n_646), .A2(n_648), .B1(n_673), .B2(n_676), .C(n_679), .Y(n_672) );
INVx8_ASAP7_75t_L g1483 ( .A(n_647), .Y(n_1483) );
CKINVDCx6p67_ASAP7_75t_R g1474 ( .A(n_649), .Y(n_1474) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g1441 ( .A(n_651), .B(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_652), .B(n_1493), .Y(n_1492) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
CKINVDCx8_ASAP7_75t_R g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_670), .B1(n_672), .B2(n_682), .Y(n_656) );
BUFx2_ASAP7_75t_L g828 ( .A(n_658), .Y(n_828) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx3_ASAP7_75t_L g796 ( .A(n_660), .Y(n_796) );
INVx1_ASAP7_75t_L g883 ( .A(n_660), .Y(n_883) );
OR2x6_ASAP7_75t_L g1503 ( .A(n_660), .B(n_1501), .Y(n_1503) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g678 ( .A(n_661), .Y(n_678) );
INVx1_ASAP7_75t_L g820 ( .A(n_661), .Y(n_820) );
INVx1_ASAP7_75t_L g1057 ( .A(n_661), .Y(n_1057) );
BUFx4f_ASAP7_75t_L g1452 ( .A(n_661), .Y(n_1452) );
BUFx4f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g1508 ( .A(n_665), .Y(n_1508) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g1094 ( .A(n_667), .Y(n_1094) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g969 ( .A(n_668), .Y(n_969) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI33xp33_ASAP7_75t_L g1554 ( .A1(n_671), .A2(n_683), .A3(n_1555), .B1(n_1559), .B2(n_1561), .B3(n_1563), .Y(n_1554) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g795 ( .A(n_675), .Y(n_795) );
INVx2_ASAP7_75t_L g932 ( .A(n_675), .Y(n_932) );
INVx1_ASAP7_75t_L g1506 ( .A(n_675), .Y(n_1506) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_682), .A2(n_793), .B1(n_1449), .B2(n_1455), .Y(n_1448) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
XNOR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_763), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx4f_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_732), .C(n_741), .D(n_751), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_728), .C(n_730), .Y(n_720) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx3_ASAP7_75t_L g913 ( .A(n_727), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_730), .A2(n_912), .B1(n_920), .B2(n_929), .C(n_930), .Y(n_911) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_734), .Y(n_914) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
BUFx3_ASAP7_75t_L g780 ( .A(n_737), .Y(n_780) );
INVx4_ASAP7_75t_L g1486 ( .A(n_737), .Y(n_1486) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .C(n_750), .Y(n_741) );
BUFx3_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_744), .Y(n_940) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g824 ( .A(n_748), .Y(n_824) );
BUFx3_ASAP7_75t_L g934 ( .A(n_748), .Y(n_934) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .C(n_759), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI22xp5_ASAP7_75t_SL g792 ( .A1(n_753), .A2(n_793), .B1(n_794), .B2(n_798), .Y(n_792) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
XNOR2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
NAND3x1_ASAP7_75t_SL g765 ( .A(n_766), .B(n_777), .C(n_802), .Y(n_765) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g926 ( .A(n_780), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g794 ( .A1(n_782), .A2(n_784), .B1(n_795), .B2(n_796), .C(n_797), .Y(n_794) );
OAI22xp5_ASAP7_75t_SL g915 ( .A1(n_789), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_915) );
INVx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g798 ( .A1(n_795), .A2(n_796), .B1(n_799), .B2(n_800), .C(n_801), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_795), .A2(n_882), .B1(n_959), .B2(n_960), .C(n_961), .Y(n_958) );
OAI221xp5_ASAP7_75t_L g931 ( .A1(n_796), .A2(n_916), .B1(n_917), .B2(n_932), .C(n_933), .Y(n_931) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_796), .A2(n_897), .B1(n_936), .B2(n_938), .C(n_939), .Y(n_935) );
BUFx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g885 ( .A(n_810), .Y(n_885) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_868), .C(n_878), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_837), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_818), .B2(n_821), .C(n_822), .Y(n_815) );
OAI22xp33_ASAP7_75t_L g851 ( .A1(n_816), .A2(n_821), .B1(n_852), .B2(n_854), .Y(n_851) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_817), .A2(n_965), .B1(n_966), .B2(n_967), .C(n_968), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g1449 ( .A1(n_817), .A2(n_1450), .B1(n_1451), .B2(n_1453), .C(n_1454), .Y(n_1449) );
OAI221xp5_ASAP7_75t_L g1455 ( .A1(n_817), .A2(n_966), .B1(n_1456), .B2(n_1457), .C(n_1458), .Y(n_1455) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx2_ASAP7_75t_L g966 ( .A(n_820), .Y(n_966) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B1(n_830), .B2(n_831), .C(n_832), .Y(n_827) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g1445 ( .A(n_836), .Y(n_1445) );
OAI33xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_842), .A3(n_851), .B1(n_856), .B2(n_862), .B3(n_867), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI33xp33_ASAP7_75t_L g970 ( .A1(n_840), .A2(n_971), .A3(n_974), .B1(n_980), .B2(n_985), .B3(n_991), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_847), .B2(n_850), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g1484 ( .A1(n_844), .A2(n_1485), .B1(n_1486), .B2(n_1487), .C(n_1488), .Y(n_1484) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_SL g976 ( .A(n_845), .Y(n_976) );
INVx2_ASAP7_75t_L g982 ( .A(n_845), .Y(n_982) );
BUFx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_852), .A2(n_857), .B1(n_858), .B2(n_861), .Y(n_856) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g1050 ( .A(n_855), .Y(n_1050) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_864), .B1(n_865), .B2(n_866), .Y(n_862) );
INVx1_ASAP7_75t_L g929 ( .A(n_867), .Y(n_929) );
BUFx3_ASAP7_75t_L g928 ( .A(n_871), .Y(n_928) );
BUFx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g919 ( .A(n_872), .Y(n_919) );
BUFx3_ASAP7_75t_L g1480 ( .A(n_872), .Y(n_1480) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_944), .B2(n_945), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_911), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_907), .B(n_910), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI22xp33_ASAP7_75t_SL g924 ( .A1(n_925), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g997 ( .A(n_947), .Y(n_997) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_956), .C(n_992), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_970), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_959), .A2(n_960), .B1(n_972), .B2(n_973), .Y(n_971) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_974) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI22xp5_ASAP7_75t_SL g980 ( .A1(n_981), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_982), .A2(n_1476), .B1(n_1477), .B2(n_1478), .Y(n_1475) );
OAI22xp33_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_988), .B1(n_989), .B2(n_990), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1223 ( .A1(n_998), .A2(n_1224), .B1(n_1229), .B2(n_1230), .Y(n_1223) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1118), .B1(n_1205), .B2(n_1206), .Y(n_1001) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1002), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1060), .B1(n_1116), .B2(n_1117), .Y(n_1003) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1004), .Y(n_1116) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1007), .Y(n_1052) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1014), .Y(n_1048) );
INVxp67_ASAP7_75t_L g1054 ( .A(n_1018), .Y(n_1054) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_1024), .Y(n_1059) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_1027), .B(n_1047), .C(n_1053), .Y(n_1046) );
AND4x1_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1033), .C(n_1037), .D(n_1040), .Y(n_1027) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
NAND3xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1035), .C(n_1036), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g1191 ( .A(n_1036), .B(n_1192), .C(n_1193), .Y(n_1191) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1043), .Y(n_1159) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1043), .Y(n_1560) );
INVx4_ASAP7_75t_L g1562 ( .A(n_1043), .Y(n_1562) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1057), .Y(n_1068) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1060), .Y(n_1117) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
NAND3xp33_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1070), .C(n_1073), .Y(n_1063) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1099), .Y(n_1089) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1102), .Y(n_1153) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1112), .Y(n_1156) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1112), .Y(n_1548) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1114), .Y(n_1549) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1118), .Y(n_1205) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_1121), .A2(n_1165), .B1(n_1166), .B2(n_1204), .Y(n_1120) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1121), .Y(n_1204) );
NAND3xp33_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1141), .C(n_1144), .Y(n_1134) );
NAND4xp25_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1151), .C(n_1157), .D(n_1162), .Y(n_1146) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1167), .Y(n_1203) );
NAND3xp33_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1182), .C(n_1184), .Y(n_1179) );
NAND4xp25_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1191), .C(n_1194), .D(n_1199), .Y(n_1187) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
OAI22xp33_ASAP7_75t_L g1307 ( .A1(n_1202), .A2(n_1308), .B1(n_1309), .B2(n_1310), .Y(n_1307) );
OAI221xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1428), .B1(n_1430), .B2(n_1509), .C(n_1515), .Y(n_1207) );
AND4x1_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1341), .C(n_1376), .D(n_1406), .Y(n_1208) );
A2O1A1Ixp33_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1294), .B(n_1295), .C(n_1325), .Y(n_1209) );
OAI211xp5_ASAP7_75t_SL g1210 ( .A1(n_1211), .A2(n_1243), .B(n_1273), .C(n_1276), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1233), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1212), .B(n_1291), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1212), .B(n_1234), .Y(n_1322) );
AND2x4_ASAP7_75t_SL g1417 ( .A(n_1212), .B(n_1233), .Y(n_1417) );
INVx2_ASAP7_75t_SL g1212 ( .A(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1213), .B(n_1233), .Y(n_1289) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1213), .Y(n_1294) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1214), .Y(n_1306) );
BUFx3_ASAP7_75t_L g1429 ( .A(n_1214), .Y(n_1429) );
AND2x4_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1218), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1215), .B(n_1218), .Y(n_1236) );
HB1xp67_ASAP7_75t_L g1568 ( .A(n_1215), .Y(n_1568) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
AND2x4_ASAP7_75t_L g1222 ( .A(n_1216), .B(n_1218), .Y(n_1222) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1217), .B(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1219), .Y(n_1228) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_1224), .A2(n_1231), .B1(n_1260), .B2(n_1261), .Y(n_1259) );
BUFx3_ASAP7_75t_L g1309 ( .A(n_1224), .Y(n_1309) );
BUFx6f_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1226), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1226), .Y(n_1240) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1227), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1567 ( .A(n_1228), .Y(n_1567) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1231), .Y(n_1311) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1232), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1233), .B(n_1268), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1233), .B(n_1292), .Y(n_1330) );
OAI221xp5_ASAP7_75t_L g1377 ( .A1(n_1233), .A2(n_1359), .B1(n_1378), .B2(n_1380), .C(n_1382), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1233), .B(n_1343), .Y(n_1385) );
CKINVDCx6p67_ASAP7_75t_R g1233 ( .A(n_1234), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1234), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1234), .B(n_1268), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1234), .B(n_1347), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1393 ( .A1(n_1234), .A2(n_1274), .B1(n_1394), .B2(n_1397), .C(n_1399), .Y(n_1393) );
A2O1A1Ixp33_ASAP7_75t_L g1407 ( .A1(n_1234), .A2(n_1361), .B(n_1408), .C(n_1409), .Y(n_1407) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_1234), .A2(n_1301), .B1(n_1353), .B2(n_1410), .C(n_1411), .Y(n_1409) );
OR2x6_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1237), .Y(n_1234) );
AND2x4_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1240), .Y(n_1238) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1240), .B(n_1242), .Y(n_1241) );
AOI211xp5_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1252), .B(n_1262), .C(n_1266), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1244), .B(n_1320), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1244), .B(n_1264), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1244), .B(n_1253), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1248), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1245), .B(n_1264), .Y(n_1263) );
INVx4_ASAP7_75t_L g1271 ( .A(n_1245), .Y(n_1271) );
INVx3_ASAP7_75t_L g1284 ( .A(n_1245), .Y(n_1284) );
NOR2xp67_ASAP7_75t_SL g1335 ( .A(n_1245), .B(n_1336), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_1245), .B(n_1370), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1245), .B(n_1253), .Y(n_1391) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1245), .B(n_1268), .Y(n_1419) );
AND2x4_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1248), .B(n_1275), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1248), .B(n_1286), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1248), .B(n_1257), .Y(n_1336) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1248), .B(n_1257), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1390 ( .A(n_1248), .B(n_1391), .Y(n_1390) );
BUFx3_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1249), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1249), .B(n_1286), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1249), .B(n_1264), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1249), .B(n_1253), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1249), .B(n_1320), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_1249), .B(n_1374), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1251), .Y(n_1249) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_1252), .A2(n_1339), .B(n_1340), .Y(n_1338) );
AOI21xp5_ASAP7_75t_L g1404 ( .A1(n_1252), .A2(n_1340), .B(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1253), .B(n_1299), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1253), .B(n_1284), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1257), .Y(n_1253) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1254), .Y(n_1265) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1254), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1254), .B(n_1258), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1257), .B(n_1265), .Y(n_1272) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1257), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1257), .B(n_1300), .Y(n_1403) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1258), .B(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1264), .B(n_1271), .Y(n_1275) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1264), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1264), .B(n_1299), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1272), .Y(n_1266) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1267), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1271), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g1292 ( .A(n_1268), .Y(n_1292) );
INVx1_ASAP7_75t_SL g1302 ( .A(n_1268), .Y(n_1302) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1268), .Y(n_1337) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1268), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1271), .B(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1271), .B(n_1300), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1271), .B(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1271), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1271), .B(n_1354), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1271), .B(n_1301), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1271), .B(n_1314), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1272), .B(n_1300), .Y(n_1360) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1272), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1272), .B(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_1275), .A2(n_1279), .B1(n_1328), .B2(n_1330), .C(n_1331), .Y(n_1327) );
A2O1A1Ixp33_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1280), .B(n_1281), .C(n_1287), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1279), .B(n_1319), .Y(n_1332) );
A2O1A1Ixp33_ASAP7_75t_L g1400 ( .A1(n_1279), .A2(n_1303), .B(n_1401), .C(n_1404), .Y(n_1400) );
INVxp67_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1285), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1283), .B(n_1330), .Y(n_1340) );
A2O1A1Ixp33_ASAP7_75t_L g1421 ( .A1(n_1283), .A2(n_1422), .B(n_1423), .C(n_1424), .Y(n_1421) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1284), .B(n_1351), .Y(n_1350) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1284), .B(n_1360), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1284), .B(n_1344), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1284), .B(n_1403), .Y(n_1402) );
NOR2x1_ASAP7_75t_L g1329 ( .A(n_1286), .B(n_1300), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1286), .B(n_1300), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1290), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1293), .Y(n_1290) );
AOI321xp33_ASAP7_75t_L g1341 ( .A1(n_1291), .A2(n_1301), .A3(n_1342), .B1(n_1345), .B2(n_1348), .C(n_1358), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1291), .B(n_1362), .Y(n_1361) );
NOR2xp33_ASAP7_75t_L g1380 ( .A(n_1291), .B(n_1381), .Y(n_1380) );
INVx3_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1292), .B(n_1379), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1292), .B(n_1417), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1293), .B(n_1304), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1326 ( .A(n_1293), .B(n_1304), .Y(n_1326) );
AOI21xp5_ASAP7_75t_SL g1406 ( .A1(n_1293), .A2(n_1407), .B(n_1415), .Y(n_1406) );
NOR3xp33_ASAP7_75t_L g1418 ( .A(n_1293), .B(n_1419), .C(n_1420), .Y(n_1418) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1294), .B(n_1314), .Y(n_1313) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1294), .Y(n_1356) );
INVxp67_ASAP7_75t_SL g1295 ( .A(n_1296), .Y(n_1295) );
OAI211xp5_ASAP7_75t_L g1325 ( .A1(n_1296), .A2(n_1326), .B(n_1327), .C(n_1333), .Y(n_1325) );
AOI221xp5_ASAP7_75t_L g1296 ( .A1(n_1297), .A2(n_1312), .B1(n_1313), .B2(n_1315), .C(n_1316), .Y(n_1296) );
OAI21xp33_ASAP7_75t_SL g1297 ( .A1(n_1298), .A2(n_1301), .B(n_1303), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1300), .B(n_1320), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1300), .B(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1301), .Y(n_1387) );
A2O1A1Ixp33_ASAP7_75t_L g1348 ( .A1(n_1303), .A2(n_1349), .B(n_1352), .C(n_1355), .Y(n_1348) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1303), .Y(n_1371) );
BUFx3_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1304), .Y(n_1347) );
AOI21xp5_ASAP7_75t_L g1363 ( .A1(n_1304), .A2(n_1364), .B(n_1365), .Y(n_1363) );
AOI31xp33_ASAP7_75t_L g1415 ( .A1(n_1304), .A2(n_1416), .A3(n_1421), .B(n_1425), .Y(n_1415) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1312), .Y(n_1388) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1313), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1313), .B(n_1324), .Y(n_1399) );
AOI21xp33_ASAP7_75t_L g1368 ( .A1(n_1314), .A2(n_1369), .B(n_1371), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1315), .B(n_1414), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_1317), .A2(n_1318), .B1(n_1321), .B2(n_1323), .Y(n_1316) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1317), .Y(n_1424) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1320), .Y(n_1370) );
NAND2xp5_ASAP7_75t_SL g1397 ( .A(n_1321), .B(n_1398), .Y(n_1397) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1416 ( .A1(n_1322), .A2(n_1334), .B1(n_1335), .B2(n_1417), .C(n_1418), .Y(n_1416) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
OAI21xp5_ASAP7_75t_L g1367 ( .A1(n_1328), .A2(n_1330), .B(n_1335), .Y(n_1367) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1329), .Y(n_1351) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
O2A1O1Ixp33_ASAP7_75t_L g1333 ( .A1(n_1334), .A2(n_1335), .B(n_1337), .C(n_1338), .Y(n_1333) );
NAND2xp5_ASAP7_75t_SL g1383 ( .A(n_1336), .B(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1337), .Y(n_1398) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1339), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1344), .Y(n_1342) );
AOI331xp33_ASAP7_75t_L g1358 ( .A1(n_1345), .A2(n_1359), .A3(n_1361), .B1(n_1363), .B2(n_1367), .B3(n_1368), .C1(n_1372), .Y(n_1358) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVxp67_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1354), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1357), .Y(n_1355) );
NOR2xp33_ASAP7_75t_L g1386 ( .A(n_1360), .B(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1375), .Y(n_1373) );
AOI21xp5_ASAP7_75t_L g1376 ( .A1(n_1377), .A2(n_1388), .B(n_1389), .Y(n_1376) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1379), .Y(n_1408) );
AOI21xp5_ASAP7_75t_SL g1382 ( .A1(n_1383), .A2(n_1385), .B(n_1386), .Y(n_1382) );
OAI21xp33_ASAP7_75t_L g1411 ( .A1(n_1384), .A2(n_1412), .B(n_1413), .Y(n_1411) );
OAI211xp5_ASAP7_75t_SL g1389 ( .A1(n_1390), .A2(n_1392), .B(n_1393), .C(n_1400), .Y(n_1389) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1390), .Y(n_1410) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1405), .Y(n_1423) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
CKINVDCx5p33_ASAP7_75t_R g1428 ( .A(n_1429), .Y(n_1428) );
HB1xp67_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
AND4x1_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1443), .C(n_1469), .D(n_1498), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1435), .Y(n_1433) );
OR2x6_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1441), .Y(n_1435) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
NOR3xp33_ASAP7_75t_SL g1443 ( .A(n_1444), .B(n_1448), .C(n_1459), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1446), .Y(n_1444) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVx2_ASAP7_75t_SL g1465 ( .A(n_1447), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1447), .B(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
OAI21xp33_ASAP7_75t_L g1479 ( .A1(n_1453), .A2(n_1480), .B(n_1481), .Y(n_1479) );
INVx2_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx2_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
NAND2x1p5_ASAP7_75t_L g1462 ( .A(n_1463), .B(n_1465), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
OAI31xp33_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1473), .A3(n_1482), .B(n_1496), .Y(n_1469) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1492), .B1(n_1494), .B2(n_1495), .Y(n_1490) );
BUFx8_ASAP7_75t_SL g1496 ( .A(n_1497), .Y(n_1496) );
NOR2xp33_ASAP7_75t_L g1498 ( .A(n_1499), .B(n_1504), .Y(n_1498) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1501), .B(n_1506), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1501), .B(n_1508), .Y(n_1507) );
CKINVDCx14_ASAP7_75t_R g1509 ( .A(n_1510), .Y(n_1509) );
INVx4_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
CKINVDCx5p33_ASAP7_75t_R g1517 ( .A(n_1518), .Y(n_1517) );
A2O1A1Ixp33_ASAP7_75t_L g1565 ( .A1(n_1519), .A2(n_1566), .B(n_1568), .C(n_1569), .Y(n_1565) );
INVxp33_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
HB1xp67_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
NAND4xp25_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1535), .C(n_1544), .D(n_1554), .Y(n_1523) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1531), .Y(n_1525) );
AO21x1_ASAP7_75t_SL g1535 ( .A1(n_1536), .A2(n_1540), .B(n_1543), .Y(n_1535) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
HB1xp67_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
endmodule