module fake_netlist_5_2389_n_1893 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1893);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1893;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1817;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_6),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_81),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_104),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_36),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_138),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_77),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_4),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_56),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_29),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_114),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_21),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_20),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_110),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_78),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_84),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_10),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_74),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_64),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_14),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_21),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_67),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_130),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_38),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_66),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_59),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_63),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_1),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_51),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_52),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_40),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_92),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_56),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_14),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_76),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_44),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_86),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_63),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_65),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_59),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_50),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_61),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_58),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_115),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_142),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_55),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_116),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_98),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_123),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_65),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_97),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_47),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_128),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_69),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_41),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_88),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_131),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_52),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_89),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_91),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_153),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_16),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_157),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_79),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_49),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_143),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_4),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_8),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_167),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_61),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_87),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_161),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_75),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_168),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_146),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_94),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_83),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_35),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_29),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_124),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_113),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_46),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_57),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_163),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_80),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_19),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_133),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_7),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_134),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_132),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_45),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_17),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_144),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_125),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_39),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_23),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_140),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_55),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_139),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_70),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_26),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_156),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_15),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_22),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_147),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_53),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_150),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_121),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_126),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_16),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_95),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_106),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_27),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_24),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_93),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_105),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_82),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_0),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_129),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_31),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_25),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_20),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_60),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_47),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_50),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_49),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_18),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_219),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_171),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_183),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_173),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_176),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_192),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_214),
.Y(n_348)
);

BUFx2_ASAP7_75t_SL g349 ( 
.A(n_223),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_214),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_214),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_214),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_180),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_266),
.B(n_220),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_266),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_172),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_179),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_281),
.B(n_0),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_281),
.B(n_2),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_220),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_220),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_234),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_233),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_233),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_181),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_233),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_249),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_237),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_237),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_182),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_237),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_2),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_244),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_184),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_312),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_186),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_265),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_244),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_262),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_244),
.B(n_3),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_196),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_274),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_274),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_199),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_177),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_274),
.B(n_5),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_200),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_203),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_197),
.B(n_262),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_180),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_205),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_193),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_193),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_282),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_194),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_198),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_187),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_282),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_180),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_198),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_202),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_213),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_202),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_265),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_215),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_208),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_208),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_225),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_217),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_405),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

BUFx8_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_210),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_363),
.B(n_358),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_407),
.A2(n_270),
.B1(n_339),
.B2(n_230),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_386),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_348),
.B(n_330),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_379),
.B(n_294),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_348),
.B(n_330),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_341),
.B(n_294),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_366),
.B(n_195),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_355),
.B(n_195),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_355),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_403),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_418),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_418),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_362),
.B(n_195),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_366),
.B(n_211),
.Y(n_463)
);

BUFx8_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_341),
.B(n_243),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_365),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_359),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_364),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_365),
.B(n_217),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_350),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_412),
.A2(n_310),
.B1(n_275),
.B2(n_221),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_417),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_350),
.B(n_211),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_421),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_375),
.B(n_211),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_359),
.B(n_375),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_351),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_369),
.Y(n_489)
);

CKINVDCx8_ASAP7_75t_R g490 ( 
.A(n_349),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_387),
.B(n_226),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_371),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_423),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_371),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_351),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_352),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_352),
.B(n_251),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_423),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_431),
.B(n_342),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_457),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_497),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_497),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_442),
.B(n_448),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_431),
.B(n_344),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_345),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

AOI22x1_ASAP7_75t_L g512 ( 
.A1(n_442),
.A2(n_406),
.B1(n_380),
.B2(n_373),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_346),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_498),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_432),
.Y(n_518)
);

CKINVDCx6p67_ASAP7_75t_R g519 ( 
.A(n_465),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_490),
.B(n_361),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_442),
.B(n_251),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_466),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_490),
.B(n_370),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_467),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_473),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_443),
.B(n_376),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g529 ( 
.A(n_465),
.B(n_389),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_473),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_490),
.B(n_382),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_470),
.B(n_353),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_457),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_470),
.B(n_385),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_448),
.B(n_387),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_487),
.B(n_390),
.Y(n_537)
);

NOR3xp33_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_395),
.C(n_389),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_467),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_470),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_473),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_473),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_470),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_464),
.B(n_393),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_426),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_487),
.B(n_396),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_457),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_429),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_464),
.B(n_398),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_474),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_464),
.B(n_400),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_445),
.B(n_404),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_464),
.B(n_416),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_474),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_461),
.B(n_349),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_448),
.B(n_422),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_463),
.B(n_401),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_428),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_463),
.B(n_353),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_461),
.A2(n_395),
.B1(n_356),
.B2(n_406),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_463),
.B(n_354),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_486),
.B(n_354),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_457),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_445),
.B(n_190),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_480),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_486),
.B(n_357),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_476),
.Y(n_576)
);

NOR2x1p5_ASAP7_75t_L g577 ( 
.A(n_475),
.B(n_272),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_457),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_464),
.B(n_419),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_480),
.Y(n_580)
);

AND2x2_ASAP7_75t_SL g581 ( 
.A(n_486),
.B(n_251),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_480),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_476),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_433),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_495),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_435),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_495),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_464),
.B(n_411),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_495),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_461),
.B(n_408),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_461),
.B(n_357),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_265),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_461),
.B(n_373),
.Y(n_593)
);

BUFx4f_ASAP7_75t_L g594 ( 
.A(n_476),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_461),
.B(n_441),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_435),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_434),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_495),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_383),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_441),
.B(n_391),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_437),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_475),
.B(n_380),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_476),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_441),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_437),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_440),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_440),
.Y(n_609)
);

INVxp33_ASAP7_75t_L g610 ( 
.A(n_430),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_498),
.B(n_265),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_430),
.Y(n_612)
);

BUFx4f_ASAP7_75t_L g613 ( 
.A(n_476),
.Y(n_613)
);

AOI21x1_ASAP7_75t_L g614 ( 
.A1(n_449),
.A2(n_356),
.B(n_402),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_441),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_462),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_441),
.B(n_391),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_462),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_469),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_469),
.B(n_343),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_444),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_468),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_478),
.B(n_383),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_428),
.B(n_243),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_471),
.B(n_347),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_444),
.B(n_394),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_476),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_SL g628 ( 
.A(n_434),
.B(n_372),
.C(n_367),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_L g629 ( 
.A(n_444),
.B(n_394),
.C(n_206),
.Y(n_629)
);

AO21x2_ASAP7_75t_L g630 ( 
.A1(n_484),
.A2(n_185),
.B(n_174),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_430),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_444),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_428),
.B(n_243),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_428),
.A2(n_384),
.B1(n_377),
.B2(n_333),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_468),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_L g637 ( 
.A(n_472),
.B(n_178),
.C(n_204),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_428),
.A2(n_229),
.B1(n_280),
.B2(n_240),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_428),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_472),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_444),
.B(n_212),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_468),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_444),
.B(n_477),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_479),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_479),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_476),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_R g648 ( 
.A(n_484),
.B(n_191),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_481),
.B(n_243),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_477),
.B(n_269),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_498),
.B(n_265),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_507),
.B(n_265),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_509),
.B(n_510),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_503),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_515),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_581),
.B(n_484),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_581),
.B(n_488),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_538),
.A2(n_484),
.B1(n_283),
.B2(n_498),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_621),
.B(n_488),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_537),
.B(n_484),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_650),
.A2(n_273),
.B1(n_247),
.B2(n_253),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_536),
.B(n_481),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_563),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_599),
.A2(n_273),
.B1(n_242),
.B2(n_247),
.Y(n_666)
);

A2O1A1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_529),
.A2(n_280),
.B(n_304),
.C(n_301),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_563),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_603),
.B(n_482),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_621),
.B(n_488),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_605),
.Y(n_671)
);

OAI221xp5_ASAP7_75t_L g672 ( 
.A1(n_567),
.A2(n_268),
.B1(n_229),
.B2(n_231),
.C(n_239),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_513),
.B(n_484),
.Y(n_673)
);

NOR2x1p5_ASAP7_75t_L g674 ( 
.A(n_519),
.B(n_209),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_605),
.B(n_482),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_595),
.B(n_488),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_503),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_638),
.A2(n_283),
.B1(n_185),
.B2(n_188),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_536),
.B(n_488),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_566),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_603),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_529),
.B(n_488),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_504),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_507),
.B(n_546),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_504),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_507),
.B(n_283),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_216),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_517),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_SL g689 ( 
.A1(n_597),
.A2(n_278),
.B1(n_340),
.B2(n_338),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_517),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_620),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_507),
.B(n_488),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_555),
.B(n_483),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_560),
.B(n_218),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_518),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_507),
.A2(n_590),
.B1(n_593),
.B2(n_522),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_625),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_526),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_566),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_507),
.B(n_488),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_607),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_561),
.B(n_222),
.Y(n_704)
);

BUFx8_ASAP7_75t_L g705 ( 
.A(n_522),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_525),
.B(n_224),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_518),
.B(n_483),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_565),
.B(n_496),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_521),
.B(n_524),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_519),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_518),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_568),
.B(n_496),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_539),
.B(n_626),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_SL g714 ( 
.A(n_539),
.B(n_325),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_522),
.A2(n_572),
.B1(n_599),
.B2(n_648),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_570),
.B(n_496),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_539),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_526),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_530),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_575),
.B(n_496),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_632),
.B(n_496),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_572),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_531),
.B(n_227),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_530),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_541),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_541),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_512),
.B(n_236),
.C(n_235),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_533),
.B(n_496),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_522),
.B(n_498),
.Y(n_729)
);

O2A1O1Ixp5_ASAP7_75t_L g730 ( 
.A1(n_632),
.A2(n_644),
.B(n_642),
.C(n_591),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_600),
.A2(n_438),
.B(n_427),
.Y(n_731)
);

NAND2x1_ASAP7_75t_L g732 ( 
.A(n_502),
.B(n_477),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_528),
.B(n_241),
.Y(n_733)
);

INVxp33_ASAP7_75t_L g734 ( 
.A(n_512),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_606),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_542),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_533),
.B(n_522),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_533),
.B(n_496),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_522),
.B(n_496),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_615),
.B(n_617),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_615),
.B(n_228),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_540),
.B(n_477),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_626),
.B(n_485),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_542),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_553),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_651),
.B(n_232),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_577),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_609),
.B(n_238),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_535),
.B(n_246),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_609),
.B(n_245),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_553),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_616),
.B(n_248),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_599),
.A2(n_284),
.B1(n_188),
.B2(n_329),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_626),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_599),
.A2(n_260),
.B1(n_332),
.B2(n_267),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_252),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_540),
.B(n_489),
.Y(n_757)
);

INVxp33_ASAP7_75t_L g758 ( 
.A(n_628),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_557),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_616),
.B(n_489),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_557),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_618),
.B(n_489),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_618),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_626),
.B(n_254),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_619),
.A2(n_286),
.B(n_231),
.C(n_239),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_619),
.B(n_489),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_558),
.A2(n_293),
.B1(n_329),
.B2(n_328),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_634),
.B(n_545),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_SL g769 ( 
.A1(n_597),
.A2(n_297),
.B1(n_337),
.B2(n_336),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_624),
.B(n_498),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_489),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_549),
.B(n_493),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_544),
.B(n_485),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_559),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_550),
.B(n_552),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_584),
.B(n_493),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_586),
.B(n_493),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_596),
.B(n_256),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_601),
.B(n_259),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_640),
.B(n_493),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_645),
.B(n_493),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_646),
.Y(n_782)
);

INVx8_ASAP7_75t_L g783 ( 
.A(n_558),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_633),
.B(n_602),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_612),
.B(n_491),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_500),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_505),
.B(n_276),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_514),
.B(n_498),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_543),
.B(n_498),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_602),
.B(n_174),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_630),
.A2(n_293),
.B1(n_207),
.B2(n_242),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_558),
.B(n_491),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_622),
.B(n_189),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_558),
.A2(n_284),
.B1(n_328),
.B2(n_207),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_622),
.B(n_189),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_610),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_636),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_636),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_551),
.B(n_264),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_641),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_630),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_L g802 ( 
.A(n_554),
.B(n_494),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_641),
.B(n_253),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_592),
.A2(n_499),
.B(n_494),
.C(n_286),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_643),
.B(n_649),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_623),
.A2(n_263),
.B1(n_279),
.B2(n_255),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_556),
.A2(n_305),
.B1(n_287),
.B2(n_288),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_643),
.B(n_255),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_649),
.B(n_257),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_635),
.B(n_271),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_623),
.B(n_499),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_630),
.B(n_257),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_534),
.B(n_258),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_520),
.B(n_298),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_614),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_559),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_562),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_520),
.B(n_299),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_614),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_562),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_534),
.B(n_578),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_576),
.A2(n_438),
.B(n_459),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_573),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_573),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_654),
.B(n_534),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_684),
.B(n_588),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_664),
.B(n_578),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_691),
.B(n_623),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_702),
.B(n_579),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_693),
.B(n_578),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_734),
.A2(n_564),
.B(n_639),
.C(n_637),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_655),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_653),
.A2(n_594),
.B(n_576),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_SL g834 ( 
.A(n_710),
.B(n_697),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_655),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_653),
.A2(n_662),
.B(n_673),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_677),
.Y(n_837)
);

BUFx12f_ASAP7_75t_L g838 ( 
.A(n_656),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_702),
.B(n_516),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_683),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_686),
.A2(n_679),
.B(n_740),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_696),
.B(n_520),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_672),
.A2(n_291),
.B(n_301),
.C(n_240),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_715),
.B(n_520),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_704),
.B(n_608),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_703),
.B(n_610),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_608),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_733),
.B(n_608),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_681),
.B(n_502),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_785),
.B(n_502),
.Y(n_850)
);

AOI21xp33_ASAP7_75t_L g851 ( 
.A1(n_687),
.A2(n_810),
.B(n_723),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_686),
.A2(n_594),
.B(n_576),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_659),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_665),
.B(n_520),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_740),
.A2(n_613),
.B(n_594),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_707),
.B(n_631),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_737),
.A2(n_613),
.B(n_571),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_669),
.B(n_631),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_657),
.B(n_547),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_665),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_658),
.A2(n_613),
.B(n_571),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_734),
.A2(n_709),
.B(n_799),
.C(n_667),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_717),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_665),
.A2(n_321),
.B1(n_258),
.B2(n_263),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_811),
.B(n_285),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_749),
.B(n_647),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_668),
.A2(n_647),
.B1(n_309),
.B2(n_317),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_675),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_675),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_730),
.A2(n_580),
.B(n_574),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_680),
.B(n_647),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_671),
.A2(n_303),
.B1(n_311),
.B2(n_314),
.Y(n_872)
);

CKINVDCx10_ASAP7_75t_R g873 ( 
.A(n_689),
.Y(n_873)
);

AND2x2_ASAP7_75t_SL g874 ( 
.A(n_784),
.B(n_277),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_796),
.B(n_289),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_783),
.B(n_547),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_658),
.A2(n_571),
.B(n_569),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_801),
.B(n_547),
.Y(n_878)
);

OAI21xp33_ASAP7_75t_L g879 ( 
.A1(n_714),
.A2(n_292),
.B(n_290),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_699),
.B(n_700),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_683),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_678),
.A2(n_652),
.B(n_611),
.C(n_592),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_692),
.A2(n_569),
.B(n_548),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_685),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_706),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_801),
.B(n_547),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_661),
.A2(n_589),
.B(n_582),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_815),
.A2(n_580),
.B(n_574),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_667),
.A2(n_652),
.B(n_611),
.C(n_321),
.Y(n_889)
);

OAI321xp33_ASAP7_75t_L g890 ( 
.A1(n_806),
.A2(n_304),
.A3(n_261),
.B1(n_268),
.B2(n_291),
.C(n_250),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_711),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_747),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_701),
.A2(n_569),
.B(n_548),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_783),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_783),
.B(n_277),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_754),
.B(n_279),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_L g897 ( 
.A(n_769),
.B(n_307),
.C(n_300),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_708),
.A2(n_547),
.B(n_548),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_712),
.A2(n_548),
.B(n_604),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_756),
.A2(n_758),
.B(n_764),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_716),
.A2(n_548),
.B(n_604),
.Y(n_901)
);

OAI321xp33_ASAP7_75t_L g902 ( 
.A1(n_663),
.A2(n_250),
.A3(n_261),
.B1(n_381),
.B2(n_378),
.C(n_374),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_754),
.B(n_374),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_720),
.A2(n_627),
.B(n_604),
.Y(n_904)
);

BUFx12f_ASAP7_75t_L g905 ( 
.A(n_695),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_685),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_675),
.B(n_812),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_735),
.A2(n_763),
.B(n_819),
.C(n_722),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_688),
.Y(n_909)
);

AO21x1_ASAP7_75t_L g910 ( 
.A1(n_682),
.A2(n_589),
.B(n_582),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_812),
.B(n_583),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_728),
.A2(n_738),
.B(n_721),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_721),
.A2(n_627),
.B(n_604),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_768),
.B(n_585),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_753),
.A2(n_598),
.B(n_587),
.C(n_585),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_782),
.B(n_587),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_702),
.A2(n_320),
.B1(n_322),
.B2(n_324),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_778),
.B(n_295),
.C(n_302),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_688),
.Y(n_919)
);

AOI21xp33_ASAP7_75t_L g920 ( 
.A1(n_758),
.A2(n_308),
.B(n_313),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_775),
.B(n_598),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_690),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_739),
.A2(n_627),
.B(n_604),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_SL g924 ( 
.A(n_710),
.B(n_325),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_690),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_743),
.B(n_316),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_676),
.A2(n_627),
.B(n_583),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_713),
.B(n_323),
.C(n_327),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_786),
.B(n_506),
.Y(n_929)
);

O2A1O1Ixp5_ASAP7_75t_L g930 ( 
.A1(n_682),
.A2(n_506),
.B(n_508),
.C(n_523),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_676),
.A2(n_508),
.B(n_511),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_792),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_727),
.B(n_318),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_773),
.A2(n_399),
.B(n_397),
.C(n_378),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_698),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_812),
.B(n_511),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_661),
.A2(n_627),
.B(n_583),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_802),
.A2(n_523),
.B(n_449),
.C(n_381),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_748),
.B(n_750),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_805),
.A2(n_762),
.B(n_760),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_792),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_748),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_670),
.A2(n_583),
.B(n_438),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_779),
.B(n_583),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_670),
.A2(n_438),
.B(n_527),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_821),
.A2(n_757),
.B(n_742),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_792),
.B(n_516),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_805),
.A2(n_771),
.B(n_766),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_784),
.A2(n_438),
.B(n_527),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_797),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_746),
.B(n_425),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_798),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_698),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_729),
.A2(n_438),
.B(n_527),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_729),
.A2(n_438),
.B(n_527),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_746),
.B(n_425),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_732),
.A2(n_438),
.B(n_527),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_791),
.A2(n_306),
.B1(n_325),
.B2(n_334),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_765),
.A2(n_392),
.B(n_397),
.C(n_399),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_814),
.A2(n_438),
.B(n_532),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_814),
.A2(n_532),
.B(n_516),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_818),
.A2(n_532),
.B(n_516),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_787),
.A2(n_325),
.B1(n_532),
.B2(n_516),
.Y(n_963)
);

AO21x1_ASAP7_75t_L g964 ( 
.A1(n_767),
.A2(n_392),
.B(n_402),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_750),
.B(n_752),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_718),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_818),
.A2(n_532),
.B(n_425),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_787),
.A2(n_460),
.B1(n_424),
.B2(n_450),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_783),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_718),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_752),
.B(n_425),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_731),
.A2(n_427),
.B(n_459),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_788),
.A2(n_427),
.B(n_459),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_789),
.A2(n_427),
.B(n_459),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_772),
.A2(n_776),
.B(n_777),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_705),
.B(n_424),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_765),
.A2(n_331),
.B(n_335),
.C(n_450),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_800),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_719),
.Y(n_979)
);

CKINVDCx6p67_ASAP7_75t_R g980 ( 
.A(n_741),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_719),
.B(n_436),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_780),
.A2(n_436),
.B(n_458),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_781),
.A2(n_436),
.B(n_458),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_724),
.Y(n_984)
);

AOI22x1_ASAP7_75t_L g985 ( 
.A1(n_724),
.A2(n_436),
.B1(n_458),
.B2(n_456),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_666),
.A2(n_460),
.B(n_424),
.C(n_450),
.Y(n_986)
);

BUFx24_ASAP7_75t_L g987 ( 
.A(n_705),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_725),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_705),
.B(n_460),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_741),
.A2(n_458),
.B(n_456),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_SL g991 ( 
.A(n_794),
.B(n_306),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_790),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_755),
.A2(n_451),
.B1(n_455),
.B2(n_452),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_674),
.B(n_306),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_770),
.B(n_452),
.C(n_455),
.Y(n_995)
);

BUFx4f_ASAP7_75t_L g996 ( 
.A(n_820),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_660),
.A2(n_452),
.B1(n_455),
.B2(n_451),
.Y(n_997)
);

AND3x4_ASAP7_75t_L g998 ( 
.A(n_725),
.B(n_456),
.C(n_454),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_807),
.B(n_5),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_726),
.Y(n_1000)
);

AOI22x1_ASAP7_75t_SL g1001 ( 
.A1(n_823),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_726),
.B(n_456),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_770),
.A2(n_454),
.B(n_447),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_736),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_736),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_813),
.A2(n_454),
.B(n_447),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_744),
.B(n_454),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_744),
.B(n_447),
.Y(n_1008)
);

AOI21x1_ASAP7_75t_L g1009 ( 
.A1(n_822),
.A2(n_447),
.B(n_446),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_804),
.A2(n_453),
.B(n_451),
.C(n_446),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_745),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_824),
.B(n_453),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_745),
.A2(n_446),
.B(n_439),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_751),
.B(n_453),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_793),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_851),
.A2(n_795),
.B1(n_803),
.B2(n_808),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_999),
.A2(n_809),
.B1(n_824),
.B2(n_816),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_885),
.B(n_817),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_868),
.B(n_759),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_838),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_862),
.A2(n_817),
.B(n_816),
.C(n_774),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_868),
.B(n_761),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_860),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_999),
.A2(n_874),
.B1(n_900),
.B2(n_939),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_894),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_939),
.A2(n_965),
.B1(n_942),
.B2(n_907),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_853),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_856),
.B(n_761),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_862),
.A2(n_759),
.B(n_751),
.C(n_446),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_837),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_846),
.B(n_9),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_850),
.B(n_439),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_874),
.A2(n_439),
.B1(n_12),
.B2(n_13),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_858),
.B(n_11),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_909),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_965),
.B(n_439),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_894),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_SL g1038 ( 
.A1(n_826),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_1038)
);

OA22x2_ASAP7_75t_L g1039 ( 
.A1(n_828),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_833),
.A2(n_836),
.B(n_852),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_894),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_869),
.B(n_159),
.Y(n_1042)
);

AND2x2_ASAP7_75t_SL g1043 ( 
.A(n_876),
.B(n_158),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_850),
.B(n_24),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_909),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_853),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_920),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_869),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_926),
.B(n_28),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_941),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_966),
.Y(n_1051)
);

BUFx10_ASAP7_75t_L g1052 ( 
.A(n_926),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_859),
.A2(n_845),
.B(n_907),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_992),
.B(n_30),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_834),
.B(n_905),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_992),
.B(n_30),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_881),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_825),
.A2(n_68),
.B1(n_152),
.B2(n_151),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_932),
.B(n_155),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1015),
.B(n_31),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_1004),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_987),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_908),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_941),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_875),
.B(n_33),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_944),
.A2(n_148),
.B(n_145),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_922),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_892),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_SL g1069 ( 
.A1(n_826),
.A2(n_34),
.B(n_37),
.C(n_38),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_894),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_932),
.B(n_71),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_R g1072 ( 
.A(n_969),
.B(n_43),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_936),
.A2(n_141),
.B(n_122),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_980),
.B(n_101),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_880),
.B(n_43),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_966),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_865),
.B(n_44),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_849),
.B(n_45),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_847),
.A2(n_118),
.B(n_117),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_1004),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_911),
.A2(n_112),
.B1(n_108),
.B2(n_100),
.Y(n_1081)
);

AOI22x1_ASAP7_75t_L g1082 ( 
.A1(n_855),
.A2(n_99),
.B1(n_72),
.B2(n_53),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_933),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_841),
.A2(n_62),
.B(n_48),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_863),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_911),
.A2(n_46),
.B1(n_48),
.B2(n_54),
.Y(n_1086)
);

BUFx2_ASAP7_75t_SL g1087 ( 
.A(n_891),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_979),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_883),
.A2(n_893),
.B(n_866),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_848),
.A2(n_57),
.B(n_58),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_849),
.B(n_60),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_857),
.A2(n_62),
.B(n_861),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_979),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_998),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_903),
.B(n_827),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_903),
.B(n_921),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_908),
.A2(n_842),
.B1(n_829),
.B2(n_844),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_925),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_996),
.B(n_1004),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_896),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_928),
.A2(n_933),
.B1(n_918),
.B2(n_947),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_831),
.A2(n_977),
.B(n_843),
.C(n_897),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_947),
.B(n_996),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_877),
.A2(n_844),
.B(n_842),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_898),
.A2(n_923),
.B(n_901),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_832),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_991),
.B(n_879),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_899),
.A2(n_912),
.B(n_888),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_904),
.A2(n_946),
.B(n_830),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_835),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_854),
.A2(n_914),
.B(n_975),
.Y(n_1111)
);

CKINVDCx11_ASAP7_75t_R g1112 ( 
.A(n_895),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_SL g1113 ( 
.A1(n_977),
.A2(n_843),
.B(n_878),
.C(n_886),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_854),
.A2(n_886),
.B(n_878),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_927),
.A2(n_913),
.B(n_951),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_840),
.B(n_884),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_956),
.A2(n_948),
.B(n_940),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_895),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_906),
.B(n_919),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_895),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_897),
.B(n_924),
.C(n_958),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_998),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_937),
.A2(n_971),
.B(n_870),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_829),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_839),
.A2(n_871),
.B(n_931),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_950),
.A2(n_978),
.B1(n_952),
.B2(n_916),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_839),
.A2(n_929),
.B(n_955),
.Y(n_1128)
);

NOR2xp67_ASAP7_75t_L g1129 ( 
.A(n_872),
.B(n_994),
.Y(n_1129)
);

AO21x1_ASAP7_75t_L g1130 ( 
.A1(n_976),
.A2(n_989),
.B(n_864),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_890),
.A2(n_928),
.B(n_934),
.C(n_989),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_934),
.A2(n_976),
.B(n_917),
.C(n_958),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_954),
.A2(n_1007),
.B(n_1002),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_935),
.B(n_953),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_970),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_984),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_988),
.A2(n_1011),
.B1(n_1000),
.B2(n_1005),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1012),
.B(n_1014),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1012),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_995),
.B(n_959),
.Y(n_1140)
);

CKINVDCx14_ASAP7_75t_R g1141 ( 
.A(n_873),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_887),
.Y(n_1142)
);

AO21x1_ASAP7_75t_L g1143 ( 
.A1(n_990),
.A2(n_995),
.B(n_915),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1014),
.Y(n_1144)
);

NAND2x1_ASAP7_75t_L g1145 ( 
.A(n_981),
.B(n_1008),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_867),
.A2(n_963),
.B1(n_964),
.B2(n_993),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_902),
.B(n_938),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_910),
.B(n_997),
.Y(n_1148)
);

OR2x6_ASAP7_75t_SL g1149 ( 
.A(n_1001),
.B(n_882),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1009),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_961),
.A2(n_962),
.B(n_967),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_930),
.A2(n_949),
.B(n_974),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1003),
.A2(n_973),
.B(n_1010),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_968),
.B(n_1010),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_972),
.B(n_943),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_959),
.B(n_889),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_960),
.A2(n_945),
.B(n_982),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_983),
.B(n_986),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_985),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1013),
.A2(n_654),
.B1(n_851),
.B2(n_862),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1006),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_957),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_SL g1163 ( 
.A1(n_833),
.A2(n_639),
.B(n_564),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_851),
.B(n_654),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_851),
.B(n_654),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_838),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_894),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_851),
.A2(n_654),
.B1(n_862),
.B2(n_907),
.Y(n_1168)
);

OAI21xp33_ASAP7_75t_L g1169 ( 
.A1(n_851),
.A2(n_654),
.B(n_509),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_838),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_838),
.Y(n_1171)
);

AO21x1_ASAP7_75t_L g1172 ( 
.A1(n_851),
.A2(n_654),
.B(n_826),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_894),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1030),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1085),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1057),
.Y(n_1176)
);

INVx5_ASAP7_75t_L g1177 ( 
.A(n_1025),
.Y(n_1177)
);

OA21x2_ASAP7_75t_L g1178 ( 
.A1(n_1117),
.A2(n_1040),
.B(n_1104),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1028),
.B(n_1165),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_1170),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1067),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1098),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1165),
.A2(n_1169),
.B(n_1107),
.C(n_1164),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1025),
.B(n_1037),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1164),
.B(n_1026),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1168),
.A2(n_1024),
.B(n_1107),
.C(n_1049),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1109),
.A2(n_1089),
.B(n_1108),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1024),
.B(n_1018),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1102),
.A2(n_1122),
.B(n_1132),
.C(n_1131),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1077),
.B(n_1065),
.C(n_1078),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1105),
.A2(n_1151),
.B(n_1152),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1068),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1027),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1046),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1018),
.B(n_1096),
.Y(n_1195)
);

AO32x2_ASAP7_75t_L g1196 ( 
.A1(n_1097),
.A2(n_1160),
.A3(n_1086),
.B1(n_1137),
.B2(n_1127),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1033),
.A2(n_1123),
.B1(n_1094),
.B2(n_1043),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1034),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1025),
.B(n_1037),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1101),
.A2(n_1091),
.B(n_1078),
.C(n_1077),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1106),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1172),
.A2(n_1143),
.A3(n_1092),
.B(n_1130),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1033),
.A2(n_1123),
.B1(n_1094),
.B2(n_1043),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_SL g1204 ( 
.A(n_1123),
.B(n_1062),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1053),
.A2(n_1111),
.B(n_1128),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1065),
.B(n_1091),
.C(n_1047),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1100),
.B(n_1050),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1052),
.B(n_1046),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1163),
.A2(n_1124),
.B(n_1133),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1158),
.A2(n_1115),
.A3(n_1016),
.B(n_1126),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1083),
.A2(n_1123),
.B1(n_1031),
.B2(n_1039),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1032),
.A2(n_1155),
.B(n_1153),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1155),
.A2(n_1157),
.B(n_1148),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_1112),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1021),
.A2(n_1029),
.B(n_1150),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1055),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_1084),
.A2(n_1044),
.B(n_1063),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1031),
.B(n_1064),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1154),
.A2(n_1114),
.B(n_1158),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1025),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1087),
.B(n_1103),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1145),
.A2(n_1036),
.B(n_1113),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1021),
.A2(n_1036),
.B(n_1147),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1142),
.A2(n_1162),
.A3(n_1090),
.B(n_1125),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_SL g1225 ( 
.A1(n_1075),
.A2(n_1140),
.B(n_1156),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1146),
.A2(n_1129),
.B(n_1095),
.C(n_1054),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1134),
.B(n_1139),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1110),
.B(n_1017),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1055),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1023),
.A2(n_1099),
.B(n_1017),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1144),
.B(n_1045),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1056),
.A2(n_1060),
.B(n_1058),
.C(n_1071),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1136),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1019),
.A2(n_1022),
.B(n_1042),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1150),
.A2(n_1019),
.B(n_1022),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1125),
.B(n_1048),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1066),
.A2(n_1079),
.A3(n_1138),
.B(n_1081),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1118),
.B(n_1121),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_SL g1240 ( 
.A1(n_1071),
.A2(n_1042),
.B(n_1059),
.C(n_1120),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1116),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1039),
.B(n_1035),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1171),
.Y(n_1243)
);

AOI221xp5_ASAP7_75t_L g1244 ( 
.A1(n_1074),
.A2(n_1073),
.B1(n_1020),
.B2(n_1166),
.C(n_1120),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1082),
.A2(n_1080),
.B(n_1119),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1103),
.B(n_1048),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1051),
.A2(n_1088),
.B(n_1076),
.C(n_1093),
.Y(n_1247)
);

BUFx2_ASAP7_75t_R g1248 ( 
.A(n_1061),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1038),
.A2(n_1069),
.B(n_1159),
.Y(n_1249)
);

NOR2xp67_ASAP7_75t_L g1250 ( 
.A(n_1161),
.B(n_1080),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1061),
.B(n_1119),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1135),
.A2(n_1037),
.B(n_1041),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1072),
.A2(n_1135),
.A3(n_1041),
.B(n_1070),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1135),
.A2(n_1037),
.B(n_1041),
.C(n_1070),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1173),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1135),
.B(n_1070),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1141),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1070),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1167),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1167),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1167),
.A2(n_1173),
.B(n_1074),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1167),
.A2(n_1040),
.B(n_1105),
.Y(n_1262)
);

OAI22x1_ASAP7_75t_L g1263 ( 
.A1(n_1173),
.A2(n_1165),
.B1(n_1122),
.B2(n_654),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1173),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1040),
.A2(n_1105),
.B(n_1109),
.Y(n_1265)
);

AOI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1036),
.A2(n_826),
.B(n_1126),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1030),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1097),
.A2(n_1172),
.A3(n_1143),
.B(n_1040),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1165),
.B(n_654),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1165),
.B(n_654),
.C(n_851),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1030),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1165),
.A2(n_654),
.B(n_851),
.C(n_1169),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1040),
.A2(n_1105),
.B(n_1109),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1055),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1165),
.A2(n_654),
.B(n_851),
.C(n_1169),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1030),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1030),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1030),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1281)
);

CKINVDCx9p33_ASAP7_75t_R g1282 ( 
.A(n_1170),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1097),
.A2(n_1172),
.A3(n_1143),
.B(n_1040),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1097),
.A2(n_1172),
.A3(n_1143),
.B(n_1040),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1030),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_SL g1287 ( 
.A(n_1043),
.B(n_654),
.Y(n_1287)
);

OAI22x1_ASAP7_75t_L g1288 ( 
.A1(n_1165),
.A2(n_1122),
.B1(n_654),
.B2(n_1164),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1040),
.A2(n_1108),
.B(n_1117),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1290)
);

BUFx10_ASAP7_75t_L g1291 ( 
.A(n_1031),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1165),
.A2(n_654),
.B1(n_851),
.B2(n_1169),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1169),
.A2(n_654),
.B(n_851),
.C(n_1165),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1165),
.B(n_654),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1164),
.B(n_858),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1165),
.B(n_654),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1165),
.A2(n_1168),
.B(n_654),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1040),
.A2(n_1105),
.B(n_1109),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_SL g1299 ( 
.A(n_1043),
.B(n_654),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1025),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1165),
.B(n_654),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1030),
.Y(n_1302)
);

AOI221x1_ASAP7_75t_L g1303 ( 
.A1(n_1165),
.A2(n_1169),
.B1(n_654),
.B2(n_851),
.C(n_1168),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1030),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1097),
.A2(n_1172),
.A3(n_1143),
.B(n_1040),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1165),
.B(n_654),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1165),
.A2(n_654),
.B1(n_1024),
.B2(n_1033),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1040),
.A2(n_1105),
.B(n_1109),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1165),
.A2(n_654),
.B(n_851),
.C(n_1169),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1165),
.B(n_654),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1030),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1165),
.A2(n_654),
.B(n_851),
.C(n_1169),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1040),
.A2(n_1105),
.B(n_1109),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1165),
.B(n_654),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1028),
.B(n_856),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1164),
.B(n_858),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1040),
.A2(n_1105),
.B(n_1109),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1097),
.A2(n_1172),
.A3(n_1143),
.B(n_1040),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1165),
.A2(n_654),
.B1(n_851),
.B2(n_1169),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1164),
.B(n_858),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1165),
.B(n_654),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_SL g1325 ( 
.A(n_1020),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1097),
.A2(n_1172),
.A3(n_1143),
.B(n_1040),
.Y(n_1326)
);

AOI211x1_ASAP7_75t_L g1327 ( 
.A1(n_1169),
.A2(n_851),
.B(n_806),
.C(n_1164),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1028),
.B(n_856),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1040),
.A2(n_836),
.B(n_654),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1117),
.A2(n_1040),
.B(n_1104),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1112),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1025),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1165),
.B(n_654),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1112),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1325),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1207),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1294),
.A2(n_1296),
.B1(n_1301),
.B2(n_1307),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1307),
.A2(n_1190),
.B1(n_1270),
.B2(n_1297),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1190),
.A2(n_1200),
.B1(n_1322),
.B2(n_1292),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1175),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1207),
.Y(n_1341)
);

INVx11_ASAP7_75t_L g1342 ( 
.A(n_1180),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1269),
.B(n_1311),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1270),
.A2(n_1315),
.B1(n_1333),
.B2(n_1306),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_L g1345 ( 
.A(n_1273),
.B(n_1276),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1306),
.A2(n_1206),
.B1(n_1310),
.B2(n_1313),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1287),
.A2(n_1299),
.B1(n_1324),
.B2(n_1206),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1297),
.A2(n_1288),
.B1(n_1299),
.B2(n_1287),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1211),
.A2(n_1197),
.B1(n_1203),
.B2(n_1188),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1197),
.A2(n_1203),
.B1(n_1183),
.B2(n_1295),
.Y(n_1350)
);

BUFx8_ASAP7_75t_SL g1351 ( 
.A(n_1257),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1300),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1179),
.A2(n_1185),
.B1(n_1291),
.B2(n_1263),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1291),
.A2(n_1217),
.B1(n_1317),
.B2(n_1323),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1239),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1303),
.A2(n_1195),
.B1(n_1198),
.B2(n_1236),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1277),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1177),
.Y(n_1358)
);

CKINVDCx11_ASAP7_75t_R g1359 ( 
.A(n_1214),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1180),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1233),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1293),
.B(n_1316),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1275),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1218),
.A2(n_1219),
.B1(n_1328),
.B2(n_1241),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1177),
.Y(n_1365)
);

INVx8_ASAP7_75t_L g1366 ( 
.A(n_1177),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1189),
.A2(n_1226),
.B1(n_1327),
.B2(n_1208),
.Y(n_1367)
);

BUFx8_ASAP7_75t_L g1368 ( 
.A(n_1325),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1244),
.A2(n_1286),
.B1(n_1242),
.B2(n_1201),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1174),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1223),
.A2(n_1334),
.B1(n_1331),
.B2(n_1186),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1228),
.A2(n_1227),
.B1(n_1312),
.B2(n_1181),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1216),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1258),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1192),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1176),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1227),
.B(n_1194),
.Y(n_1377)
);

INVxp33_ASAP7_75t_SL g1378 ( 
.A(n_1204),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1182),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1229),
.A2(n_1221),
.B1(n_1304),
.B2(n_1302),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1250),
.A2(n_1221),
.B1(n_1243),
.B2(n_1246),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1223),
.A2(n_1280),
.B1(n_1279),
.B2(n_1267),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1228),
.A2(n_1249),
.B1(n_1221),
.B2(n_1250),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1231),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1249),
.A2(n_1212),
.B1(n_1272),
.B2(n_1290),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_SL g1386 ( 
.A(n_1259),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1251),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1251),
.Y(n_1388)
);

BUFx2_ASAP7_75t_SL g1389 ( 
.A(n_1300),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1278),
.A2(n_1283),
.B1(n_1308),
.B2(n_1281),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1300),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1318),
.A2(n_1329),
.B1(n_1321),
.B2(n_1230),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1234),
.A2(n_1213),
.B1(n_1289),
.B2(n_1222),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1261),
.A2(n_1237),
.B1(n_1256),
.B2(n_1264),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1256),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1224),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1248),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1240),
.A2(n_1237),
.B1(n_1264),
.B2(n_1260),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1247),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1253),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1289),
.A2(n_1178),
.B1(n_1330),
.B2(n_1205),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1282),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1232),
.A2(n_1254),
.B1(n_1255),
.B2(n_1184),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1184),
.A2(n_1199),
.B1(n_1252),
.B2(n_1332),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1199),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1268),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1178),
.A2(n_1330),
.B1(n_1215),
.B2(n_1187),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1220),
.A2(n_1209),
.B1(n_1225),
.B2(n_1266),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1235),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1196),
.A2(n_1262),
.B1(n_1245),
.B2(n_1191),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1210),
.B(n_1285),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1268),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1196),
.A2(n_1285),
.B1(n_1320),
.B2(n_1305),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1202),
.A2(n_1238),
.B1(n_1326),
.B2(n_1320),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1268),
.B(n_1326),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1210),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_1238),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1202),
.A2(n_1238),
.B1(n_1326),
.B2(n_1320),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1210),
.B(n_1305),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1265),
.A2(n_1298),
.B(n_1274),
.Y(n_1420)
);

BUFx8_ASAP7_75t_L g1421 ( 
.A(n_1202),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1309),
.A2(n_1314),
.B1(n_1319),
.B2(n_1305),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1284),
.A2(n_1296),
.B1(n_1301),
.B2(n_1294),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1285),
.A2(n_654),
.B1(n_1165),
.B2(n_1296),
.Y(n_1424)
);

INVx6_ASAP7_75t_L g1425 ( 
.A(n_1177),
.Y(n_1425)
);

CKINVDCx6p67_ASAP7_75t_R g1426 ( 
.A(n_1282),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1294),
.A2(n_1301),
.B1(n_1296),
.B2(n_1307),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1177),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1175),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1294),
.A2(n_654),
.B(n_851),
.Y(n_1430)
);

BUFx8_ASAP7_75t_L g1431 ( 
.A(n_1325),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1175),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1207),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1307),
.A2(n_1269),
.B1(n_1315),
.B2(n_1311),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1180),
.Y(n_1435)
);

BUFx8_ASAP7_75t_SL g1436 ( 
.A(n_1257),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1177),
.B(n_1258),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1177),
.Y(n_1438)
);

BUFx5_ASAP7_75t_L g1439 ( 
.A(n_1241),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1294),
.A2(n_654),
.B1(n_1165),
.B2(n_1296),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1214),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1271),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1177),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1177),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1294),
.A2(n_1301),
.B1(n_1296),
.B2(n_1307),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1177),
.Y(n_1446)
);

BUFx8_ASAP7_75t_L g1447 ( 
.A(n_1325),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1207),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1193),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1177),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1193),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1294),
.A2(n_654),
.B1(n_1301),
.B2(n_1296),
.Y(n_1452)
);

OAI22x1_ASAP7_75t_L g1453 ( 
.A1(n_1190),
.A2(n_1165),
.B1(n_1296),
.B2(n_1294),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1175),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1257),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1294),
.A2(n_654),
.B1(n_1301),
.B2(n_1296),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1294),
.A2(n_654),
.B1(n_1301),
.B2(n_1296),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1294),
.A2(n_654),
.B1(n_1165),
.B2(n_1296),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1294),
.A2(n_1301),
.B1(n_1296),
.B2(n_1307),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1271),
.Y(n_1460)
);

OAI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1294),
.A2(n_654),
.B(n_1165),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1409),
.B(n_1400),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1338),
.B(n_1423),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1440),
.A2(n_1339),
.B1(n_1349),
.B2(n_1350),
.Y(n_1464)
);

OAI21xp33_ASAP7_75t_L g1465 ( 
.A1(n_1461),
.A2(n_1456),
.B(n_1452),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1366),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1415),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1337),
.A2(n_1427),
.B1(n_1445),
.B2(n_1459),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1338),
.B(n_1423),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1408),
.B(n_1417),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1345),
.A2(n_1346),
.B1(n_1367),
.B2(n_1424),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1377),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1401),
.A2(n_1407),
.B(n_1392),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1439),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1395),
.B(n_1348),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1348),
.B(n_1387),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1396),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1388),
.B(n_1376),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1449),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1430),
.A2(n_1452),
.B(n_1456),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1421),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1359),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1406),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1401),
.A2(n_1407),
.B(n_1392),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1390),
.A2(n_1410),
.B(n_1393),
.Y(n_1486)
);

BUFx2_ASAP7_75t_SL g1487 ( 
.A(n_1450),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1411),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1422),
.A2(n_1420),
.B(n_1413),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1413),
.A2(n_1419),
.B(n_1418),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1405),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1421),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1380),
.B(n_1414),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1453),
.B(n_1416),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1439),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1458),
.B(n_1457),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1370),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1379),
.B(n_1398),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1450),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1372),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1372),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1457),
.B(n_1343),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1405),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1384),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1444),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1460),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1357),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1366),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1450),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1362),
.B(n_1344),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1351),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1451),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1390),
.A2(n_1393),
.B(n_1385),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1434),
.B(n_1337),
.Y(n_1515)
);

AO31x2_ASAP7_75t_L g1516 ( 
.A1(n_1403),
.A2(n_1399),
.A3(n_1404),
.B(n_1410),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1385),
.A2(n_1382),
.B(n_1383),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1353),
.B(n_1364),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1354),
.A2(n_1383),
.B(n_1382),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1358),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1354),
.A2(n_1364),
.B(n_1369),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1366),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1369),
.A2(n_1437),
.B(n_1442),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1436),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1355),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1434),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1394),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1427),
.B(n_1459),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1361),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1394),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1445),
.B(n_1371),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1429),
.B(n_1378),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1356),
.B(n_1371),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1356),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1381),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1365),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1425),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1340),
.A2(n_1432),
.B1(n_1454),
.B2(n_1341),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1336),
.B(n_1448),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1433),
.A2(n_1402),
.B(n_1397),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1352),
.B(n_1391),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1443),
.A2(n_1446),
.B(n_1389),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1443),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1473),
.B(n_1373),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1529),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1468),
.B(n_1426),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1497),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1497),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1464),
.A2(n_1363),
.B(n_1360),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1468),
.B(n_1335),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1490),
.B(n_1428),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1464),
.A2(n_1455),
.B(n_1335),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1511),
.B(n_1447),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1514),
.A2(n_1438),
.B(n_1374),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1462),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1496),
.A2(n_1375),
.B1(n_1435),
.B2(n_1368),
.Y(n_1556)
);

NAND4xp25_ASAP7_75t_SL g1557 ( 
.A(n_1481),
.B(n_1447),
.C(n_1368),
.D(n_1431),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_SL g1558 ( 
.A1(n_1481),
.A2(n_1431),
.B(n_1342),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1490),
.B(n_1488),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1469),
.A2(n_1441),
.B1(n_1386),
.B2(n_1438),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1465),
.A2(n_1386),
.B(n_1515),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1465),
.A2(n_1472),
.B(n_1531),
.C(n_1503),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1539),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_SL g1564 ( 
.A1(n_1534),
.A2(n_1526),
.B(n_1532),
.C(n_1506),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1479),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1462),
.B(n_1492),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1534),
.A2(n_1485),
.B(n_1474),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1540),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_SL g1571 ( 
.A1(n_1533),
.A2(n_1515),
.B(n_1492),
.C(n_1535),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1486),
.A2(n_1474),
.B(n_1485),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1531),
.A2(n_1521),
.B(n_1533),
.C(n_1517),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_SL g1574 ( 
.A(n_1512),
.B(n_1524),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1463),
.B(n_1470),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1490),
.B(n_1488),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

AO32x2_ASAP7_75t_L g1578 ( 
.A1(n_1491),
.A2(n_1504),
.A3(n_1520),
.B1(n_1490),
.B2(n_1484),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1521),
.A2(n_1517),
.B(n_1528),
.C(n_1470),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1521),
.A2(n_1517),
.B(n_1528),
.C(n_1463),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1483),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1494),
.B(n_1526),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1480),
.B(n_1513),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1518),
.A2(n_1498),
.B(n_1527),
.C(n_1530),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1540),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1494),
.B(n_1493),
.Y(n_1586)
);

CKINVDCx8_ASAP7_75t_R g1587 ( 
.A(n_1487),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1493),
.B(n_1508),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1535),
.A2(n_1538),
.B1(n_1540),
.B2(n_1482),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1508),
.B(n_1507),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1479),
.B(n_1498),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1479),
.B(n_1505),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1525),
.A2(n_1502),
.B(n_1501),
.C(n_1530),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1493),
.B(n_1479),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1486),
.A2(n_1474),
.B(n_1485),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1523),
.A2(n_1518),
.B(n_1519),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1482),
.B(n_1542),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1482),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1559),
.B(n_1576),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1572),
.B(n_1489),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1566),
.B(n_1505),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1572),
.B(n_1489),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1577),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1585),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1572),
.B(n_1489),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1547),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1548),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1578),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1595),
.B(n_1568),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1566),
.B(n_1516),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1595),
.B(n_1489),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1555),
.B(n_1475),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1555),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1595),
.B(n_1467),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1592),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1516),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1568),
.B(n_1596),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1545),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1557),
.A2(n_1519),
.B1(n_1493),
.B2(n_1499),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1570),
.B(n_1516),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1565),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1559),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1597),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1578),
.B(n_1471),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1552),
.A2(n_1519),
.B1(n_1499),
.B2(n_1539),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1576),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_SL g1628 ( 
.A(n_1587),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1578),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1578),
.B(n_1471),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1615),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1616),
.B(n_1579),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1615),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1619),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1615),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1626),
.B(n_1562),
.C(n_1573),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1599),
.B(n_1551),
.Y(n_1637)
);

AOI33xp33_ASAP7_75t_L g1638 ( 
.A1(n_1618),
.A2(n_1582),
.A3(n_1575),
.B1(n_1571),
.B2(n_1593),
.B3(n_1586),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1588),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1624),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1624),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1551),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1625),
.B(n_1588),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1625),
.B(n_1630),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1616),
.B(n_1622),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1606),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1622),
.B(n_1579),
.Y(n_1648)
);

OAI221xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1626),
.A2(n_1562),
.B1(n_1573),
.B2(n_1584),
.C(n_1580),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1614),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1603),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1624),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1630),
.B(n_1594),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1620),
.A2(n_1519),
.B1(n_1589),
.B2(n_1582),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1630),
.B(n_1594),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1606),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1620),
.A2(n_1549),
.B1(n_1560),
.B2(n_1558),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1606),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1598),
.Y(n_1659)
);

INVx5_ASAP7_75t_SL g1660 ( 
.A(n_1612),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1618),
.A2(n_1580),
.B1(n_1584),
.B2(n_1561),
.C(n_1571),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_SL g1662 ( 
.A(n_1610),
.B(n_1553),
.C(n_1554),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1604),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1599),
.B(n_1591),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1608),
.B(n_1586),
.Y(n_1665)
);

AOI21xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1618),
.A2(n_1556),
.B(n_1583),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1600),
.A2(n_1495),
.B(n_1478),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1608),
.B(n_1567),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1613),
.B(n_1575),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1606),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1607),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1644),
.B(n_1629),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1634),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1631),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1647),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1631),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1637),
.B(n_1642),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1644),
.B(n_1629),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1656),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1644),
.B(n_1629),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1671),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1648),
.B(n_1613),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1665),
.B(n_1629),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1663),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1663),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1656),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1665),
.B(n_1600),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1665),
.B(n_1600),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1640),
.B(n_1602),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1640),
.B(n_1602),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1636),
.A2(n_1617),
.B1(n_1621),
.B2(n_1627),
.C(n_1602),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1651),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1671),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1648),
.B(n_1613),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1651),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1637),
.B(n_1642),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1642),
.B(n_1617),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1645),
.B(n_1627),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1581),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1631),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1670),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1633),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1645),
.B(n_1604),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1633),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1701),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1691),
.B(n_1653),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1697),
.B(n_1666),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1701),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1687),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1687),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1689),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1697),
.B(n_1638),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1705),
.A2(n_1636),
.B1(n_1661),
.B2(n_1657),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1689),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1698),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1675),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1676),
.B(n_1679),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1685),
.B(n_1638),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1680),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1673),
.A2(n_1661),
.B1(n_1654),
.B2(n_1662),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_L g1727 ( 
.A(n_1676),
.B(n_1649),
.C(n_1662),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1674),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1674),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1677),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1677),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1679),
.B(n_1685),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1675),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1682),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.B(n_1664),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1700),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1709),
.B(n_1619),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1688),
.B(n_1664),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1688),
.B(n_1664),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1691),
.B(n_1653),
.Y(n_1740)
);

OAI33xp33_ASAP7_75t_L g1741 ( 
.A1(n_1704),
.A2(n_1646),
.A3(n_1669),
.B1(n_1544),
.B2(n_1670),
.B3(n_1601),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1675),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1691),
.B(n_1653),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1692),
.B(n_1686),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1682),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1680),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1703),
.B(n_1669),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1601),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1692),
.B(n_1655),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1703),
.B(n_1633),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1684),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1673),
.A2(n_1649),
.B(n_1654),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1704),
.B(n_1635),
.Y(n_1753)
);

NOR3xp33_ASAP7_75t_L g1754 ( 
.A(n_1713),
.B(n_1718),
.C(n_1752),
.Y(n_1754)
);

NAND4xp25_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1657),
.C(n_1564),
.D(n_1550),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1727),
.B(n_1639),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1726),
.B(n_1581),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1639),
.Y(n_1758)
);

NAND2x1_ASAP7_75t_L g1759 ( 
.A(n_1725),
.B(n_1659),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1741),
.A2(n_1597),
.B1(n_1611),
.B2(n_1605),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1744),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1716),
.B(n_1639),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1712),
.B(n_1692),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1717),
.B(n_1643),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_1715),
.B(n_1550),
.C(n_1564),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1720),
.B(n_1643),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1744),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1711),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1728),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1711),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1712),
.B(n_1686),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1728),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1574),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1729),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1729),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1721),
.B(n_1643),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1730),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1723),
.B(n_1655),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1723),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1746),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1730),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1655),
.Y(n_1783)
);

NAND4xp25_ASAP7_75t_SL g1784 ( 
.A(n_1732),
.B(n_1702),
.C(n_1686),
.D(n_1598),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1714),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1746),
.B(n_1678),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1732),
.B(n_1668),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1735),
.B(n_1678),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1740),
.B(n_1672),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1748),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1771),
.Y(n_1791)
);

OA22x2_ASAP7_75t_L g1792 ( 
.A1(n_1757),
.A2(n_1659),
.B1(n_1751),
.B2(n_1745),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1781),
.Y(n_1793)
);

OAI32xp33_ASAP7_75t_L g1794 ( 
.A1(n_1756),
.A2(n_1735),
.A3(n_1739),
.B1(n_1738),
.B2(n_1747),
.Y(n_1794)
);

NAND4xp25_ASAP7_75t_L g1795 ( 
.A(n_1780),
.B(n_1739),
.C(n_1738),
.D(n_1734),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1740),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1781),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1758),
.B(n_1747),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1771),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1774),
.B(n_1753),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1761),
.B(n_1743),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1765),
.B(n_1743),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1760),
.A2(n_1628),
.B1(n_1749),
.B2(n_1660),
.Y(n_1803)
);

INVx1_ASAP7_75t_SL g1804 ( 
.A(n_1768),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1755),
.B(n_1769),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1759),
.B(n_1734),
.C(n_1731),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1770),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1759),
.A2(n_1784),
.B(n_1768),
.Y(n_1808)
);

AOI21xp33_ASAP7_75t_L g1809 ( 
.A1(n_1786),
.A2(n_1753),
.B(n_1733),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1770),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1773),
.A2(n_1611),
.B(n_1605),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1773),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1776),
.B(n_1733),
.C(n_1722),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1766),
.A2(n_1611),
.B(n_1605),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1761),
.A2(n_1767),
.B1(n_1762),
.B2(n_1764),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1792),
.A2(n_1778),
.B(n_1777),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1793),
.B(n_1767),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1797),
.B(n_1763),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1804),
.B(n_1801),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1791),
.B(n_1763),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1799),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1806),
.Y(n_1822)
);

AOI32xp33_ASAP7_75t_L g1823 ( 
.A1(n_1805),
.A2(n_1772),
.A3(n_1789),
.B1(n_1787),
.B2(n_1783),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1790),
.A2(n_1779),
.B1(n_1775),
.B2(n_1782),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1805),
.B(n_1772),
.Y(n_1825)
);

AOI21xp33_ASAP7_75t_L g1826 ( 
.A1(n_1792),
.A2(n_1786),
.B(n_1782),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1800),
.B(n_1789),
.Y(n_1827)
);

AOI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1795),
.A2(n_1775),
.B(n_1788),
.C(n_1722),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1807),
.Y(n_1829)
);

OAI211xp5_ASAP7_75t_L g1830 ( 
.A1(n_1808),
.A2(n_1788),
.B(n_1742),
.C(n_1587),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1802),
.A2(n_1742),
.B(n_1646),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1800),
.B(n_1750),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1796),
.B(n_1749),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1810),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1812),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1819),
.B(n_1820),
.Y(n_1836)
);

O2A1O1Ixp33_ASAP7_75t_SL g1837 ( 
.A1(n_1822),
.A2(n_1794),
.B(n_1809),
.C(n_1803),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1820),
.B(n_1815),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1829),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1829),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1822),
.A2(n_1798),
.B1(n_1813),
.B2(n_1811),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1817),
.Y(n_1842)
);

INVxp33_ASAP7_75t_L g1843 ( 
.A(n_1832),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1830),
.A2(n_1811),
.B(n_1814),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1832),
.A2(n_1628),
.B1(n_1567),
.B2(n_1546),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1818),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1821),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1843),
.B(n_1825),
.Y(n_1848)
);

NAND4xp25_ASAP7_75t_L g1849 ( 
.A(n_1836),
.B(n_1838),
.C(n_1837),
.D(n_1842),
.Y(n_1849)
);

NOR3xp33_ASAP7_75t_L g1850 ( 
.A(n_1846),
.B(n_1827),
.C(n_1824),
.Y(n_1850)
);

NOR4xp25_ASAP7_75t_L g1851 ( 
.A(n_1840),
.B(n_1835),
.C(n_1826),
.D(n_1834),
.Y(n_1851)
);

NAND3xp33_ASAP7_75t_L g1852 ( 
.A(n_1841),
.B(n_1824),
.C(n_1816),
.Y(n_1852)
);

AOI32xp33_ASAP7_75t_L g1853 ( 
.A1(n_1841),
.A2(n_1828),
.A3(n_1833),
.B1(n_1823),
.B2(n_1696),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1844),
.A2(n_1831),
.B1(n_1750),
.B2(n_1696),
.C(n_1695),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1839),
.B(n_1672),
.Y(n_1855)
);

NAND4xp75_ASAP7_75t_L g1856 ( 
.A(n_1847),
.B(n_1696),
.C(n_1695),
.D(n_1672),
.Y(n_1856)
);

NOR3xp33_ASAP7_75t_L g1857 ( 
.A(n_1837),
.B(n_1509),
.C(n_1466),
.Y(n_1857)
);

NAND3xp33_ASAP7_75t_L g1858 ( 
.A(n_1845),
.B(n_1543),
.C(n_1537),
.Y(n_1858)
);

OAI211xp5_ASAP7_75t_L g1859 ( 
.A1(n_1852),
.A2(n_1695),
.B(n_1522),
.C(n_1466),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1857),
.B(n_1678),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1851),
.A2(n_1652),
.B(n_1708),
.C(n_1706),
.Y(n_1861)
);

NOR4xp25_ASAP7_75t_L g1862 ( 
.A(n_1849),
.B(n_1710),
.C(n_1708),
.D(n_1706),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1850),
.A2(n_1609),
.B1(n_1681),
.B2(n_1683),
.C(n_1707),
.Y(n_1863)
);

OAI211xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1853),
.A2(n_1621),
.B(n_1563),
.C(n_1707),
.Y(n_1864)
);

O2A1O1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1848),
.A2(n_1652),
.B(n_1710),
.C(n_1706),
.Y(n_1865)
);

OAI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1862),
.A2(n_1854),
.B1(n_1855),
.B2(n_1858),
.C(n_1856),
.Y(n_1866)
);

NOR2x1p5_ASAP7_75t_L g1867 ( 
.A(n_1859),
.B(n_1522),
.Y(n_1867)
);

OAI322xp33_ASAP7_75t_L g1868 ( 
.A1(n_1861),
.A2(n_1710),
.A3(n_1708),
.B1(n_1652),
.B2(n_1694),
.C1(n_1699),
.C2(n_1690),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1863),
.A2(n_1640),
.B1(n_1683),
.B2(n_1681),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1865),
.B(n_1860),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1864),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1859),
.B(n_1684),
.Y(n_1872)
);

XNOR2xp5_ASAP7_75t_L g1873 ( 
.A(n_1867),
.B(n_1546),
.Y(n_1873)
);

XNOR2xp5_ASAP7_75t_L g1874 ( 
.A(n_1866),
.B(n_1522),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1870),
.B(n_1690),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1871),
.Y(n_1876)
);

XNOR2xp5_ASAP7_75t_L g1877 ( 
.A(n_1872),
.B(n_1541),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1874),
.A2(n_1868),
.B(n_1869),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1876),
.B(n_1693),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1875),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1880),
.B(n_1873),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1881),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1882),
.A2(n_1878),
.B(n_1879),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1882),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1884),
.A2(n_1877),
.B1(n_1681),
.B2(n_1683),
.Y(n_1885)
);

OAI22x1_ASAP7_75t_L g1886 ( 
.A1(n_1883),
.A2(n_1509),
.B1(n_1466),
.B2(n_1520),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1886),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1885),
.A2(n_1699),
.B(n_1694),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1887),
.B(n_1693),
.Y(n_1889)
);

OAI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1889),
.A2(n_1888),
.B1(n_1641),
.B2(n_1536),
.Y(n_1890)
);

XNOR2xp5_ASAP7_75t_L g1891 ( 
.A(n_1890),
.B(n_1487),
.Y(n_1891)
);

OAI221xp5_ASAP7_75t_R g1892 ( 
.A1(n_1891),
.A2(n_1641),
.B1(n_1660),
.B2(n_1650),
.C(n_1667),
.Y(n_1892)
);

AOI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1536),
.B(n_1500),
.C(n_1510),
.Y(n_1893)
);


endmodule