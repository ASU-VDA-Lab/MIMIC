module fake_ariane_2374_n_1651 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1651);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1651;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_SL g159 ( 
.A(n_106),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_82),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_25),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_51),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_54),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_100),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_58),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_80),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_56),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_81),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_27),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_99),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_50),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_89),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_49),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_116),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_9),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_15),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_0),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_41),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_11),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_121),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_25),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_38),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_91),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_33),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_3),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_84),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_131),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_15),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_3),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_51),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_28),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_145),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_13),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_74),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_75),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_62),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_1),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_138),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_55),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_23),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_137),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_76),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_63),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_86),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_107),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_152),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_127),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_156),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_21),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_37),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_85),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_115),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_19),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_151),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_27),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_139),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_130),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_154),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_17),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_117),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_105),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_37),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_102),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_149),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_73),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_119),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_110),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_71),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_18),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_109),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_45),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_45),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_118),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_111),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_46),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_46),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_67),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_2),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_147),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_77),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_90),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_30),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_6),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_14),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_132),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_83),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_79),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_26),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_61),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_64),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_69),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_0),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_135),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_142),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_146),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_103),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_24),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_41),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_32),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_141),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_60),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_16),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_87),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_113),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_88),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_43),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_16),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_223),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_186),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_181),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_265),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_309),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_161),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_161),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_169),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_169),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_246),
.B(n_2),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_183),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_257),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_188),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_201),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_222),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_183),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_205),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_210),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_205),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_166),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_186),
.B(n_5),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_224),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_5),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_243),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_248),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_163),
.B(n_6),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_164),
.B(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_249),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_167),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_243),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_261),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_167),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_262),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_291),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_291),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_317),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_165),
.B(n_9),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_172),
.B(n_10),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_317),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_206),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_174),
.B(n_12),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_223),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_206),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_223),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_209),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_236),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_177),
.B(n_12),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_236),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_209),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_167),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_278),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_278),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_263),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_234),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_236),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_283),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_271),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_234),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_283),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_160),
.B(n_150),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_263),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_271),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_263),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_271),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_168),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_305),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_275),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_168),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_171),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_312),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_171),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_305),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_331),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

BUFx10_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_379),
.B(n_175),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_330),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_320),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_330),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_371),
.A2(n_192),
.B(n_190),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_333),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_380),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_159),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_397),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_159),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_333),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_393),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_347),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_334),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_198),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_348),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_342),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_346),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_366),
.B(n_180),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_350),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_351),
.B(n_178),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_356),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_362),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_334),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_367),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_369),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_398),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_357),
.A2(n_189),
.B(n_184),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_338),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_374),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_358),
.B(n_208),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_325),
.B(n_320),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_406),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_378),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_349),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_379),
.B(n_175),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_338),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_344),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_352),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_335),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_344),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_370),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_419),
.B(n_324),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_426),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_426),
.B(n_400),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_447),
.B(n_322),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_R g493 ( 
.A(n_418),
.B(n_345),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_440),
.A2(n_329),
.B1(n_328),
.B2(n_409),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_434),
.B(n_326),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_411),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_434),
.B(n_326),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_466),
.A2(n_328),
.B1(n_329),
.B2(n_401),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_434),
.B(n_190),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_434),
.B(n_381),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_466),
.A2(n_394),
.B1(n_381),
.B2(n_401),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_486),
.A2(n_390),
.B1(n_353),
.B2(n_268),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_432),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_466),
.A2(n_473),
.B1(n_486),
.B2(n_480),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_434),
.B(n_383),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_428),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_383),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_440),
.A2(n_385),
.B1(n_399),
.B2(n_394),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_426),
.B(n_405),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_414),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_439),
.A2(n_385),
.B1(n_399),
.B2(n_392),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_445),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_392),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_427),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_443),
.B(n_173),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_449),
.B(n_345),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_448),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_434),
.B(n_192),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_457),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_457),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_443),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_449),
.B(n_198),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_458),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_466),
.A2(n_275),
.B1(n_167),
.B2(n_293),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_438),
.B(n_355),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_L g543 ( 
.A(n_485),
.B(n_215),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_485),
.B(n_215),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_419),
.B(n_227),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_419),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_466),
.A2(n_275),
.B1(n_293),
.B2(n_239),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_434),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_415),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_478),
.A2(n_480),
.B1(n_481),
.B2(n_477),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_438),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_252),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_421),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_485),
.B(n_217),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_465),
.B(n_355),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_421),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_459),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_453),
.A2(n_410),
.B1(n_404),
.B2(n_395),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_421),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_414),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_413),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_439),
.B(n_176),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_441),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_477),
.B(n_476),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_473),
.A2(n_293),
.B1(n_214),
.B2(n_268),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_464),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_478),
.A2(n_361),
.B1(n_375),
.B2(n_220),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_417),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_465),
.B(n_361),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_424),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_481),
.B(n_375),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_485),
.B(n_226),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_488),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_416),
.B(n_233),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_460),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_460),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_482),
.B(n_235),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_446),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_417),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_454),
.B(n_173),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_472),
.Y(n_590)
);

CKINVDCx6p67_ASAP7_75t_R g591 ( 
.A(n_472),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_453),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_471),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_485),
.B(n_237),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_485),
.A2(n_214),
.B1(n_196),
.B2(n_296),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_422),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_422),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_448),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_423),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_448),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_460),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_460),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_454),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_460),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_476),
.B(n_185),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_469),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_448),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_469),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_424),
.B(n_456),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_430),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_430),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_430),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_461),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_469),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_456),
.B(n_196),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_469),
.B(n_456),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_467),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_437),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_454),
.B(n_185),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_469),
.B(n_241),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_469),
.B(n_245),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_437),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_437),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_483),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_541),
.A2(n_469),
.B1(n_450),
.B2(n_462),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_552),
.A2(n_456),
.B(n_462),
.C(n_463),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_569),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_525),
.B(n_475),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_568),
.B(n_479),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_583),
.A2(n_429),
.B(n_470),
.C(n_463),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_512),
.B(n_554),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_497),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_492),
.B(n_462),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_490),
.B(n_462),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_499),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_530),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_SL g640 ( 
.A(n_494),
.B(n_517),
.C(n_526),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_490),
.B(n_463),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_575),
.B(n_484),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_586),
.A2(n_479),
.B1(n_463),
.B2(n_470),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_536),
.B(n_470),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_470),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_537),
.A2(n_455),
.B1(n_450),
.B2(n_487),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_525),
.B(n_455),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_582),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_568),
.B(n_429),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_497),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_606),
.B(n_450),
.Y(n_651)
);

O2A1O1Ixp5_ASAP7_75t_L g652 ( 
.A1(n_568),
.A2(n_450),
.B(n_276),
.C(n_433),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_569),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_498),
.B(n_433),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_606),
.B(n_474),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_515),
.B(n_474),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_491),
.B(n_474),
.Y(n_657)
);

INVx8_ASAP7_75t_L g658 ( 
.A(n_608),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_545),
.B(n_444),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_520),
.B(n_391),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_548),
.A2(n_444),
.B1(n_442),
.B2(n_436),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_496),
.B(n_444),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_616),
.B(n_620),
.C(n_576),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_503),
.A2(n_442),
.B1(n_436),
.B2(n_435),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_590),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_522),
.B(n_242),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_506),
.B(n_511),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_567),
.B(n_242),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_523),
.B(n_318),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_570),
.B(n_429),
.Y(n_670)
);

NOR2x1_ASAP7_75t_L g671 ( 
.A(n_489),
.B(n_250),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_505),
.A2(n_319),
.B1(n_318),
.B2(n_315),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_519),
.B(n_319),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_524),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_498),
.B(n_195),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_618),
.A2(n_296),
.B1(n_314),
.B2(n_264),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_582),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_580),
.B(n_197),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_529),
.B(n_199),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_537),
.A2(n_316),
.B1(n_253),
.B2(n_313),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_612),
.A2(n_281),
.B(n_306),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_500),
.B(n_200),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_528),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_553),
.B(n_202),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_618),
.A2(n_314),
.B1(n_258),
.B2(n_274),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_564),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_507),
.B(n_207),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_505),
.A2(n_304),
.B(n_300),
.C(n_279),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_553),
.B(n_216),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_SL g690 ( 
.A(n_547),
.B(n_218),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_533),
.B(n_219),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_577),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_535),
.B(n_225),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_572),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_542),
.B(n_238),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g696 ( 
.A(n_524),
.B(n_254),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_539),
.B(n_256),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_627),
.B(n_266),
.C(n_267),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_588),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_538),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_537),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_540),
.B(n_560),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_526),
.Y(n_703)
);

BUFx8_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_513),
.B(n_273),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_561),
.B(n_277),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_566),
.B(n_280),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_537),
.A2(n_282),
.B1(n_284),
.B2(n_307),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_587),
.B(n_288),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_618),
.A2(n_294),
.B1(n_303),
.B2(n_299),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_527),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_618),
.A2(n_182),
.B1(n_286),
.B2(n_211),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_579),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_513),
.B(n_17),
.Y(n_714)
);

BUFx6f_ASAP7_75t_SL g715 ( 
.A(n_573),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_547),
.B(n_170),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_549),
.B(n_18),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_527),
.B(n_179),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_595),
.B(n_187),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_R g720 ( 
.A(n_493),
.B(n_191),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_591),
.B(n_20),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_538),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_578),
.B(n_182),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_573),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_588),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_549),
.B(n_20),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_527),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_549),
.B(n_21),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_573),
.B(n_589),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_618),
.B(n_215),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_579),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_601),
.B(n_193),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_589),
.B(n_194),
.Y(n_733)
);

INVx8_ASAP7_75t_L g734 ( 
.A(n_608),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_495),
.B(n_215),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_592),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_556),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_573),
.A2(n_608),
.B1(n_556),
.B2(n_596),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_618),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_589),
.B(n_203),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_622),
.B(n_204),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_622),
.B(n_212),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_622),
.B(n_308),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_543),
.A2(n_302),
.B(n_298),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_562),
.B(n_182),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_574),
.B(n_247),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_251),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_593),
.B(n_244),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_608),
.A2(n_255),
.B1(n_297),
.B2(n_292),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_598),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_495),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_495),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_591),
.B(n_240),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_531),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_599),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_581),
.A2(n_232),
.B(n_289),
.C(n_213),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_510),
.B(n_259),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_613),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_594),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_510),
.B(n_231),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_619),
.B(n_29),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_510),
.B(n_260),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_594),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_613),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_614),
.B(n_228),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_501),
.B(n_502),
.Y(n_766)
);

BUFx12f_ASAP7_75t_L g767 ( 
.A(n_504),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_614),
.B(n_221),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_597),
.A2(n_310),
.B1(n_286),
.B2(n_211),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_615),
.A2(n_215),
.B1(n_270),
.B2(n_269),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_615),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_714),
.A2(n_596),
.B(n_543),
.C(n_544),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_649),
.A2(n_544),
.B(n_501),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_633),
.A2(n_619),
.B(n_558),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_656),
.B(n_621),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_714),
.A2(n_565),
.B1(n_603),
.B2(n_607),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_638),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_705),
.A2(n_603),
.B(n_565),
.C(n_607),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_667),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_670),
.A2(n_559),
.B(n_555),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_686),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_766),
.A2(n_502),
.B(n_508),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_644),
.A2(n_508),
.B(n_514),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_705),
.A2(n_603),
.B(n_565),
.C(n_607),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_636),
.A2(n_521),
.B1(n_514),
.B2(n_534),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_674),
.B(n_621),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_735),
.A2(n_605),
.B(n_609),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_655),
.B(n_625),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_662),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_703),
.B(n_516),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_645),
.A2(n_514),
.B(n_521),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_713),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_629),
.A2(n_559),
.B(n_555),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_647),
.B(n_625),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_651),
.A2(n_521),
.B(n_534),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_764),
.B(n_626),
.Y(n_796)
);

AOI21x1_ASAP7_75t_L g797 ( 
.A1(n_735),
.A2(n_611),
.B(n_617),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_771),
.Y(n_798)
);

OAI21xp33_ASAP7_75t_L g799 ( 
.A1(n_709),
.A2(n_518),
.B(n_563),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_637),
.A2(n_518),
.B(n_516),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_713),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_729),
.B(n_626),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_646),
.B(n_546),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_646),
.B(n_546),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_641),
.A2(n_516),
.B(n_563),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_702),
.A2(n_563),
.B1(n_571),
.B2(n_584),
.Y(n_806)
);

AO21x1_ASAP7_75t_L g807 ( 
.A1(n_634),
.A2(n_571),
.B(n_584),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_657),
.B(n_550),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_643),
.B(n_551),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_694),
.B(n_624),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_729),
.B(n_531),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_686),
.B(n_584),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_630),
.Y(n_813)
);

OAI21xp33_ASAP7_75t_L g814 ( 
.A1(n_675),
.A2(n_624),
.B(n_623),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_632),
.A2(n_604),
.B(n_602),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_652),
.A2(n_610),
.B(n_604),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_639),
.B(n_610),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_660),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_659),
.A2(n_509),
.B(n_585),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_675),
.B(n_504),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_695),
.B(n_532),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_680),
.B(n_600),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_680),
.B(n_600),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_745),
.A2(n_532),
.B1(n_504),
.B2(n_546),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_653),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_682),
.B(n_711),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_682),
.B(n_504),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_752),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_684),
.B(n_532),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_708),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_640),
.B(n_600),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_761),
.A2(n_504),
.B(n_532),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_708),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_761),
.A2(n_585),
.B1(n_509),
.B2(n_546),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_654),
.A2(n_600),
.B(n_531),
.C(n_272),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_631),
.A2(n_678),
.B(n_669),
.C(n_691),
.Y(n_836)
);

BUFx12f_ASAP7_75t_L g837 ( 
.A(n_763),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_739),
.B(n_532),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_720),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_642),
.B(n_532),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_724),
.B(n_35),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_719),
.A2(n_270),
.B(n_215),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_715),
.A2(n_270),
.B1(n_36),
.B2(n_38),
.Y(n_843)
);

AOI33xp33_ASAP7_75t_L g844 ( 
.A1(n_737),
.A2(n_35),
.A3(n_39),
.B1(n_42),
.B2(n_43),
.B3(n_44),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_724),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_732),
.A2(n_747),
.B(n_748),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_679),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_727),
.B(n_52),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_654),
.B(n_52),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_704),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_731),
.B(n_53),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_SL g852 ( 
.A(n_663),
.B(n_270),
.C(n_57),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_739),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_753),
.B(n_59),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_751),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_701),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_759),
.B(n_114),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_664),
.B(n_136),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_693),
.A2(n_697),
.B(n_706),
.C(n_707),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_692),
.A2(n_725),
.B(n_699),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_721),
.B(n_712),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_736),
.A2(n_750),
.B(n_755),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_673),
.A2(n_768),
.B(n_765),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_717),
.A2(n_726),
.B1(n_728),
.B2(n_710),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_665),
.B(n_648),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_715),
.A2(n_738),
.B1(n_701),
.B2(n_672),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_758),
.Y(n_867)
);

INVx5_ASAP7_75t_L g868 ( 
.A(n_767),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_687),
.A2(n_689),
.B(n_726),
.C(n_728),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_681),
.A2(n_688),
.B(n_756),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_671),
.A2(n_668),
.B(n_666),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_704),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_723),
.B(n_718),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_664),
.B(n_661),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_658),
.B(n_734),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_749),
.B(n_710),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_658),
.B(n_734),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_635),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_685),
.A2(n_676),
.B1(n_712),
.B2(n_628),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_650),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_730),
.A2(n_742),
.B(n_740),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_658),
.B(n_743),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_733),
.A2(n_741),
.B(n_752),
.Y(n_883)
);

OAI321xp33_ASAP7_75t_L g884 ( 
.A1(n_685),
.A2(n_676),
.A3(n_745),
.B1(n_762),
.B2(n_760),
.C(n_757),
.Y(n_884)
);

INVx3_ASAP7_75t_SL g885 ( 
.A(n_723),
.Y(n_885)
);

OA21x2_ASAP7_75t_L g886 ( 
.A1(n_683),
.A2(n_722),
.B(n_700),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_720),
.B(n_698),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_628),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_746),
.B(n_690),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_754),
.B(n_744),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_770),
.B(n_769),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_770),
.B(n_769),
.Y(n_892)
);

CKINVDCx10_ASAP7_75t_R g893 ( 
.A(n_677),
.Y(n_893)
);

AOI22x1_ASAP7_75t_L g894 ( 
.A1(n_696),
.A2(n_485),
.B1(n_549),
.B2(n_547),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_667),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_656),
.B(n_490),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_694),
.B(n_330),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_640),
.B(n_620),
.C(n_616),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_646),
.B(n_729),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_L g902 ( 
.A1(n_709),
.A2(n_580),
.B(n_492),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_640),
.A2(n_646),
.B1(n_729),
.B2(n_705),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_714),
.A2(n_705),
.B(n_654),
.C(n_682),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_656),
.B(n_490),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_638),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_667),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_714),
.A2(n_512),
.B1(n_552),
.B2(n_480),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_752),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_656),
.B(n_490),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_640),
.A2(n_646),
.B1(n_729),
.B2(n_705),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_656),
.B(n_490),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_680),
.A2(n_552),
.B(n_580),
.C(n_708),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_767),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_714),
.A2(n_512),
.B1(n_552),
.B2(n_480),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_694),
.B(n_330),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_657),
.B(n_491),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_922)
);

O2A1O1Ixp5_ASAP7_75t_L g923 ( 
.A1(n_649),
.A2(n_568),
.B(n_513),
.C(n_505),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_656),
.B(n_490),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_771),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_656),
.B(n_490),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_SL g928 ( 
.A1(n_716),
.A2(n_649),
.B(n_636),
.C(n_633),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_656),
.B(n_490),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_752),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_649),
.A2(n_568),
.B(n_670),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_895),
.A2(n_905),
.B(n_900),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_906),
.A2(n_921),
.B(n_916),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_861),
.A2(n_818),
.B1(n_876),
.B2(n_874),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_L g936 ( 
.A(n_864),
.B(n_904),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_878),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_915),
.A2(n_902),
.B(n_864),
.C(n_869),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_779),
.B(n_896),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_922),
.A2(n_931),
.B(n_925),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_880),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_828),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_910),
.A2(n_918),
.B1(n_849),
.B2(n_909),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_813),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_828),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_920),
.B(n_898),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_786),
.B(n_919),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_897),
.B(n_907),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_774),
.A2(n_918),
.B(n_910),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_844),
.A2(n_914),
.B(n_912),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_780),
.A2(n_773),
.B(n_774),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_780),
.A2(n_793),
.B(n_787),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_789),
.B(n_924),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_927),
.B(n_929),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_825),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_793),
.A2(n_797),
.B(n_816),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_903),
.A2(n_913),
.B(n_859),
.C(n_836),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_839),
.B(n_826),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_846),
.A2(n_928),
.B(n_863),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_781),
.B(n_899),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_923),
.A2(n_772),
.B(n_778),
.Y(n_961)
);

INVx5_ASAP7_75t_L g962 ( 
.A(n_850),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_SL g963 ( 
.A1(n_879),
.A2(n_853),
.B(n_834),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_890),
.A2(n_791),
.B(n_795),
.Y(n_964)
);

OA21x2_ASAP7_75t_L g965 ( 
.A1(n_784),
.A2(n_842),
.B(n_816),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_783),
.A2(n_834),
.B(n_785),
.Y(n_966)
);

AO31x2_ASAP7_75t_L g967 ( 
.A1(n_835),
.A2(n_883),
.A3(n_776),
.B(n_820),
.Y(n_967)
);

AO31x2_ASAP7_75t_L g968 ( 
.A1(n_776),
.A2(n_827),
.A3(n_862),
.B(n_860),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_841),
.B(n_856),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_802),
.B(n_796),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_800),
.A2(n_805),
.B(n_815),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_777),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_881),
.A2(n_775),
.B(n_804),
.Y(n_973)
);

NOR2x1_ASAP7_75t_L g974 ( 
.A(n_792),
.B(n_801),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_889),
.A2(n_782),
.B(n_819),
.Y(n_975)
);

AO21x1_ASAP7_75t_L g976 ( 
.A1(n_858),
.A2(n_803),
.B(n_831),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_SL g977 ( 
.A1(n_830),
.A2(n_833),
.B(n_845),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_841),
.B(n_885),
.Y(n_978)
);

AND3x4_ASAP7_75t_L g979 ( 
.A(n_865),
.B(n_810),
.C(n_893),
.Y(n_979)
);

NAND2x1_ASAP7_75t_L g980 ( 
.A(n_828),
.B(n_911),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_872),
.B(n_875),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_870),
.A2(n_809),
.B(n_832),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_806),
.A2(n_788),
.B(n_799),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_867),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_814),
.A2(n_840),
.B(n_817),
.C(n_852),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_808),
.Y(n_986)
);

AOI21x1_ASAP7_75t_SL g987 ( 
.A1(n_851),
.A2(n_848),
.B(n_821),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_837),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_887),
.B(n_866),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_871),
.A2(n_894),
.B(n_901),
.Y(n_990)
);

OAI21x1_ASAP7_75t_SL g991 ( 
.A1(n_798),
.A2(n_926),
.B(n_882),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_847),
.A2(n_873),
.B(n_884),
.C(n_823),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_794),
.B(n_792),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_908),
.B(n_801),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_812),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_888),
.A2(n_829),
.B1(n_891),
.B2(n_892),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_911),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_855),
.B(n_930),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_911),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_877),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_838),
.A2(n_886),
.B(n_822),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_811),
.B(n_855),
.Y(n_1002)
);

AOI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_843),
.A2(n_824),
.B(n_854),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_930),
.A2(n_838),
.B(n_857),
.Y(n_1004)
);

AND2x6_ASAP7_75t_SL g1005 ( 
.A(n_790),
.B(n_868),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_868),
.A2(n_932),
.B(n_931),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_868),
.A2(n_568),
.B(n_864),
.Y(n_1007)
);

NAND2x1_ASAP7_75t_L g1008 ( 
.A(n_868),
.B(n_917),
.Y(n_1008)
);

OA21x2_ASAP7_75t_L g1009 ( 
.A1(n_917),
.A2(n_900),
.B(n_895),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_917),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_917),
.A2(n_932),
.B(n_931),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_904),
.A2(n_915),
.B(n_902),
.C(n_864),
.Y(n_1012)
);

INVx8_ASAP7_75t_L g1013 ( 
.A(n_850),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_895),
.A2(n_649),
.B(n_931),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_779),
.B(n_896),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_895),
.A2(n_932),
.B(n_931),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_904),
.A2(n_915),
.B(n_902),
.C(n_864),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_910),
.A2(n_918),
.B1(n_904),
.B2(n_864),
.Y(n_1020)
);

OR2x6_ASAP7_75t_L g1021 ( 
.A(n_850),
.B(n_658),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_864),
.A2(n_918),
.B(n_910),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_864),
.A2(n_918),
.B(n_910),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_SL g1025 ( 
.A1(n_904),
.A2(n_864),
.B(n_879),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_841),
.B(n_739),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_779),
.B(n_896),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_920),
.B(n_491),
.Y(n_1029)
);

BUFx8_ASAP7_75t_SL g1030 ( 
.A(n_837),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_779),
.B(n_896),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_779),
.B(n_896),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_850),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_895),
.A2(n_932),
.B(n_931),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_920),
.B(n_491),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_902),
.B(n_709),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_920),
.B(n_491),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_807),
.A2(n_864),
.A3(n_900),
.B(n_895),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_828),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_895),
.A2(n_932),
.B(n_931),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_868),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_875),
.B(n_877),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_828),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_875),
.B(n_877),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_813),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_813),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_904),
.A2(n_864),
.B(n_633),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_779),
.B(n_896),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_828),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_868),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_813),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_895),
.A2(n_649),
.B(n_931),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_850),
.Y(n_1055)
);

AO31x2_ASAP7_75t_L g1056 ( 
.A1(n_807),
.A2(n_864),
.A3(n_900),
.B(n_895),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_828),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_828),
.Y(n_1058)
);

AO21x1_ASAP7_75t_L g1059 ( 
.A1(n_864),
.A2(n_918),
.B(n_910),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_818),
.B(n_499),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_902),
.A2(n_526),
.B1(n_703),
.B2(n_898),
.Y(n_1061)
);

INVx6_ASAP7_75t_L g1062 ( 
.A(n_850),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_SL g1063 ( 
.A1(n_904),
.A2(n_864),
.B(n_879),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_813),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_864),
.A2(n_568),
.B(n_904),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_828),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_861),
.A2(n_745),
.B1(n_333),
.B2(n_334),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_868),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_989),
.B(n_947),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_1023),
.A2(n_949),
.B(n_957),
.C(n_1020),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_946),
.B(n_1029),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_939),
.B(n_1015),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_1013),
.Y(n_1073)
);

INVx3_ASAP7_75t_SL g1074 ( 
.A(n_1013),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1020),
.A2(n_1023),
.B1(n_949),
.B2(n_1063),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1012),
.A2(n_1017),
.B1(n_1061),
.B2(n_938),
.Y(n_1076)
);

AO21x2_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_1019),
.B(n_1018),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1036),
.B(n_1039),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_R g1079 ( 
.A(n_962),
.B(n_1062),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_962),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_969),
.B(n_978),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_L g1082 ( 
.A(n_979),
.B(n_1043),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_972),
.B(n_1060),
.Y(n_1083)
);

OAI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_936),
.A2(n_1025),
.B(n_1019),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_943),
.A2(n_1026),
.B1(n_1067),
.B2(n_1015),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1022),
.A2(n_1059),
.B1(n_943),
.B2(n_977),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_944),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_1013),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_994),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_937),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_939),
.B(n_1028),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1028),
.B(n_1050),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_958),
.B(n_1050),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1026),
.B(n_1021),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_1010),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_SL g1096 ( 
.A(n_1026),
.B(n_992),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_962),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_984),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_941),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_1021),
.B(n_981),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1065),
.A2(n_1027),
.B(n_1024),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1047),
.B(n_1048),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_970),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_945),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1018),
.A2(n_1037),
.B(n_1035),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_960),
.B(n_953),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1053),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_954),
.B(n_948),
.Y(n_1109)
);

OAI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1024),
.A2(n_1037),
.B1(n_1027),
.B2(n_1035),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_1008),
.B(n_963),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1000),
.B(n_986),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1049),
.A2(n_1064),
.B(n_950),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_L g1114 ( 
.A(n_1062),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_935),
.B(n_1000),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_985),
.B(n_959),
.C(n_961),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1026),
.B(n_1044),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1003),
.A2(n_982),
.B(n_1007),
.C(n_990),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1046),
.B(n_993),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_996),
.B(n_998),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_966),
.A2(n_983),
.B(n_964),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_975),
.A2(n_940),
.B(n_973),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1002),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_998),
.B(n_1045),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_945),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_974),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_942),
.B(n_1045),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_995),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_951),
.A2(n_956),
.B(n_952),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_971),
.A2(n_933),
.B(n_934),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_976),
.A2(n_991),
.B(n_942),
.C(n_1041),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_1030),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1041),
.B(n_1057),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1057),
.B(n_1068),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_1052),
.B(n_1004),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1052),
.A2(n_1066),
.B1(n_1058),
.B2(n_1051),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1016),
.A2(n_1042),
.B(n_1034),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1033),
.A2(n_1055),
.B1(n_988),
.B2(n_1058),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_997),
.B(n_1066),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_999),
.B(n_1051),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1001),
.A2(n_1011),
.B(n_1006),
.C(n_980),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1058),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1005),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_1005),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1009),
.A2(n_965),
.B1(n_1054),
.B2(n_1014),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1009),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_967),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1040),
.B(n_1056),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_987),
.B(n_1040),
.C(n_967),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_968),
.A2(n_1020),
.B1(n_1023),
.B2(n_949),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_968),
.A2(n_936),
.B(n_1020),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1026),
.B(n_875),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1060),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1060),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_SL g1155 ( 
.A1(n_1023),
.A2(n_1020),
.B(n_1038),
.C(n_1018),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1061),
.B(n_989),
.Y(n_1156)
);

INVx3_ASAP7_75t_SL g1157 ( 
.A(n_1013),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1061),
.B(n_989),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1010),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1026),
.B(n_875),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_946),
.B(n_939),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1060),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_1026),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1026),
.B(n_875),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_946),
.B(n_1029),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1023),
.A2(n_949),
.B(n_982),
.Y(n_1166)
);

AOI221x1_ASAP7_75t_L g1167 ( 
.A1(n_1023),
.A2(n_1020),
.B1(n_1063),
.B2(n_1025),
.C(n_1017),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_955),
.Y(n_1168)
);

AND2x4_ASAP7_75t_SL g1169 ( 
.A(n_1021),
.B(n_524),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_940),
.A2(n_1023),
.B(n_1019),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1010),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1013),
.Y(n_1172)
);

OR2x6_ASAP7_75t_L g1173 ( 
.A(n_1021),
.B(n_658),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1026),
.B(n_875),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_936),
.A2(n_1020),
.B(n_1023),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_972),
.Y(n_1176)
);

INVx3_ASAP7_75t_SL g1177 ( 
.A(n_1013),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_946),
.B(n_939),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1023),
.A2(n_1022),
.B(n_1059),
.C(n_1020),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1020),
.A2(n_1023),
.B1(n_949),
.B2(n_1025),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_989),
.B(n_330),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_955),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_946),
.B(n_1029),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1026),
.B(n_875),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_936),
.A2(n_1020),
.B(n_1023),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_947),
.B(n_1060),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1026),
.B(n_875),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1030),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_946),
.B(n_939),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1030),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1023),
.A2(n_904),
.B(n_915),
.C(n_902),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_945),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_946),
.B(n_1029),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_1023),
.A2(n_1022),
.B(n_1059),
.C(n_1020),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1023),
.A2(n_904),
.B(n_915),
.C(n_902),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1069),
.B(n_1093),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1103),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1086),
.A2(n_1167),
.B1(n_1075),
.B2(n_1180),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1108),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1094),
.B(n_1163),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1073),
.Y(n_1201)
);

BUFx4f_ASAP7_75t_L g1202 ( 
.A(n_1074),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1137),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1163),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1087),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1147),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1099),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1071),
.B(n_1165),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1188),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1181),
.A2(n_1156),
.B1(n_1158),
.B2(n_1096),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_1132),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1086),
.A2(n_1180),
.B1(n_1075),
.B2(n_1110),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1168),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1129),
.A2(n_1118),
.B(n_1116),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1183),
.B(n_1193),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1172),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1182),
.Y(n_1217)
);

NOR2x1_ASAP7_75t_R g1218 ( 
.A(n_1190),
.B(n_1114),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1084),
.A2(n_1076),
.B1(n_1085),
.B2(n_1106),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1084),
.A2(n_1106),
.B1(n_1175),
.B2(n_1185),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1145),
.A2(n_1135),
.B(n_1148),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1186),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1123),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1090),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1100),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1080),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1078),
.B(n_1081),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1112),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1083),
.B(n_1161),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1080),
.Y(n_1230)
);

CKINVDCx11_ASAP7_75t_R g1231 ( 
.A(n_1157),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1151),
.A2(n_1102),
.B(n_1147),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1119),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1072),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1102),
.A2(n_1130),
.B(n_1116),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1177),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1178),
.B(n_1189),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1096),
.A2(n_1150),
.B1(n_1115),
.B2(n_1077),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1105),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1150),
.A2(n_1109),
.B1(n_1092),
.B2(n_1091),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1166),
.A2(n_1107),
.B1(n_1146),
.B2(n_1104),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1089),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1153),
.B(n_1154),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1124),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1097),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1162),
.B(n_1169),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1170),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1166),
.A2(n_1144),
.B1(n_1117),
.B2(n_1120),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1070),
.A2(n_1195),
.B1(n_1191),
.B2(n_1176),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1149),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1149),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1098),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1128),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1101),
.A2(n_1174),
.B1(n_1184),
.B2(n_1164),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1139),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1160),
.B2(n_1152),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1105),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1126),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1095),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1179),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1127),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1184),
.A2(n_1187),
.B1(n_1173),
.B2(n_1082),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1133),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1113),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1194),
.A2(n_1155),
.B(n_1131),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1187),
.B(n_1111),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1111),
.Y(n_1267)
);

CKINVDCx8_ASAP7_75t_R g1268 ( 
.A(n_1095),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1140),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1095),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1134),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1192),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1088),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1192),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1159),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1125),
.B(n_1138),
.Y(n_1276)
);

CKINVDCx16_ASAP7_75t_R g1277 ( 
.A(n_1138),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1171),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1125),
.B(n_1142),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1136),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1141),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1171),
.A2(n_1023),
.B1(n_1059),
.B2(n_1022),
.Y(n_1282)
);

AO21x1_ASAP7_75t_L g1283 ( 
.A1(n_1079),
.A2(n_1020),
.B(n_943),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1079),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1156),
.B(n_1158),
.Y(n_1285)
);

BUFx8_ASAP7_75t_L g1286 ( 
.A(n_1114),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1103),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1086),
.A2(n_1020),
.B1(n_1023),
.B2(n_1167),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1103),
.Y(n_1289)
);

AO21x1_ASAP7_75t_L g1290 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_943),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1103),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1103),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1080),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1103),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1147),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1086),
.A2(n_1070),
.B1(n_1020),
.B2(n_1075),
.Y(n_1296)
);

AO21x1_ASAP7_75t_L g1297 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_943),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1163),
.B(n_1094),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1211),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1265),
.A2(n_1198),
.B(n_1212),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1211),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1210),
.A2(n_1296),
.B1(n_1198),
.B2(n_1288),
.Y(n_1302)
);

BUFx2_ASAP7_75t_SL g1303 ( 
.A(n_1283),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1199),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_SL g1305 ( 
.A(n_1209),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1251),
.B(n_1238),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1238),
.B(n_1250),
.Y(n_1307)
);

AO21x1_ASAP7_75t_SL g1308 ( 
.A1(n_1220),
.A2(n_1219),
.B(n_1250),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1212),
.A2(n_1247),
.B(n_1240),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1214),
.B(n_1197),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1288),
.A2(n_1297),
.B1(n_1290),
.B2(n_1219),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1281),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1266),
.B(n_1267),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1232),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1271),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1255),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1281),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1214),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1286),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1214),
.B(n_1287),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1240),
.A2(n_1260),
.B(n_1221),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1289),
.B(n_1291),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1206),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1206),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1242),
.B(n_1196),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1295),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1295),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1235),
.A2(n_1220),
.B(n_1280),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1203),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1258),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1205),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1207),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1229),
.B(n_1237),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1234),
.B(n_1245),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1264),
.A2(n_1203),
.B(n_1249),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1223),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1282),
.A2(n_1254),
.B(n_1262),
.Y(n_1338)
);

AOI221xp5_ASAP7_75t_L g1339 ( 
.A1(n_1285),
.A2(n_1253),
.B1(n_1282),
.B2(n_1263),
.C(n_1261),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1285),
.A2(n_1241),
.B1(n_1269),
.B2(n_1225),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1243),
.B(n_1269),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1222),
.B(n_1244),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1228),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1208),
.B(n_1215),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_SL g1345 ( 
.A(n_1286),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1233),
.B(n_1227),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1213),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1217),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1224),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1272),
.B(n_1274),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1248),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1257),
.B(n_1246),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1279),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1256),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1286),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1262),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1310),
.B(n_1320),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1320),
.B(n_1239),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1332),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1332),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1309),
.B(n_1252),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1323),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1338),
.B(n_1298),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1309),
.B(n_1239),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1323),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1303),
.B(n_1201),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1318),
.B(n_1200),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1327),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1312),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1324),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1309),
.B(n_1226),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1315),
.B(n_1293),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1312),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1317),
.B(n_1230),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1328),
.B(n_1201),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1324),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1317),
.B(n_1216),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1313),
.B(n_1284),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1326),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1302),
.A2(n_1278),
.B1(n_1275),
.B2(n_1204),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1328),
.B(n_1216),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1303),
.B(n_1273),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1307),
.B(n_1306),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1300),
.A2(n_1278),
.B1(n_1275),
.B2(n_1204),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1326),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1300),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1343),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1388),
.B(n_1358),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1388),
.B(n_1304),
.Y(n_1390)
);

OA211x2_ASAP7_75t_L g1391 ( 
.A1(n_1385),
.A2(n_1311),
.B(n_1339),
.C(n_1345),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1358),
.B(n_1300),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1358),
.B(n_1373),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1373),
.B(n_1305),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1384),
.B(n_1353),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1387),
.B(n_1331),
.C(n_1337),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1384),
.B(n_1368),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1384),
.B(n_1353),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1372),
.A2(n_1329),
.B(n_1365),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1368),
.B(n_1376),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1368),
.B(n_1334),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1381),
.A2(n_1344),
.B1(n_1355),
.B2(n_1299),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1387),
.B(n_1351),
.C(n_1337),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1376),
.B(n_1308),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1325),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1382),
.B(n_1308),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1325),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1382),
.B(n_1336),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1375),
.B(n_1322),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1365),
.A2(n_1352),
.B(n_1338),
.Y(n_1410)
);

OAI21xp33_ASAP7_75t_L g1411 ( 
.A1(n_1370),
.A2(n_1351),
.B(n_1340),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1375),
.B(n_1330),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1367),
.B(n_1316),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1374),
.B(n_1314),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1363),
.B(n_1342),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1367),
.A2(n_1355),
.B1(n_1301),
.B2(n_1352),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1360),
.A2(n_1335),
.B1(n_1333),
.B2(n_1357),
.C(n_1321),
.Y(n_1417)
);

OR2x2_ASAP7_75t_SL g1418 ( 
.A(n_1362),
.B(n_1346),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1383),
.A2(n_1349),
.B(n_1356),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1363),
.B(n_1354),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1366),
.B(n_1354),
.Y(n_1421)
);

AOI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1360),
.A2(n_1321),
.B1(n_1348),
.B2(n_1347),
.C(n_1350),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1370),
.A2(n_1374),
.B(n_1359),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1371),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1361),
.A2(n_1321),
.B1(n_1348),
.B2(n_1347),
.C(n_1350),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1371),
.B(n_1341),
.Y(n_1426)
);

AND2x4_ASAP7_75t_SL g1427 ( 
.A(n_1401),
.B(n_1379),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1400),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1392),
.B(n_1377),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1389),
.B(n_1377),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1397),
.B(n_1400),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1424),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1424),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1420),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1399),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1421),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1426),
.B(n_1380),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1405),
.B(n_1380),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1404),
.B(n_1379),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1415),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1390),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1407),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1393),
.B(n_1386),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1399),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1418),
.B(n_1386),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1418),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1414),
.Y(n_1447)
);

NAND2x1p5_ASAP7_75t_L g1448 ( 
.A(n_1406),
.B(n_1362),
.Y(n_1448)
);

AND2x4_ASAP7_75t_SL g1449 ( 
.A(n_1395),
.B(n_1379),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1409),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1410),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1410),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1395),
.B(n_1398),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1412),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1408),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1423),
.B(n_1369),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1413),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1410),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1432),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1441),
.B(n_1423),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1449),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1433),
.Y(n_1462)
);

INVxp67_ASAP7_75t_SL g1463 ( 
.A(n_1456),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1433),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1431),
.B(n_1406),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1434),
.Y(n_1466)
);

INVx3_ASAP7_75t_SL g1467 ( 
.A(n_1445),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1431),
.B(n_1414),
.Y(n_1468)
);

NOR2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1455),
.B(n_1319),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1428),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1435),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1449),
.B(n_1427),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1434),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1437),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1448),
.B(n_1364),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1427),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1435),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1438),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1444),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1436),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1417),
.C(n_1396),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1440),
.B(n_1422),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1428),
.B(n_1403),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1439),
.B(n_1403),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1438),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_1439),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1443),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1443),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1487),
.B(n_1453),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1471),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1480),
.B(n_1450),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1478),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1459),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1482),
.B(n_1450),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1484),
.B(n_1454),
.Y(n_1496)
);

NAND4xp25_ASAP7_75t_L g1497 ( 
.A(n_1481),
.B(n_1391),
.C(n_1394),
.D(n_1236),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1460),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1469),
.B(n_1202),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1487),
.B(n_1439),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1472),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1471),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1472),
.B(n_1485),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1469),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1486),
.B(n_1429),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1474),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1463),
.A2(n_1411),
.B(n_1445),
.Y(n_1508)
);

NAND2xp67_ASAP7_75t_L g1509 ( 
.A(n_1477),
.B(n_1451),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1461),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1467),
.A2(n_1391),
.B1(n_1411),
.B2(n_1402),
.Y(n_1512)
);

AOI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1466),
.A2(n_1458),
.B(n_1452),
.Y(n_1513)
);

CKINVDCx8_ASAP7_75t_R g1514 ( 
.A(n_1485),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1488),
.B(n_1457),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1488),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1467),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1467),
.B(n_1447),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1483),
.B(n_1446),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_SL g1520 ( 
.A(n_1475),
.B(n_1461),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1430),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1509),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1500),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1521),
.B(n_1473),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1490),
.B(n_1483),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_1483),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1517),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1499),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1521),
.B(n_1473),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1514),
.Y(n_1532)
);

NAND2x1_ASAP7_75t_SL g1533 ( 
.A(n_1518),
.B(n_1470),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1497),
.B(n_1319),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1498),
.B(n_1462),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1518),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1510),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1494),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1504),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1493),
.B(n_1462),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1510),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1506),
.B(n_1464),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1507),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1504),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1497),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1501),
.B(n_1476),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1501),
.B(n_1476),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1503),
.B(n_1468),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1534),
.B(n_1512),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1531),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1536),
.B(n_1516),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1548),
.A2(n_1512),
.B(n_1532),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1531),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1532),
.B(n_1231),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1523),
.B(n_1503),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1514),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1527),
.B(n_1492),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1539),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1539),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1537),
.Y(n_1565)
);

AOI21xp33_ASAP7_75t_L g1566 ( 
.A1(n_1535),
.A2(n_1502),
.B(n_1491),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1532),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1540),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1532),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1540),
.Y(n_1570)
);

XNOR2x1_ASAP7_75t_L g1571 ( 
.A(n_1546),
.B(n_1551),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1547),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1550),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1547),
.Y(n_1574)
);

NAND2x1_ASAP7_75t_SL g1575 ( 
.A(n_1541),
.B(n_1519),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1535),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1499),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1534),
.A2(n_1519),
.B1(n_1508),
.B2(n_1416),
.Y(n_1578)
);

OAI221xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1537),
.A2(n_1506),
.B1(n_1515),
.B2(n_1446),
.C(n_1419),
.Y(n_1579)
);

NOR2x1p5_ASAP7_75t_SL g1580 ( 
.A(n_1567),
.B(n_1543),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1573),
.B(n_1523),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1565),
.Y(n_1582)
);

NOR3xp33_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1528),
.C(n_1536),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1561),
.B(n_1356),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1569),
.B(n_1538),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1571),
.B(n_1546),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1565),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1555),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1559),
.B(n_1544),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1560),
.B(n_1553),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1553),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1554),
.A2(n_1544),
.B(n_1542),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1559),
.B(n_1550),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1571),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1558),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1562),
.B(n_1524),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1552),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1556),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1563),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1586),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1594),
.A2(n_1592),
.B(n_1554),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1583),
.A2(n_1578),
.B1(n_1577),
.B2(n_1522),
.Y(n_1602)
);

AND4x1_ASAP7_75t_L g1603 ( 
.A(n_1584),
.B(n_1577),
.C(n_1552),
.D(n_1576),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1589),
.A2(n_1579),
.B(n_1566),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1596),
.A2(n_1528),
.B1(n_1529),
.B2(n_1522),
.Y(n_1605)
);

OAI31xp33_ASAP7_75t_L g1606 ( 
.A1(n_1589),
.A2(n_1529),
.A3(n_1522),
.B(n_1519),
.Y(n_1606)
);

AOI21xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1585),
.A2(n_1499),
.B(n_1541),
.Y(n_1607)
);

CKINVDCx16_ASAP7_75t_R g1608 ( 
.A(n_1593),
.Y(n_1608)
);

NOR2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1596),
.B(n_1528),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1582),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1597),
.B(n_1564),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_L g1612 ( 
.A(n_1601),
.B(n_1587),
.Y(n_1612)
);

NAND3xp33_ASAP7_75t_SL g1613 ( 
.A(n_1604),
.B(n_1593),
.C(n_1591),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1608),
.B(n_1590),
.Y(n_1614)
);

INVxp33_ASAP7_75t_L g1615 ( 
.A(n_1602),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1600),
.B(n_1598),
.C(n_1597),
.Y(n_1616)
);

XNOR2x2_ASAP7_75t_L g1617 ( 
.A(n_1610),
.B(n_1591),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1609),
.B(n_1588),
.Y(n_1618)
);

NOR3xp33_ASAP7_75t_L g1619 ( 
.A(n_1600),
.B(n_1528),
.C(n_1595),
.Y(n_1619)
);

NOR3xp33_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1599),
.C(n_1570),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1607),
.B(n_1611),
.C(n_1572),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1622)
);

OAI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1616),
.A2(n_1575),
.B(n_1606),
.C(n_1533),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_L g1624 ( 
.A(n_1613),
.B(n_1218),
.C(n_1568),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1614),
.B(n_1603),
.Y(n_1625)
);

AOI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1621),
.A2(n_1574),
.B(n_1580),
.C(n_1541),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1622),
.B(n_1581),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1625),
.A2(n_1615),
.B1(n_1620),
.B2(n_1619),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1623),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1626),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1624),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1622),
.B(n_1581),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1627),
.Y(n_1633)
);

NAND4xp75_ASAP7_75t_L g1634 ( 
.A(n_1628),
.B(n_1618),
.C(n_1580),
.D(n_1617),
.Y(n_1634)
);

AOI32xp33_ASAP7_75t_L g1635 ( 
.A1(n_1629),
.A2(n_1590),
.A3(n_1541),
.B1(n_1525),
.B2(n_1529),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1632),
.Y(n_1636)
);

NOR2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1630),
.B(n_1209),
.Y(n_1637)
);

NOR2xp67_ASAP7_75t_L g1638 ( 
.A(n_1636),
.B(n_1236),
.Y(n_1638)
);

NAND2x1p5_ASAP7_75t_L g1639 ( 
.A(n_1633),
.B(n_1631),
.Y(n_1639)
);

NAND4xp75_ASAP7_75t_L g1640 ( 
.A(n_1634),
.B(n_1525),
.C(n_1526),
.D(n_1543),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1639),
.B(n_1543),
.Y(n_1641)
);

NOR2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1641),
.B(n_1640),
.Y(n_1642)
);

OAI22x1_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1637),
.B1(n_1638),
.B2(n_1635),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1642),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1644),
.A2(n_1530),
.B1(n_1524),
.B2(n_1545),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1643),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1646),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1647),
.Y(n_1648)
);

AOI322xp5_ASAP7_75t_L g1649 ( 
.A1(n_1648),
.A2(n_1645),
.A3(n_1549),
.B1(n_1519),
.B2(n_1542),
.C1(n_1513),
.C2(n_1526),
.Y(n_1649)
);

OAI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1649),
.A2(n_1533),
.B1(n_1268),
.B2(n_1549),
.C(n_1231),
.Y(n_1650)
);

AOI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1270),
.B(n_1259),
.C(n_1549),
.Y(n_1651)
);


endmodule