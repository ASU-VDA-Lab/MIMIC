module fake_jpeg_8204_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_9),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_43),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_18),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_22),
.B1(n_21),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_58),
.B1(n_63),
.B2(n_66),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_33),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_23),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_22),
.B1(n_19),
.B2(n_31),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_38),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_73),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_24),
.B1(n_29),
.B2(n_25),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_96),
.B(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_80),
.Y(n_106)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_88),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_48),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_42),
.C(n_28),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_23),
.B1(n_31),
.B2(n_16),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_23),
.B1(n_31),
.B2(n_27),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_107),
.A2(n_18),
.B(n_28),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_69),
.B1(n_52),
.B2(n_30),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_112),
.B1(n_120),
.B2(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_48),
.B1(n_61),
.B2(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_80),
.B1(n_98),
.B2(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_67),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_48),
.B1(n_69),
.B2(n_52),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_93),
.B1(n_77),
.B2(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_87),
.B1(n_82),
.B2(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_131),
.B(n_132),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_100),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_133),
.B(n_140),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_137),
.B1(n_148),
.B2(n_118),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_89),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_138),
.C(n_101),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_81),
.B1(n_68),
.B2(n_94),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_81),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_146),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_143),
.B(n_144),
.Y(n_193)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_88),
.B1(n_78),
.B2(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_113),
.B1(n_116),
.B2(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_19),
.B1(n_16),
.B2(n_27),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_151),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_17),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_158),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_19),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_109),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_42),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_108),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_18),
.B(n_28),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_116),
.B(n_125),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_17),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_42),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_165),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_163),
.A2(n_168),
.B1(n_177),
.B2(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_108),
.B1(n_115),
.B2(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_183),
.B1(n_192),
.B2(n_2),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_175),
.B(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_182),
.C(n_179),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_101),
.B(n_109),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_108),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_108),
.B1(n_113),
.B2(n_103),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_189),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_4),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_103),
.B1(n_18),
.B2(n_28),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_18),
.B1(n_28),
.B2(n_30),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_104),
.C(n_28),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_104),
.B1(n_30),
.B2(n_28),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_18),
.B1(n_104),
.B2(n_10),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_138),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_203),
.C(n_206),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_194),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_172),
.B1(n_193),
.B2(n_163),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_130),
.B(n_156),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_208),
.B(n_217),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_142),
.C(n_152),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_142),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_192),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_148),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_210),
.B(n_213),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_8),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_221),
.B1(n_171),
.B2(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_166),
.B(n_8),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_178),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_161),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_11),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_225),
.B(n_238),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_186),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_199),
.C(n_210),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_231),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_195),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_234),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_189),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_173),
.B1(n_164),
.B2(n_165),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_205),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_242),
.B1(n_218),
.B2(n_213),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_199),
.B(n_214),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_173),
.B1(n_164),
.B2(n_184),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_221),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_12),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_248),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_12),
.C(n_14),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_249),
.B(n_252),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_228),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_209),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_211),
.B(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_211),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_266),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_232),
.C(n_231),
.Y(n_275)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_219),
.B1(n_222),
.B2(n_7),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_236),
.B1(n_248),
.B2(n_11),
.Y(n_282)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_232),
.B1(n_234),
.B2(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_224),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_278),
.C(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_283),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_227),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_265),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_246),
.C(n_230),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_11),
.Y(n_283)
);

XOR2x1_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_250),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_293),
.B1(n_13),
.B2(n_15),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_287),
.B(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_257),
.B(n_264),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_261),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.C(n_275),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_259),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_253),
.B(n_256),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_258),
.B(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_276),
.B1(n_272),
.B2(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_273),
.B1(n_271),
.B2(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_268),
.B1(n_274),
.B2(n_278),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_15),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_285),
.C(n_15),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_289),
.B(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_294),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_304),
.C(n_300),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_306),
.B(n_307),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_308),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_319),
.B(n_310),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_312),
.A2(n_311),
.B1(n_277),
.B2(n_309),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_318),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_321),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_315),
.Y(n_326)
);


endmodule