module fake_jpeg_23835_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_35),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_12),
.B1(n_18),
.B2(n_16),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_16),
.B1(n_19),
.B2(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_12),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_44),
.B1(n_29),
.B2(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_45),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_29),
.Y(n_47)
);

OAI22x1_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_11),
.B1(n_19),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_35),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_44),
.C(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_53),
.B1(n_39),
.B2(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.C(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_45),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_52),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_60),
.B1(n_63),
.B2(n_50),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_70),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_44),
.Y(n_74)
);


endmodule