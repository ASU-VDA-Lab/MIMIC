module fake_aes_7753_n_730 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_730);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_730;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_49), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_33), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_10), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_5), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_18), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_1), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_50), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_78), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_4), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_8), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_47), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_26), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_41), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_25), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_4), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_31), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_24), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_56), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_57), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_46), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_61), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_60), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_63), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_22), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_16), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_14), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_1), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_9), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_18), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_58), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_42), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_34), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_36), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_69), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_51), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_43), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_128), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_86), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_96), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_104), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
NOR2x1_ASAP7_75t_L g142 ( .A(n_121), .B(n_37), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_117), .B(n_0), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_120), .B(n_123), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_87), .B(n_0), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_93), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_106), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_101), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_90), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_100), .B(n_2), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_113), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_89), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_84), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_101), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_107), .B(n_6), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_108), .B(n_7), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_109), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_92), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_111), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_129), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_110), .B(n_11), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_91), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_111), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_116), .Y(n_173) );
NOR2x1_ASAP7_75t_L g174 ( .A(n_116), .B(n_44), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_98), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_102), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_135), .B(n_118), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_176), .B(n_118), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_147), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_176), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_176), .B(n_131), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_176), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_171), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_171), .B(n_140), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_159), .B(n_131), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_147), .B(n_119), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_149), .B(n_119), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_147), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_173), .B(n_122), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_150), .B(n_122), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_139), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_140), .B(n_130), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_134), .Y(n_207) );
INVx8_ASAP7_75t_L g208 ( .A(n_169), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_125), .B1(n_130), .B2(n_126), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_173), .B(n_112), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_173), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_143), .B(n_125), .C(n_126), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_159), .B(n_105), .Y(n_216) );
XOR2xp5_ASAP7_75t_L g217 ( .A(n_160), .B(n_11), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_157), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_138), .B(n_105), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_132), .B(n_112), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_152), .B(n_103), .Y(n_223) );
BUFx4_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_157), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_163), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_163), .Y(n_229) );
NOR2xp67_ASAP7_75t_L g230 ( .A(n_153), .B(n_98), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_132), .B(n_124), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_154), .B(n_124), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_175), .B(n_115), .Y(n_237) );
NAND3x1_ASAP7_75t_L g238 ( .A(n_151), .B(n_99), .C(n_103), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_167), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_167), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_155), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_197), .A2(n_156), .B(n_172), .C(n_168), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_203), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_201), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_190), .A2(n_162), .B1(n_158), .B2(n_166), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_243), .B(n_170), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_223), .B(n_145), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
NOR2x1p5_ASAP7_75t_L g253 ( .A(n_207), .B(n_134), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_214), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_223), .B(n_145), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_198), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_243), .B(n_165), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_178), .B(n_145), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_178), .A2(n_162), .B1(n_174), .B2(n_142), .Y(n_263) );
AOI22xp5_ASAP7_75t_SL g264 ( .A1(n_217), .A2(n_160), .B1(n_127), .B2(n_115), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
NOR3xp33_ASAP7_75t_SL g266 ( .A(n_207), .B(n_114), .C(n_99), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_197), .A2(n_114), .B(n_97), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_198), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_210), .B(n_12), .C(n_13), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_208), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_208), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_178), .B(n_12), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_195), .B(n_15), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_236), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_195), .B(n_16), .Y(n_276) );
NOR2x1p5_ASAP7_75t_SL g277 ( .A(n_193), .B(n_81), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_182), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_211), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_181), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_211), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_211), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_187), .B(n_53), .Y(n_283) );
NOR3xp33_ASAP7_75t_SL g284 ( .A(n_221), .B(n_17), .C(n_20), .Y(n_284) );
OR2x6_ASAP7_75t_L g285 ( .A(n_208), .B(n_17), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_181), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_196), .B(n_21), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_182), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_208), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_227), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_195), .B(n_21), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_197), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_195), .B(n_22), .Y(n_295) );
INVx5_ASAP7_75t_L g296 ( .A(n_211), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_236), .Y(n_297) );
AO22x1_ASAP7_75t_L g298 ( .A1(n_187), .A2(n_23), .B1(n_27), .B2(n_28), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_191), .B(n_29), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_196), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_208), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_228), .Y(n_302) );
INVx5_ASAP7_75t_L g303 ( .A(n_211), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_217), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_200), .B(n_30), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_222), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_224), .Y(n_307) );
NAND3xp33_ASAP7_75t_SL g308 ( .A(n_204), .B(n_32), .C(n_35), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_200), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_179), .B(n_38), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_179), .B(n_39), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_216), .B(n_40), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_235), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_228), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_246), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_258), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_271), .B(n_183), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_258), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_245), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_274), .A2(n_238), .B1(n_233), .B2(n_215), .Y(n_322) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_271), .B(n_183), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_256), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g325 ( .A1(n_300), .A2(n_230), .B1(n_237), .B2(n_222), .C1(n_231), .C2(n_213), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_274), .B(n_185), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_274), .B(n_185), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_295), .A2(n_237), .B1(n_231), .B2(n_222), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_250), .B(n_231), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_294), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_287), .B(n_237), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_297), .B(n_224), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_295), .A2(n_242), .B1(n_184), .B2(n_234), .Y(n_334) );
INVx5_ASAP7_75t_L g335 ( .A(n_285), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_295), .A2(n_238), .B1(n_242), .B2(n_228), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_307), .B(n_234), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_289), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_244), .A2(n_192), .B(n_232), .C(n_225), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_244), .A2(n_192), .B(n_232), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_285), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_248), .B(n_234), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_287), .B(n_188), .Y(n_343) );
BUFx8_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_261), .A2(n_188), .B(n_225), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_309), .B(n_186), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_275), .A2(n_186), .B1(n_220), .B2(n_219), .C(n_218), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_292), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
INVx5_ASAP7_75t_L g350 ( .A(n_285), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_260), .Y(n_351) );
NOR2xp67_ASAP7_75t_L g352 ( .A(n_263), .B(n_48), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_262), .B(n_189), .Y(n_353) );
INVx5_ASAP7_75t_L g354 ( .A(n_289), .Y(n_354) );
INVx5_ASAP7_75t_L g355 ( .A(n_302), .Y(n_355) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_306), .B(n_276), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_272), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_265), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_262), .B(n_241), .Y(n_359) );
AND2x6_ASAP7_75t_L g360 ( .A(n_269), .B(n_189), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_302), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_302), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_311), .B(n_312), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_273), .B(n_235), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_315), .Y(n_366) );
INVx8_ASAP7_75t_L g367 ( .A(n_272), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_270), .A2(n_241), .B(n_220), .C(n_219), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_290), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_315), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_290), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_322), .A2(n_266), .B1(n_284), .B2(n_293), .C(n_251), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_342), .A2(n_253), .B1(n_301), .B2(n_291), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_358), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_329), .A2(n_301), .B1(n_255), .B2(n_251), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_317), .A2(n_255), .B1(n_280), .B2(n_286), .Y(n_376) );
NOR3xp33_ASAP7_75t_SL g377 ( .A(n_368), .B(n_308), .C(n_299), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_316), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_319), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_331), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_331), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_330), .B(n_305), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_344), .Y(n_384) );
INVx4_ASAP7_75t_L g385 ( .A(n_319), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_267), .B(n_313), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_332), .B(n_278), .Y(n_387) );
NAND3xp33_ASAP7_75t_SL g388 ( .A(n_325), .B(n_283), .C(n_252), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_339), .A2(n_218), .B(n_180), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_320), .B(n_304), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_333), .A2(n_278), .B1(n_288), .B2(n_254), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_319), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_324), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_344), .A2(n_288), .B1(n_180), .B2(n_194), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_344), .A2(n_209), .B1(n_194), .B2(n_199), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_319), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_321), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_319), .B(n_277), .Y(n_400) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_341), .B(n_298), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_321), .B(n_264), .Y(n_402) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_336), .A2(n_209), .B(n_199), .C(n_202), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_356), .A2(n_332), .B1(n_335), .B2(n_350), .Y(n_404) );
AND2x6_ASAP7_75t_L g405 ( .A(n_327), .B(n_259), .Y(n_405) );
O2A1O1Ixp5_ASAP7_75t_SL g406 ( .A1(n_340), .A2(n_202), .B(n_212), .C(n_277), .Y(n_406) );
OR2x6_ASAP7_75t_L g407 ( .A(n_385), .B(n_367), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_394), .A2(n_212), .A3(n_337), .B1(n_239), .B2(n_229), .B3(n_226), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_372), .A2(n_356), .B1(n_335), .B2(n_350), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_386), .A2(n_368), .B(n_363), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_380), .B(n_335), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_372), .A2(n_350), .B1(n_335), .B2(n_352), .Y(n_414) );
INVx4_ASAP7_75t_SL g415 ( .A(n_405), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_378), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_405), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_402), .A2(n_346), .B1(n_353), .B2(n_334), .C(n_357), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_375), .A2(n_350), .B1(n_335), .B2(n_367), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_384), .A2(n_350), .B1(n_367), .B2(n_369), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_377), .B(n_365), .C(n_363), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_381), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_383), .A2(n_388), .B(n_386), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_367), .B1(n_327), .B2(n_328), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_373), .A2(n_376), .B(n_378), .C(n_384), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_405), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_391), .A2(n_371), .B1(n_369), .B2(n_327), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_328), .B1(n_343), .B2(n_359), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
AOI222xp33_ASAP7_75t_L g433 ( .A1(n_399), .A2(n_343), .B1(n_347), .B2(n_328), .C1(n_349), .C2(n_338), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_401), .A2(n_323), .B1(n_318), .B2(n_326), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_388), .A2(n_338), .B1(n_349), .B2(n_364), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_410), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_410), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_421), .A2(n_377), .B(n_401), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_416), .B(n_394), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_423), .B(n_406), .C(n_403), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_433), .A2(n_401), .B1(n_387), .B2(n_374), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_428), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_428), .Y(n_445) );
OAI211xp5_ASAP7_75t_SL g446 ( .A1(n_429), .A2(n_392), .B(n_404), .C(n_395), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_430), .A2(n_374), .B1(n_389), .B2(n_393), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_418), .B(n_395), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_422), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_425), .A2(n_379), .B(n_393), .C(n_387), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_422), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_426), .A2(n_387), .B1(n_403), .B2(n_389), .C(n_396), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_424), .B(n_390), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_436), .B(n_390), .Y(n_455) );
NAND2xp33_ASAP7_75t_R g456 ( .A(n_407), .B(n_400), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_427), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_431), .Y(n_461) );
NAND2xp33_ASAP7_75t_R g462 ( .A(n_407), .B(n_400), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_427), .B(n_390), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_436), .B(n_390), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_435), .A2(n_345), .B1(n_397), .B2(n_379), .C(n_338), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_413), .B(n_379), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_413), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_430), .B(n_405), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_411), .Y(n_471) );
AOI211xp5_ASAP7_75t_L g472 ( .A1(n_419), .A2(n_400), .B(n_326), .C(n_348), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_411), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_454), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_454), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_453), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_458), .B(n_411), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_437), .B(n_432), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_443), .B(n_412), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_443), .B(n_412), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_440), .B(n_425), .Y(n_482) );
AND2x4_ASAP7_75t_SL g483 ( .A(n_467), .B(n_407), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_461), .B(n_415), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_449), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_469), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_451), .B(n_432), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_467), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_451), .B(n_431), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_457), .B(n_431), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_457), .B(n_431), .Y(n_492) );
INVx4_ASAP7_75t_L g493 ( .A(n_461), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_460), .B(n_431), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_460), .B(n_434), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_464), .B(n_431), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_447), .A2(n_409), .A3(n_421), .B(n_414), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_464), .B(n_415), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_444), .B(n_417), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_438), .B(n_415), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_455), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_438), .B(n_415), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_448), .B(n_420), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_441), .A2(n_406), .B(n_400), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_444), .B(n_417), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_468), .B(n_415), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_439), .A2(n_417), .B1(n_407), .B2(n_385), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_441), .B(n_365), .C(n_398), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_468), .B(n_407), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g511 ( .A1(n_442), .A2(n_385), .B1(n_398), .B2(n_323), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_445), .B(n_398), .Y(n_512) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_472), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_446), .A2(n_408), .B1(n_349), .B2(n_385), .C(n_398), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_445), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_469), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_455), .Y(n_517) );
OR2x2_ASAP7_75t_SL g518 ( .A(n_470), .B(n_348), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_471), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_463), .B(n_382), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_463), .B(n_382), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_465), .B(n_382), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_465), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_442), .A2(n_405), .B1(n_365), .B2(n_348), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_472), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_502), .B(n_473), .Y(n_526) );
OA222x2_ASAP7_75t_L g527 ( .A1(n_512), .A2(n_456), .B1(n_462), .B2(n_461), .C1(n_473), .C2(n_471), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_476), .B(n_450), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_502), .B(n_452), .Y(n_530) );
NAND2xp33_ASAP7_75t_SL g531 ( .A(n_511), .B(n_405), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_517), .B(n_466), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_517), .B(n_365), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_523), .B(n_226), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_495), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_523), .B(n_239), .Y(n_536) );
AOI33xp33_ASAP7_75t_L g537 ( .A1(n_524), .A2(n_193), .A3(n_205), .B1(n_206), .B2(n_229), .B3(n_370), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
NAND2xp33_ASAP7_75t_R g539 ( .A(n_499), .B(n_52), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_482), .B(n_405), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_521), .B(n_206), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_485), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_521), .B(n_205), .Y(n_544) );
AOI33xp33_ASAP7_75t_L g545 ( .A1(n_508), .A2(n_370), .A3(n_366), .B1(n_361), .B2(n_257), .B3(n_268), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_489), .B(n_240), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_504), .B(n_354), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_525), .A2(n_318), .B1(n_364), .B2(n_362), .C(n_354), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_519), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_522), .B(n_240), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_489), .B(n_366), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_513), .B(n_354), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_513), .A2(n_355), .B1(n_354), .B2(n_364), .Y(n_555) );
NOR2x1_ASAP7_75t_SL g556 ( .A(n_512), .B(n_355), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_519), .Y(n_557) );
AOI22x1_ASAP7_75t_L g558 ( .A1(n_525), .A2(n_361), .B1(n_362), .B2(n_240), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_480), .B(n_362), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_522), .B(n_240), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_477), .B(n_240), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_483), .B(n_354), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_477), .B(n_235), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_480), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_515), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_474), .B(n_235), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_509), .A2(n_355), .B(n_296), .Y(n_567) );
NAND2xp33_ASAP7_75t_SL g568 ( .A(n_511), .B(n_360), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_474), .B(n_54), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_475), .B(n_519), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_483), .B(n_355), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_475), .B(n_55), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_486), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_481), .B(n_355), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_484), .B(n_492), .Y(n_576) );
NOR4xp25_ASAP7_75t_SL g577 ( .A(n_514), .B(n_59), .C(n_62), .D(n_64), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_509), .B(n_65), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_483), .B(n_68), .Y(n_579) );
NAND2x1_ASAP7_75t_L g580 ( .A(n_493), .B(n_360), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_478), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_490), .B(n_70), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_510), .B(n_360), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_508), .Y(n_584) );
AO221x1_ASAP7_75t_L g585 ( .A1(n_527), .A2(n_529), .B1(n_535), .B2(n_531), .C(n_539), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_529), .Y(n_586) );
NOR2xp67_ASAP7_75t_L g587 ( .A(n_584), .B(n_493), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_541), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_541), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_564), .B(n_497), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_584), .A2(n_510), .B1(n_499), .B2(n_514), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_565), .A2(n_505), .B(n_491), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_547), .A2(n_530), .B1(n_568), .B2(n_531), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_572), .A2(n_496), .B1(n_478), .B2(n_488), .Y(n_594) );
NOR2xp33_ASAP7_75t_R g595 ( .A(n_568), .B(n_496), .Y(n_595) );
AOI33xp33_ASAP7_75t_L g596 ( .A1(n_530), .A2(n_490), .A3(n_494), .B1(n_492), .B2(n_491), .B3(n_497), .Y(n_596) );
AOI32xp33_ASAP7_75t_L g597 ( .A1(n_578), .A2(n_501), .A3(n_503), .B1(n_507), .B2(n_506), .Y(n_597) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_554), .A2(n_505), .B(n_498), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_572), .A2(n_488), .B1(n_506), .B2(n_500), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_580), .B(n_493), .Y(n_600) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_556), .Y(n_601) );
AOI32xp33_ASAP7_75t_L g602 ( .A1(n_579), .A2(n_501), .A3(n_503), .B1(n_507), .B2(n_500), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_556), .Y(n_603) );
OAI32xp33_ASAP7_75t_L g604 ( .A1(n_528), .A2(n_493), .A3(n_520), .B1(n_516), .B2(n_486), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_540), .A2(n_498), .B1(n_520), .B2(n_516), .C(n_518), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_570), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_528), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_581), .B(n_516), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_559), .A2(n_518), .B1(n_303), .B2(n_296), .C(n_268), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_538), .Y(n_611) );
INVxp33_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_576), .B(n_484), .Y(n_613) );
NAND3xp33_ASAP7_75t_SL g614 ( .A(n_545), .B(n_71), .C(n_74), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_532), .B(n_484), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_580), .A2(n_303), .B(n_296), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_550), .B(n_75), .Y(n_617) );
NAND2x1_ASAP7_75t_L g618 ( .A(n_550), .B(n_360), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_549), .A2(n_247), .B(n_314), .C(n_257), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_548), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_526), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_576), .B(n_526), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_533), .B(n_76), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_557), .B(n_77), .Y(n_626) );
AOI211x1_ASAP7_75t_SL g627 ( .A1(n_555), .A2(n_79), .B(n_80), .C(n_247), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_R g628 ( .A1(n_574), .A2(n_249), .B(n_314), .C(n_282), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_557), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_575), .B(n_249), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_575), .B(n_282), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_532), .B(n_360), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_573), .B(n_279), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_571), .A2(n_296), .B1(n_303), .B2(n_279), .C(n_259), .Y(n_634) );
AOI211x1_ASAP7_75t_L g635 ( .A1(n_569), .A2(n_360), .B(n_296), .C(n_303), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_566), .Y(n_636) );
NOR2xp33_ASAP7_75t_R g637 ( .A(n_603), .B(n_582), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_623), .Y(n_638) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_601), .Y(n_639) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_612), .A2(n_566), .B(n_569), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g641 ( .A(n_595), .B(n_537), .C(n_577), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_586), .Y(n_642) );
XNOR2xp5_ASAP7_75t_L g643 ( .A(n_624), .B(n_593), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_614), .B(n_567), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_597), .A2(n_582), .B(n_533), .C(n_544), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_606), .B(n_563), .Y(n_646) );
XOR2x2_ASAP7_75t_L g647 ( .A(n_587), .B(n_583), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_608), .B(n_563), .Y(n_648) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_586), .B(n_546), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_607), .B(n_561), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_590), .B(n_561), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_605), .A2(n_542), .A3(n_544), .B(n_551), .Y(n_652) );
NAND2xp33_ASAP7_75t_R g653 ( .A(n_585), .B(n_573), .Y(n_653) );
NOR3xp33_ASAP7_75t_SL g654 ( .A(n_598), .B(n_552), .C(n_558), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_615), .B(n_542), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_611), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_629), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_609), .B(n_560), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_613), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_588), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_636), .B(n_560), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_620), .Y(n_662) );
XNOR2x2_ASAP7_75t_L g663 ( .A(n_635), .B(n_599), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_600), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_621), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_622), .B(n_551), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_596), .B(n_536), .Y(n_667) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_598), .A2(n_536), .B(n_534), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_589), .B(n_534), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_633), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_594), .A2(n_558), .B1(n_303), .B2(n_279), .C1(n_281), .C2(n_310), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_610), .Y(n_672) );
NAND2xp33_ASAP7_75t_L g673 ( .A(n_602), .B(n_279), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_639), .Y(n_674) );
HAxp5_ASAP7_75t_SL g675 ( .A(n_653), .B(n_591), .CON(n_675), .SN(n_675) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_664), .B(n_618), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_652), .A2(n_592), .B1(n_594), .B2(n_600), .C(n_599), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_672), .A2(n_673), .B(n_667), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g679 ( .A1(n_639), .A2(n_625), .A3(n_632), .B1(n_634), .B2(n_628), .Y(n_679) );
INVxp33_ASAP7_75t_L g680 ( .A(n_664), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_657), .B(n_632), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g682 ( .A(n_643), .B(n_627), .Y(n_682) );
NAND4xp75_ASAP7_75t_L g683 ( .A(n_644), .B(n_616), .C(n_604), .D(n_619), .Y(n_683) );
OAI21xp33_ASAP7_75t_SL g684 ( .A1(n_649), .A2(n_617), .B(n_626), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_656), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_672), .B(n_630), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_645), .A2(n_631), .B(n_279), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_668), .A2(n_654), .B(n_642), .C(n_640), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_637), .B(n_259), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_670), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_662), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_665), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_670), .B(n_259), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_646), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_660), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_654), .A2(n_281), .B(n_310), .C(n_641), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_696), .B(n_678), .C(n_688), .Y(n_697) );
INVxp33_ASAP7_75t_SL g698 ( .A(n_682), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_696), .B(n_641), .C(n_671), .D(n_655), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_690), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_690), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_679), .A2(n_648), .B(n_669), .C(n_651), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_686), .B(n_638), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_680), .Y(n_704) );
AND2x2_ASAP7_75t_SL g705 ( .A(n_675), .B(n_650), .Y(n_705) );
XNOR2x1_ASAP7_75t_L g706 ( .A(n_676), .B(n_663), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_674), .Y(n_707) );
INVxp67_ASAP7_75t_L g708 ( .A(n_693), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_680), .A2(n_647), .B(n_659), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_689), .A2(n_658), .B(n_666), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_677), .A2(n_661), .B1(n_281), .B2(n_310), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_687), .A2(n_310), .B(n_684), .C(n_692), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_685), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_683), .B(n_691), .C(n_695), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_681), .A2(n_678), .B(n_696), .C(n_679), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_694), .B(n_680), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_705), .A2(n_706), .B(n_698), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_707), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_705), .A2(n_697), .B1(n_699), .B2(n_711), .Y(n_719) );
OR3x1_ASAP7_75t_L g720 ( .A(n_700), .B(n_701), .C(n_715), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_704), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_717), .A2(n_712), .B1(n_714), .B2(n_709), .C(n_702), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_721), .Y(n_723) );
OAI222xp33_ASAP7_75t_L g724 ( .A1(n_719), .A2(n_716), .B1(n_708), .B2(n_710), .C1(n_703), .C2(n_713), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_722), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_725), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_726), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_720), .B1(n_718), .B2(n_708), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_727), .B(n_724), .Y(n_730) );
endmodule