module real_aes_350_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_0), .B(n_136), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_1), .A2(n_145), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_2), .B(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_3), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_4), .B(n_152), .Y(n_215) );
INVx1_ASAP7_75t_L g143 ( .A(n_5), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_6), .B(n_152), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_7), .B(n_156), .Y(n_480) );
INVx1_ASAP7_75t_L g514 ( .A(n_8), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g816 ( .A(n_9), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_10), .Y(n_552) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_11), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_13), .A2(n_25), .B1(n_136), .B2(n_145), .C(n_232), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_14), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_15), .B(n_136), .Y(n_135) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_16), .A2(n_131), .B(n_134), .Y(n_130) );
INVx1_ASAP7_75t_L g489 ( .A(n_17), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_18), .B(n_170), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_19), .B(n_152), .Y(n_179) );
AO21x1_ASAP7_75t_L g210 ( .A1(n_20), .A2(n_136), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g118 ( .A(n_21), .Y(n_118) );
INVx1_ASAP7_75t_L g487 ( .A(n_22), .Y(n_487) );
INVx1_ASAP7_75t_SL g497 ( .A(n_23), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_24), .B(n_137), .Y(n_580) );
NAND2x1_ASAP7_75t_L g201 ( .A(n_26), .B(n_152), .Y(n_201) );
AOI33xp33_ASAP7_75t_L g526 ( .A1(n_27), .A2(n_51), .A3(n_464), .B1(n_469), .B2(n_527), .B3(n_528), .Y(n_526) );
NAND2x1_ASAP7_75t_L g189 ( .A(n_28), .B(n_154), .Y(n_189) );
INVx1_ASAP7_75t_L g546 ( .A(n_29), .Y(n_546) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_30), .A2(n_86), .B(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g157 ( .A(n_30), .B(n_86), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_31), .B(n_472), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_32), .B(n_154), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_33), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_34), .B(n_154), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_35), .A2(n_145), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g142 ( .A(n_36), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g146 ( .A(n_36), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g463 ( .A(n_36), .Y(n_463) );
OR2x6_ASAP7_75t_L g116 ( .A(n_37), .B(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_38), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_39), .B(n_136), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_40), .B(n_472), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_41), .A2(n_156), .B1(n_163), .B2(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_42), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_43), .B(n_137), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_44), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_45), .B(n_154), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_46), .B(n_131), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_47), .B(n_137), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_48), .A2(n_145), .B(n_188), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_49), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_50), .B(n_154), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_52), .B(n_137), .Y(n_538) );
INVx1_ASAP7_75t_L g139 ( .A(n_53), .Y(n_139) );
INVx1_ASAP7_75t_L g149 ( .A(n_53), .Y(n_149) );
AND2x2_ASAP7_75t_L g539 ( .A(n_54), .B(n_170), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_55), .A2(n_72), .B1(n_461), .B2(n_472), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_56), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_57), .B(n_152), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_58), .B(n_163), .Y(n_554) );
AOI21xp5_ASAP7_75t_SL g460 ( .A1(n_59), .A2(n_461), .B(n_466), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_60), .A2(n_145), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g483 ( .A(n_61), .Y(n_483) );
AO21x1_ASAP7_75t_L g212 ( .A1(n_62), .A2(n_145), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_63), .B(n_136), .Y(n_165) );
INVx1_ASAP7_75t_L g537 ( .A(n_64), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_65), .B(n_136), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_67), .A2(n_461), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g225 ( .A(n_68), .B(n_171), .Y(n_225) );
INVx1_ASAP7_75t_L g141 ( .A(n_69), .Y(n_141) );
INVx1_ASAP7_75t_L g147 ( .A(n_69), .Y(n_147) );
AND2x2_ASAP7_75t_L g193 ( .A(n_70), .B(n_162), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_71), .B(n_472), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_73), .A2(n_785), .B1(n_789), .B2(n_791), .Y(n_788) );
OAI22xp5_ASAP7_75t_SL g802 ( .A1(n_74), .A2(n_84), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_74), .Y(n_803) );
AND2x2_ASAP7_75t_L g499 ( .A(n_75), .B(n_162), .Y(n_499) );
INVx1_ASAP7_75t_L g484 ( .A(n_76), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_77), .A2(n_461), .B(n_496), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_78), .A2(n_461), .B(n_521), .C(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g119 ( .A(n_79), .Y(n_119) );
AND2x2_ASAP7_75t_L g161 ( .A(n_80), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_81), .B(n_136), .Y(n_181) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_82), .B(n_162), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_83), .A2(n_461), .B1(n_524), .B2(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g804 ( .A(n_84), .Y(n_804) );
AND2x2_ASAP7_75t_L g211 ( .A(n_85), .B(n_156), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_87), .B(n_154), .Y(n_180) );
AND2x2_ASAP7_75t_L g205 ( .A(n_88), .B(n_162), .Y(n_205) );
INVx1_ASAP7_75t_L g467 ( .A(n_89), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_90), .B(n_152), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_91), .A2(n_145), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_92), .B(n_154), .Y(n_233) );
AND2x2_ASAP7_75t_L g530 ( .A(n_93), .B(n_162), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_94), .A2(n_95), .B1(n_786), .B2(n_787), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_94), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_95), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_96), .B(n_152), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_97), .A2(n_544), .B(n_545), .C(n_547), .Y(n_543) );
BUFx2_ASAP7_75t_L g106 ( .A(n_98), .Y(n_106) );
BUFx2_ASAP7_75t_SL g797 ( .A(n_98), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_99), .A2(n_145), .B(n_150), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_100), .B(n_137), .Y(n_470) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_810), .B(n_817), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_121), .B(n_795), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_108), .A2(n_799), .B(n_807), .Y(n_798) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_120), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g809 ( .A(n_113), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x6_ASAP7_75t_SL g449 ( .A(n_114), .B(n_116), .Y(n_449) );
OR2x6_ASAP7_75t_SL g784 ( .A(n_114), .B(n_115), .Y(n_784) );
OR2x2_ASAP7_75t_L g794 ( .A(n_114), .B(n_116), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_785), .B(n_788), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_446), .B1(n_450), .B2(n_784), .Y(n_123) );
INVx2_ASAP7_75t_L g790 ( .A(n_124), .Y(n_790) );
INVx1_ASAP7_75t_L g800 ( .A(n_124), .Y(n_800) );
INVx2_ASAP7_75t_L g806 ( .A(n_124), .Y(n_806) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_367), .Y(n_124) );
NOR3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_279), .C(n_319), .Y(n_125) );
OAI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_194), .B1(n_243), .B2(n_258), .C(n_261), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_158), .Y(n_128) );
INVx2_ASAP7_75t_L g276 ( .A(n_129), .Y(n_276) );
AND2x2_ASAP7_75t_L g306 ( .A(n_129), .B(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g244 ( .A(n_130), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g251 ( .A(n_130), .B(n_184), .Y(n_251) );
INVx2_ASAP7_75t_L g257 ( .A(n_130), .Y(n_257) );
AND2x2_ASAP7_75t_L g266 ( .A(n_130), .B(n_160), .Y(n_266) );
INVx1_ASAP7_75t_L g282 ( .A(n_130), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_130), .B(n_328), .Y(n_327) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_131), .A2(n_512), .B(n_516), .Y(n_511) );
INVx2_ASAP7_75t_SL g521 ( .A(n_131), .Y(n_521) );
BUFx4f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
AND2x4_ASAP7_75t_L g156 ( .A(n_133), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_133), .B(n_157), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_144), .B(n_156), .Y(n_134) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_142), .Y(n_136) );
INVx1_ASAP7_75t_L g485 ( .A(n_137), .Y(n_485) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
AND2x6_ASAP7_75t_L g154 ( .A(n_138), .B(n_147), .Y(n_154) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g152 ( .A(n_140), .B(n_149), .Y(n_152) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_142), .Y(n_547) );
AND2x2_ASAP7_75t_L g148 ( .A(n_143), .B(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_143), .Y(n_474) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
BUFx3_ASAP7_75t_L g475 ( .A(n_146), .Y(n_475) );
INVx2_ASAP7_75t_L g465 ( .A(n_147), .Y(n_465) );
AND2x4_ASAP7_75t_L g461 ( .A(n_148), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g469 ( .A(n_149), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B(n_155), .Y(n_150) );
INVxp67_ASAP7_75t_L g490 ( .A(n_152), .Y(n_490) );
INVxp67_ASAP7_75t_L g488 ( .A(n_154), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_155), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_155), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_155), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_155), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_155), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_155), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_155), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_155), .A2(n_467), .B(n_468), .C(n_470), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_155), .B(n_156), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_155), .A2(n_468), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_155), .A2(n_468), .B(n_514), .C(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g524 ( .A(n_155), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_155), .A2(n_468), .B(n_537), .C(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_155), .A2(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_SL g175 ( .A(n_156), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_156), .B(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_156), .A2(n_460), .B(n_471), .Y(n_459) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_172), .Y(n_158) );
INVx4_ASAP7_75t_L g247 ( .A(n_159), .Y(n_247) );
AND2x2_ASAP7_75t_L g278 ( .A(n_159), .B(n_185), .Y(n_278) );
AND2x2_ASAP7_75t_L g354 ( .A(n_159), .B(n_328), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_159), .B(n_184), .Y(n_396) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_160), .B(n_184), .Y(n_283) );
AND2x2_ASAP7_75t_L g307 ( .A(n_160), .B(n_185), .Y(n_307) );
BUFx2_ASAP7_75t_L g323 ( .A(n_160), .Y(n_323) );
NOR2x1_ASAP7_75t_SL g426 ( .A(n_160), .B(n_328), .Y(n_426) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_164), .Y(n_160) );
INVx3_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_162), .A2(n_204), .B1(n_543), .B2(n_548), .Y(n_542) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_163), .B(n_551), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_170), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_170), .Y(n_192) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_170), .A2(n_231), .B(n_235), .Y(n_230) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_170), .A2(n_231), .B(n_235), .Y(n_293) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g303 ( .A(n_172), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_172), .A2(n_370), .B1(n_372), .B2(n_374), .C(n_379), .Y(n_369) );
AND2x2_ASAP7_75t_L g389 ( .A(n_172), .B(n_282), .Y(n_389) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_184), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
INVx1_ASAP7_75t_L g298 ( .A(n_174), .Y(n_298) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_182), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_175), .B(n_183), .Y(n_182) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_175), .A2(n_176), .B(n_182), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_181), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_184), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g267 ( .A(n_184), .B(n_255), .Y(n_267) );
INVx2_ASAP7_75t_L g309 ( .A(n_184), .Y(n_309) );
AND2x2_ASAP7_75t_L g442 ( .A(n_184), .B(n_257), .Y(n_442) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_185), .Y(n_299) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_192), .A2(n_493), .B(n_499), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_226), .C(n_241), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
INVx2_ASAP7_75t_L g356 ( .A(n_196), .Y(n_356) );
AND2x2_ASAP7_75t_L g401 ( .A(n_196), .B(n_278), .Y(n_401) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g346 ( .A(n_197), .Y(n_346) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_197), .B(n_273), .Y(n_361) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_204), .B(n_205), .Y(n_197) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_198), .A2(n_204), .B(n_205), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_203), .Y(n_198) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_204), .A2(n_219), .B(n_225), .Y(n_218) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_204), .A2(n_219), .B(n_225), .Y(n_238) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_204), .A2(n_533), .B(n_539), .Y(n_532) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_204), .A2(n_533), .B(n_539), .Y(n_562) );
INVx2_ASAP7_75t_L g315 ( .A(n_206), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_206), .B(n_345), .Y(n_371) );
AND2x4_ASAP7_75t_L g404 ( .A(n_206), .B(n_351), .Y(n_404) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
AND2x2_ASAP7_75t_L g242 ( .A(n_207), .B(n_237), .Y(n_242) );
OR2x2_ASAP7_75t_L g272 ( .A(n_207), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_SL g341 ( .A(n_207), .B(n_293), .Y(n_341) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx2_ASAP7_75t_L g286 ( .A(n_208), .Y(n_286) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
OAI21x1_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_212), .B(n_216), .Y(n_209) );
INVx1_ASAP7_75t_L g217 ( .A(n_211), .Y(n_217) );
INVx2_ASAP7_75t_L g273 ( .A(n_218), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_220), .B(n_224), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_226), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_236), .Y(n_227) );
AND2x2_ASAP7_75t_L g241 ( .A(n_228), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g314 ( .A(n_228), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g399 ( .A(n_228), .Y(n_399) );
BUFx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g259 ( .A(n_229), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g378 ( .A(n_229), .B(n_238), .Y(n_378) );
AND2x2_ASAP7_75t_L g382 ( .A(n_229), .B(n_248), .Y(n_382) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g351 ( .A(n_230), .Y(n_351) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_230), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_236), .B(n_259), .Y(n_335) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_237), .B(n_260), .Y(n_445) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g249 ( .A(n_238), .B(n_240), .Y(n_249) );
AND2x2_ASAP7_75t_L g331 ( .A(n_238), .B(n_293), .Y(n_331) );
AND2x2_ASAP7_75t_L g350 ( .A(n_238), .B(n_239), .Y(n_350) );
BUFx2_ASAP7_75t_L g271 ( .A(n_239), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_239), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
BUFx3_ASAP7_75t_L g248 ( .A(n_240), .Y(n_248) );
INVxp67_ASAP7_75t_L g291 ( .A(n_240), .Y(n_291) );
INVx1_ASAP7_75t_L g264 ( .A(n_242), .Y(n_264) );
AND2x2_ASAP7_75t_L g300 ( .A(n_242), .B(n_271), .Y(n_300) );
NAND2xp33_ASAP7_75t_L g381 ( .A(n_242), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g418 ( .A(n_242), .B(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_246), .B1(n_249), .B2(n_250), .C(n_252), .Y(n_243) );
AND2x2_ASAP7_75t_L g347 ( .A(n_244), .B(n_247), .Y(n_347) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_244), .B(n_307), .Y(n_366) );
AND2x2_ASAP7_75t_L g384 ( .A(n_244), .B(n_309), .Y(n_384) );
AND2x2_ASAP7_75t_L g439 ( .A(n_244), .B(n_278), .Y(n_439) );
INVx1_ASAP7_75t_L g255 ( .A(n_245), .Y(n_255) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_245), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_246), .Y(n_391) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_247), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_247), .B(n_298), .Y(n_373) );
AND2x2_ASAP7_75t_L g340 ( .A(n_248), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g376 ( .A(n_248), .Y(n_376) );
AND2x2_ASAP7_75t_L g285 ( .A(n_249), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_249), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g427 ( .A(n_249), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_249), .B(n_351), .Y(n_437) );
AND2x4_ASAP7_75t_L g353 ( .A(n_250), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g424 ( .A(n_251), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
OR2x2_ASAP7_75t_L g295 ( .A(n_256), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g302 ( .A(n_257), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g333 ( .A(n_257), .B(n_307), .Y(n_333) );
AND2x2_ASAP7_75t_L g407 ( .A(n_257), .B(n_328), .Y(n_407) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g355 ( .A(n_259), .B(n_356), .Y(n_355) );
OAI32xp33_ASAP7_75t_L g420 ( .A1(n_259), .A2(n_421), .A3(n_423), .B1(n_424), .B2(n_427), .Y(n_420) );
AND2x4_ASAP7_75t_L g292 ( .A(n_260), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g390 ( .A(n_260), .B(n_293), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B1(n_268), .B2(n_274), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_SL g379 ( .A1(n_263), .A2(n_277), .B(n_380), .C(n_381), .Y(n_379) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g363 ( .A(n_264), .B(n_291), .Y(n_363) );
INVx1_ASAP7_75t_SL g434 ( .A(n_265), .Y(n_434) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x4_ASAP7_75t_L g337 ( .A(n_267), .B(n_276), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_267), .A2(n_416), .B1(n_417), .B2(n_418), .C(n_420), .Y(n_415) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_272), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_275), .A2(n_305), .B1(n_358), .B2(n_359), .Y(n_357) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_276), .A2(n_394), .B(n_402), .C(n_415), .Y(n_393) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g313 ( .A(n_278), .B(n_282), .Y(n_313) );
OAI211xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_284), .B(n_287), .C(n_316), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g310 ( .A(n_282), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g430 ( .A(n_282), .B(n_426), .Y(n_430) );
OAI32xp33_ASAP7_75t_L g387 ( .A1(n_283), .A2(n_388), .A3(n_390), .B1(n_391), .B2(n_392), .Y(n_387) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_286), .B(n_378), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_294), .B1(n_300), .B2(n_301), .C(n_304), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g444 ( .A(n_291), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_292), .B(n_356), .Y(n_358) );
A2O1A1O1Ixp25_ASAP7_75t_L g429 ( .A1(n_292), .A2(n_361), .B(n_377), .C(n_423), .D(n_430), .Y(n_429) );
AOI31xp33_ASAP7_75t_L g431 ( .A1(n_292), .A2(n_313), .A3(n_423), .B(n_430), .Y(n_431) );
AND2x2_ASAP7_75t_L g345 ( .A(n_293), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_295), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx2_ASAP7_75t_L g422 ( .A(n_297), .Y(n_422) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g417 ( .A(n_298), .B(n_309), .Y(n_417) );
INVx1_ASAP7_75t_L g332 ( .A(n_300), .Y(n_332) );
AND2x2_ASAP7_75t_L g317 ( .A(n_301), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AOI31xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_308), .A3(n_312), .B(n_314), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_307), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g440 ( .A(n_307), .B(n_386), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g385 ( .A(n_309), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g411 ( .A(n_309), .Y(n_411) );
INVxp67_ASAP7_75t_L g380 ( .A(n_310), .Y(n_380) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g318 ( .A(n_314), .Y(n_318) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND3xp33_ASAP7_75t_SL g319 ( .A(n_320), .B(n_336), .C(n_352), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_329), .B1(n_333), .B2(n_334), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g406 ( .A(n_323), .Y(n_406) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_327), .Y(n_386) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_327), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_327), .B(n_396), .Y(n_413) );
NAND2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVx1_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_347), .B2(n_348), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_339), .B(n_342), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_345), .A2(n_350), .B1(n_384), .B2(n_385), .C(n_387), .Y(n_383) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2x1_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g423 ( .A(n_350), .Y(n_423) );
AND2x2_ASAP7_75t_L g360 ( .A(n_351), .B(n_361), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_SL g408 ( .A1(n_351), .A2(n_409), .B(n_413), .C(n_414), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_357), .C(n_362), .Y(n_352) );
AND2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
AOI21xp33_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_364), .B(n_365), .Y(n_362) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_393), .C(n_428), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_383), .Y(n_368) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g392 ( .A(n_377), .Y(n_392) );
INVxp67_ASAP7_75t_L g416 ( .A(n_381), .Y(n_416) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g400 ( .A(n_390), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_400), .B2(n_401), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B(n_408), .Y(n_402) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g441 ( .A(n_426), .B(n_442), .Y(n_441) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_432), .B2(n_435), .C(n_438), .Y(n_428) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI31xp33_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .A3(n_441), .B(n_443), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx4_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_448), .A2(n_451), .B1(n_784), .B2(n_790), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_671), .C(n_748), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_623), .Y(n_452) );
NOR2xp67_ASAP7_75t_L g453 ( .A(n_454), .B(n_563), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_500), .B1(n_507), .B2(n_556), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_476), .Y(n_455) );
NOR2xp67_ASAP7_75t_SL g606 ( .A(n_456), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g621 ( .A(n_456), .B(n_622), .Y(n_621) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_456), .B(n_639), .Y(n_638) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_456), .B(n_679), .Y(n_678) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_457), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_457), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g613 ( .A(n_457), .Y(n_613) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_457), .Y(n_618) );
AND2x2_ASAP7_75t_L g647 ( .A(n_457), .B(n_587), .Y(n_647) );
OR2x2_ASAP7_75t_L g651 ( .A(n_457), .B(n_492), .Y(n_651) );
AND2x4_ASAP7_75t_L g664 ( .A(n_457), .B(n_622), .Y(n_664) );
NOR2x1_ASAP7_75t_SL g666 ( .A(n_457), .B(n_479), .Y(n_666) );
AND2x2_ASAP7_75t_L g694 ( .A(n_457), .B(n_572), .Y(n_694) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVxp67_ASAP7_75t_L g553 ( .A(n_461), .Y(n_553) );
NOR2x1p5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g528 ( .A(n_464), .Y(n_528) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x6_ASAP7_75t_L g468 ( .A(n_465), .B(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_468), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_482) );
INVxp67_ASAP7_75t_L g544 ( .A(n_468), .Y(n_544) );
INVx2_ASAP7_75t_L g582 ( .A(n_468), .Y(n_582) );
AND2x2_ASAP7_75t_L g473 ( .A(n_469), .B(n_474), .Y(n_473) );
INVxp33_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
INVx1_ASAP7_75t_L g555 ( .A(n_472), .Y(n_555) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g575 ( .A(n_473), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_475), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_476), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_477), .A2(n_752), .B1(n_754), .B2(n_757), .Y(n_751) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_492), .Y(n_477) );
INVx1_ASAP7_75t_L g506 ( .A(n_478), .Y(n_506) );
AND2x2_ASAP7_75t_L g609 ( .A(n_478), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g614 ( .A(n_478), .B(n_572), .Y(n_614) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g571 ( .A(n_479), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g587 ( .A(n_479), .Y(n_587) );
AND2x2_ASAP7_75t_L g620 ( .A(n_479), .B(n_492), .Y(n_620) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_486), .B(n_491), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_485), .B(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_486) );
INVx2_ASAP7_75t_L g504 ( .A(n_492), .Y(n_504) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_492), .Y(n_589) );
INVx1_ASAP7_75t_L g608 ( .A(n_492), .Y(n_608) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_492), .Y(n_677) );
INVx1_ASAP7_75t_L g689 ( .A(n_492), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI31xp33_ASAP7_75t_SL g743 ( .A1(n_501), .A2(n_744), .A3(n_745), .B(n_746), .Y(n_743) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g668 ( .A(n_503), .B(n_570), .Y(n_668) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g584 ( .A(n_504), .Y(n_584) );
AND2x4_ASAP7_75t_SL g704 ( .A(n_506), .B(n_608), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_507), .A2(n_625), .B(n_628), .Y(n_624) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
INVx2_ASAP7_75t_L g597 ( .A(n_508), .Y(n_597) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_509), .B(n_632), .Y(n_724) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g634 ( .A(n_510), .B(n_540), .Y(n_634) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVxp67_ASAP7_75t_L g559 ( .A(n_511), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_511), .B(n_520), .Y(n_594) );
AND2x4_ASAP7_75t_L g604 ( .A(n_511), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g649 ( .A(n_511), .B(n_541), .Y(n_649) );
INVx2_ASAP7_75t_L g657 ( .A(n_511), .Y(n_657) );
INVx1_ASAP7_75t_L g756 ( .A(n_511), .Y(n_756) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_511), .Y(n_765) );
INVx1_ASAP7_75t_L g702 ( .A(n_517), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_518), .B(n_531), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g558 ( .A(n_519), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g697 ( .A(n_519), .B(n_632), .Y(n_697) );
AND2x2_ASAP7_75t_L g714 ( .A(n_519), .B(n_532), .Y(n_714) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_520), .B(n_562), .Y(n_737) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_530), .Y(n_520) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_521), .A2(n_522), .B(n_530), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_529), .Y(n_522) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g660 ( .A(n_531), .B(n_558), .Y(n_660) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_540), .Y(n_531) );
INVx2_ASAP7_75t_L g566 ( .A(n_532), .Y(n_566) );
NOR2xp67_ASAP7_75t_L g747 ( .A(n_532), .B(n_540), .Y(n_747) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_532), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g663 ( .A(n_540), .B(n_567), .Y(n_663) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_541), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
AND2x4_ASAP7_75t_L g656 ( .A(n_541), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g686 ( .A(n_541), .Y(n_686) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_557), .A2(n_570), .B1(n_708), .B2(n_709), .C(n_710), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x2_ASAP7_75t_L g684 ( .A(n_558), .B(n_685), .Y(n_684) );
BUFx2_ASAP7_75t_L g727 ( .A(n_558), .Y(n_727) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g670 ( .A(n_561), .B(n_594), .Y(n_670) );
INVx3_ASAP7_75t_L g632 ( .A(n_562), .Y(n_632) );
AND2x2_ASAP7_75t_L g764 ( .A(n_562), .B(n_765), .Y(n_764) );
NAND3xp33_ASAP7_75t_SL g563 ( .A(n_564), .B(n_595), .C(n_611), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B1(n_585), .B2(n_590), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_565), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g695 ( .A(n_565), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g706 ( .A(n_565), .B(n_601), .Y(n_706) );
AND2x2_ASAP7_75t_L g776 ( .A(n_565), .B(n_649), .Y(n_776) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g605 ( .A(n_567), .Y(n_605) );
INVx1_ASAP7_75t_L g654 ( .A(n_567), .Y(n_654) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI222xp33_ASAP7_75t_L g721 ( .A1(n_569), .A2(n_722), .B1(n_723), .B2(n_725), .C1(n_726), .C2(n_728), .Y(n_721) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_583), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_570), .B(n_597), .Y(n_596) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_570), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g688 ( .A(n_571), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g744 ( .A(n_571), .B(n_618), .Y(n_744) );
INVx2_ASAP7_75t_L g610 ( .A(n_572), .Y(n_610) );
INVx1_ASAP7_75t_L g622 ( .A(n_572), .Y(n_622) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_572), .Y(n_679) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .C(n_577), .Y(n_574) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_584), .Y(n_627) );
INVx3_ASAP7_75t_L g646 ( .A(n_584), .Y(n_646) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g712 ( .A(n_586), .Y(n_712) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g699 ( .A(n_588), .Y(n_699) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g700 ( .A(n_591), .Y(n_700) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g601 ( .A(n_592), .Y(n_601) );
AND2x2_ASAP7_75t_L g719 ( .A(n_592), .B(n_604), .Y(n_719) );
AND2x2_ASAP7_75t_L g782 ( .A(n_592), .B(n_714), .Y(n_782) );
AND2x2_ASAP7_75t_L g711 ( .A(n_593), .B(n_631), .Y(n_711) );
INVx1_ASAP7_75t_L g722 ( .A(n_593), .Y(n_722) );
AND2x2_ASAP7_75t_L g739 ( .A(n_593), .B(n_686), .Y(n_739) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B1(n_602), .B2(n_606), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_598), .A2(n_612), .B(n_615), .Y(n_611) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g643 ( .A(n_601), .B(n_604), .Y(n_643) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g746 ( .A(n_604), .B(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g709 ( .A(n_607), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_608), .Y(n_637) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_609), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g682 ( .A(n_609), .Y(n_682) );
AND2x2_ASAP7_75t_L g780 ( .A(n_609), .B(n_677), .Y(n_780) );
INVx1_ASAP7_75t_L g735 ( .A(n_610), .Y(n_735) );
INVx1_ASAP7_75t_L g641 ( .A(n_612), .Y(n_641) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g730 ( .A(n_613), .Y(n_730) );
INVx4_ASAP7_75t_L g639 ( .A(n_614), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI32xp33_ASAP7_75t_L g710 ( .A1(n_617), .A2(n_711), .A3(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
AND2x2_ASAP7_75t_L g705 ( .A(n_618), .B(n_620), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_SL g768 ( .A1(n_618), .A2(n_769), .B(n_770), .C(n_772), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_620), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g772 ( .A(n_620), .Y(n_772) );
AND2x2_ASAP7_75t_L g626 ( .A(n_621), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g753 ( .A(n_621), .Y(n_753) );
AND2x2_ASAP7_75t_L g759 ( .A(n_621), .B(n_646), .Y(n_759) );
NOR3x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_640), .C(n_658), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_631), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g691 ( .A(n_631), .B(n_656), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_631), .B(n_677), .Y(n_718) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_639), .B(n_646), .Y(n_745) );
INVx2_ASAP7_75t_L g767 ( .A(n_639), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_644), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g731 ( .A1(n_641), .A2(n_732), .B1(n_736), .B2(n_738), .C(n_743), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_642), .A2(n_762), .B1(n_763), .B2(n_766), .Y(n_761) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B1(n_650), .B2(n_652), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g690 ( .A(n_646), .B(n_666), .Y(n_690) );
INVx1_ASAP7_75t_L g696 ( .A(n_646), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_646), .B(n_664), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_649), .B(n_717), .Y(n_783) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_650), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_651), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2x1_ASAP7_75t_SL g769 ( .A(n_654), .B(n_656), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_654), .B(n_754), .Y(n_775) );
OR2x2_ASAP7_75t_L g736 ( .A(n_655), .B(n_737), .Y(n_736) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g771 ( .A(n_656), .B(n_697), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_659), .B(n_665), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B(n_664), .Y(n_659) );
OR2x2_ASAP7_75t_L g723 ( .A(n_662), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g757 ( .A(n_663), .B(n_755), .Y(n_757) );
AND2x2_ASAP7_75t_SL g703 ( .A(n_664), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g713 ( .A(n_664), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B(n_669), .Y(n_665) );
AND2x2_ASAP7_75t_L g698 ( .A(n_666), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_715), .Y(n_672) );
NOR3xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_692), .C(n_707), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_680), .B(n_683), .C(n_687), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g741 ( .A(n_686), .Y(n_741) );
AND2x2_ASAP7_75t_L g754 ( .A(n_686), .B(n_755), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g762 ( .A(n_688), .Y(n_762) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_700), .B(n_701), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_697), .B2(n_698), .Y(n_693) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_694), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_705), .B2(n_706), .Y(n_701) );
INVx1_ASAP7_75t_SL g708 ( .A(n_706), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_712), .B(n_753), .Y(n_752) );
OAI22xp33_ASAP7_75t_SL g778 ( .A1(n_713), .A2(n_779), .B1(n_781), .B2(n_783), .Y(n_778) );
AOI211x1_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_720), .B(n_721), .C(n_731), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g773 ( .A1(n_733), .A2(n_774), .B(n_776), .Y(n_773) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g742 ( .A(n_737), .Y(n_742) );
NOR2xp67_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_740), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_760), .C(n_773), .D(n_777), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_758), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_768), .Y(n_760) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g813 ( .A(n_793), .B(n_814), .Y(n_813) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .Y(n_795) );
INVx1_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
OAI22xp5_ASAP7_75t_SL g799 ( .A1(n_800), .A2(n_801), .B1(n_802), .B2(n_805), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g819 ( .A(n_813), .Y(n_819) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
endmodule