module real_jpeg_7065_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_1),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_1),
.B(n_95),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_2),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_3),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_3),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_3),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_4),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_4),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_4),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_4),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_5),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_5),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_5),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_5),
.B(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_7),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_7),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_7),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_8),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_8),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_8),
.B(n_92),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_8),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_8),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_8),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_8),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_9),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_9),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_9),
.B(n_414),
.Y(n_413)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_11),
.Y(n_241)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_13),
.B(n_133),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_13),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_13),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_13),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_13),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_13),
.B(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_14),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_14),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_14),
.B(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_14),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_14),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_14),
.B(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_15),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_15),
.Y(n_412)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_197),
.B1(n_454),
.B2(n_455),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_18),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_196),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_160),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_21),
.B(n_160),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_101),
.C(n_136),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_22),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.C(n_83),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_23),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.C(n_58),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_24),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_27),
.A2(n_28),
.B1(n_109),
.B2(n_110),
.Y(n_310)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_28),
.B(n_31),
.C(n_37),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_28),
.B(n_110),
.C(n_217),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g349 ( 
.A(n_30),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_31),
.A2(n_35),
.B1(n_111),
.B2(n_115),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_31),
.B(n_111),
.C(n_147),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_31),
.A2(n_35),
.B1(n_364),
.B2(n_365),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_61),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_32),
.B(n_91),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_35),
.B(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_36),
.A2(n_37),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_40),
.Y(n_278)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_41),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_42),
.B(n_58),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.C(n_54),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_43),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_47),
.Y(n_273)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_48),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_49),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_49),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_49),
.B(n_54),
.Y(n_287)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_53),
.Y(n_172)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_53),
.Y(n_381)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_57),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_70),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_81),
.C(n_82),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_71),
.B(n_83),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_80),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_78),
.C(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_76),
.A2(n_79),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_79),
.B(n_155),
.C(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_96),
.C(n_98),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_85),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.C(n_94),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_86),
.A2(n_94),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_86),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_86),
.A2(n_234),
.B1(n_271),
.B2(n_272),
.Y(n_372)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_90),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_93),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_96),
.B(n_98),
.Y(n_299)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_101),
.B(n_136),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_117),
.C(n_125),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_103),
.B(n_110),
.C(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_109),
.A2(n_110),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_111),
.B(n_312),
.C(n_316),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_111),
.A2(n_115),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_118),
.A2(n_141),
.B1(n_259),
.B2(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_118),
.B(n_170),
.C(n_259),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_120),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_135),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_131),
.C(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_151),
.B2(n_159),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_152),
.C(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.C(n_145),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_139),
.A2(n_140),
.B1(n_144),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_144),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_145),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_160),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.CI(n_178),
.CON(n_160),
.SN(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_174),
.B2(n_175),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_170),
.A2(n_173),
.B1(n_258),
.B2(n_265),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_171),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_172),
.Y(n_354)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_192),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_197),
.Y(n_455)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_336),
.B(n_339),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_325),
.B(n_335),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_302),
.B(n_324),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_200),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_289),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_201),
.B(n_289),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_256),
.C(n_283),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_202),
.B(n_323),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g458 ( 
.A(n_202),
.Y(n_458)
);

FAx1_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_229),
.CI(n_235),
.CON(n_202),
.SN(n_202)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_203),
.B(n_229),
.C(n_235),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_216),
.C(n_222),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_204),
.B(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_213),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_206),
.B(n_209),
.C(n_213),
.Y(n_288)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_216),
.A2(n_222),
.B1(n_223),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_216),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_217),
.B(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_318)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_246),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_237),
.B(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_247),
.C(n_254),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_245),
.B(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_251),
.Y(n_388)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_252),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_255),
.B(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_255),
.B(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_255),
.B(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_283),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.C(n_268),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_257),
.A2(n_266),
.B1(n_267),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_268),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.C(n_279),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_269),
.A2(n_270),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_274),
.A2(n_275),
.B1(n_279),
.B2(n_280),
.Y(n_442)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_286),
.C(n_288),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_292),
.C(n_301),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_294),
.B1(n_300),
.B2(n_301),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_322),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_303),
.B(n_322),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_319),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_304),
.A2(n_305),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_308),
.B(n_319),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.C(n_318),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_309),
.B(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_311),
.B(n_318),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_313),
.B1(n_316),
.B2(n_317),
.Y(n_361)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_326),
.B(n_336),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_328),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_337),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_328),
.B(n_337),
.Y(n_453)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_332),
.CI(n_334),
.CON(n_328),
.SN(n_328)
);

OAI31xp33_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_450),
.A3(n_451),
.B(n_453),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_444),
.B(n_449),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_429),
.B(n_443),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_383),
.B(n_428),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_373),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_344),
.B(n_373),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_362),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_359),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_346),
.B(n_359),
.C(n_362),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.C(n_355),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_375)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_355),
.B(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_368),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_363),
.B(n_438),
.C(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.C(n_382),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_376),
.A2(n_382),
.B1(n_420),
.B2(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_380),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_382),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_422),
.B(n_427),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_408),
.B(n_421),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_393),
.B(n_407),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_404),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_404),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_399),
.B(n_403),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_399),
.Y(n_403)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_403),
.A2(n_410),
.B1(n_415),
.B2(n_416),
.Y(n_409)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_403),
.Y(n_415)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_417),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_417),
.Y(n_421)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_410),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_411),
.A2(n_413),
.B(n_415),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B(n_420),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_424),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_431),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_435),
.B2(n_436),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_437),
.C(n_440),
.Y(n_445)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.Y(n_449)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_447),
.Y(n_448)
);


endmodule