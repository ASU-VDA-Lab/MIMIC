module fake_jpeg_20003_n_300 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_17),
.B1(n_33),
.B2(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_16),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_45),
.B(n_24),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_31),
.B1(n_34),
.B2(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_20),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_18),
.B1(n_34),
.B2(n_23),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_30),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_64),
.B(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_81),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_79),
.B1(n_89),
.B2(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_83),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_82),
.B(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_60),
.B1(n_55),
.B2(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_38),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_32),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_94),
.B1(n_98),
.B2(n_97),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_32),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_97),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_96),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_33),
.B1(n_24),
.B2(n_32),
.Y(n_95)
);

OAI211xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_19),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_70),
.B(n_71),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_51),
.B(n_24),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_114),
.B(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_62),
.B1(n_51),
.B2(n_54),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_118),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_62),
.B(n_50),
.C(n_0),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_65),
.A2(n_62),
.B1(n_50),
.B2(n_2),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_5),
.C(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_7),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_91),
.B(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_100),
.B1(n_99),
.B2(n_64),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_111),
.Y(n_186)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_96),
.B1(n_86),
.B2(n_66),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_144),
.B(n_157),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_73),
.B1(n_78),
.B2(n_80),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_75),
.B1(n_88),
.B2(n_76),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_148),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_126),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_140),
.B1(n_142),
.B2(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_84),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_77),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_77),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_8),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_153),
.B(n_156),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_77),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_109),
.B(n_9),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_10),
.B(n_11),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_10),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_11),
.Y(n_188)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_135),
.A3(n_151),
.B1(n_147),
.B2(n_106),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_183),
.B(n_188),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_177),
.B1(n_159),
.B2(n_158),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_109),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_119),
.C(n_122),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_176),
.C(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_119),
.C(n_128),
.Y(n_176)
);

OAI22x1_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_111),
.B1(n_116),
.B2(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_110),
.B(n_116),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_143),
.B(n_115),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_113),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_141),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_125),
.B1(n_160),
.B2(n_108),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_177),
.Y(n_192)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_157),
.B(n_161),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_203),
.B1(n_211),
.B2(n_170),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_148),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_196),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_136),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_197),
.B(n_171),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_188),
.C(n_168),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_125),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_207),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_205),
.B1(n_210),
.B2(n_166),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_208),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_104),
.B1(n_130),
.B2(n_108),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_130),
.B1(n_104),
.B2(n_150),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_141),
.B1(n_13),
.B2(n_14),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_185),
.B(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_176),
.C(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_223),
.C(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_232),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_165),
.C(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_236),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_163),
.C(n_172),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_215),
.B(n_168),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_166),
.B1(n_164),
.B2(n_182),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_192),
.B1(n_220),
.B2(n_233),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_183),
.B1(n_190),
.B2(n_164),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_174),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_204),
.B1(n_210),
.B2(n_196),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_213),
.B1(n_205),
.B2(n_218),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_207),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_245),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_189),
.B(n_167),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_215),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

XOR2x2_ASAP7_75t_SL g248 ( 
.A(n_230),
.B(n_199),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_253),
.C(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_251),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_228),
.B(n_175),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_224),
.B(n_190),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_197),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_260),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_261),
.B1(n_239),
.B2(n_255),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_224),
.B1(n_219),
.B2(n_203),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_241),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_268),
.B(n_245),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_238),
.B(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_250),
.C(n_242),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_261),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_266),
.B1(n_259),
.B2(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_284),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_258),
.B(n_248),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_272),
.B(n_276),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_12),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_274),
.B(n_270),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_287),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_167),
.B(n_14),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_280),
.C(n_13),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_290),
.B(n_16),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_293),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_295),
.B(n_294),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_291),
.B(n_16),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_299),
.Y(n_300)
);


endmodule