module fake_jpeg_29521_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_36),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_17),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_20),
.B1(n_22),
.B2(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_23),
.B1(n_17),
.B2(n_19),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_23),
.B(n_19),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_30),
.A2(n_25),
.B1(n_1),
.B2(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_8),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_68),
.B(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_70),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_14),
.B1(n_8),
.B2(n_10),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_57),
.C(n_50),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_62),
.B(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_57),
.B1(n_45),
.B2(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_66),
.B1(n_70),
.B2(n_69),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_44),
.B(n_62),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.C(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_98),
.B(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_66),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_76),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_82),
.C(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_80),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_89),
.B(n_94),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_103),
.B(n_84),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_88),
.B(n_82),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_75),
.B1(n_78),
.B2(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_107),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_79),
.B1(n_45),
.B2(n_84),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_109),
.Y(n_113)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_111),
.B(n_100),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_108),
.B(n_109),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_113),
.C(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_112),
.Y(n_118)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_116),
.B(n_71),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_65),
.Y(n_121)
);


endmodule