module real_jpeg_3977_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_1),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_196),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_1),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_1),
.A2(n_26),
.B1(n_172),
.B2(n_272),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_92),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_92),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_2),
.A2(n_81),
.B1(n_92),
.B2(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_4),
.Y(n_415)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_6),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_6),
.B(n_10),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_7),
.A2(n_85),
.B1(n_122),
.B2(n_127),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_45),
.B1(n_85),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_7),
.A2(n_85),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_23),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_10),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_52),
.B1(n_162),
.B2(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_52),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_52),
.B1(n_183),
.B2(n_228),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_10),
.A2(n_136),
.B(n_264),
.C(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_10),
.B(n_57),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_10),
.B(n_298),
.C(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_120),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_10),
.B(n_115),
.C(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_10),
.B(n_28),
.Y(n_335)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_12),
.Y(n_412)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_410),
.B(n_413),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_145),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_18),
.B(n_140),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.C(n_138),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_19),
.B(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_54),
.C(n_87),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_20),
.A2(n_193),
.B1(n_204),
.B2(n_205),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_20),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_20),
.B(n_152),
.C(n_205),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_20),
.B(n_243),
.C(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_20),
.A2(n_204),
.B1(n_243),
.B2(n_336),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_20),
.A2(n_204),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_50),
.B2(n_53),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_21),
.A2(n_27),
.B1(n_50),
.B2(n_53),
.Y(n_230)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_24),
.Y(n_134)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_25),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_27),
.B(n_50),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_27),
.A2(n_53),
.B1(n_130),
.B2(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_27),
.A2(n_50),
.B(n_53),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_40),
.Y(n_27)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_30),
.Y(n_196)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_31),
.Y(n_264)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_33),
.Y(n_266)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_36),
.Y(n_128)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_52),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_53),
.A2(n_130),
.B(n_137),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_54),
.A2(n_87),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_54),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_54),
.B(n_230),
.C(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_54),
.A2(n_385),
.B1(n_387),
.B2(n_394),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_83),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_56),
.A2(n_69),
.B1(n_156),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_56),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_56),
.A2(n_69),
.B1(n_156),
.B2(n_161),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_56),
.A2(n_69),
.B(n_161),
.Y(n_347)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_59),
.Y(n_173)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_59),
.Y(n_177)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_66),
.Y(n_185)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_69),
.B(n_161),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_69),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_76),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_83),
.A2(n_209),
.B1(n_211),
.B2(n_242),
.Y(n_241)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_87),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B1(n_120),
.B2(n_121),
.Y(n_87)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_88),
.Y(n_388)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_94),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_95),
.A2(n_120),
.B1(n_194),
.B2(n_199),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_95),
.B(n_194),
.Y(n_389)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_97),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_96),
.A2(n_97),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_112),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_97),
.A2(n_388),
.B(n_389),
.Y(n_387)
);

AOI22x1_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_105),
.B2(n_108),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_114),
.Y(n_318)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_129),
.B(n_138),
.Y(n_407)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_139),
.B(n_194),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_405),
.B(n_409),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_376),
.B(n_402),
.Y(n_146)
);

OAI211xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_275),
.B(n_371),
.C(n_375),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_250),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_149),
.A2(n_250),
.B(n_372),
.C(n_374),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_231),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_150),
.B(n_231),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_206),
.C(n_218),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_151),
.B(n_206),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_192),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_167),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_153),
.A2(n_167),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_153),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_153),
.A2(n_260),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_154),
.A2(n_155),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_167),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_174),
.B1(n_181),
.B2(n_188),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_168),
.A2(n_223),
.B(n_226),
.Y(n_222)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_171),
.Y(n_301)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_174),
.B(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_175),
.A2(n_227),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_175),
.A2(n_227),
.B1(n_271),
.B2(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_193),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_193),
.A2(n_205),
.B1(n_220),
.B2(n_221),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_193),
.B(n_220),
.C(n_315),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_193),
.A2(n_205),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_193),
.B(n_256),
.C(n_347),
.Y(n_365)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx6_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_213),
.B2(n_217),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_213),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_217),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_213),
.A2(n_237),
.B(n_238),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_214),
.B(n_227),
.Y(n_321)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_229),
.C(n_230),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_220),
.A2(n_221),
.B1(n_294),
.B2(n_302),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_220),
.B(n_302),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_222),
.Y(n_363)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_230),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_230),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_230),
.A2(n_256),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_230),
.A2(n_256),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_230),
.A2(n_256),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_230),
.B(n_381),
.C(n_386),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_248),
.B2(n_249),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_239),
.B1(n_240),
.B2(n_247),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_239),
.B(n_247),
.C(n_249),
.Y(n_401)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_243),
.B(n_246),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_243),
.A2(n_332),
.B1(n_333),
.B2(n_336),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_243),
.Y(n_336)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_246),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_246),
.A2(n_391),
.B1(n_395),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_251),
.B(n_253),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.C(n_261),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_254),
.B(n_258),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_270),
.C(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_260),
.B(n_328),
.C(n_330),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_261),
.B(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_262),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_263),
.A2(n_269),
.B1(n_270),
.B2(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_270),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_289),
.Y(n_290)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_355),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_340),
.B(n_354),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_325),
.B(n_339),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_312),
.B(n_324),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_304),
.B(n_311),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_291),
.B(n_303),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_288),
.B(n_290),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_292),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_292),
.B(n_334),
.C(n_336),
.Y(n_350)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_322),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_338),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_338),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.B1(n_331),
.B2(n_337),
.Y(n_326)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_342),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_350),
.C(n_351),
.Y(n_367)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_358),
.B(n_366),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_358),
.C(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_362),
.C(n_364),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_362),
.A2(n_364),
.B1(n_365),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_362),
.Y(n_370)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_368),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_397),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_390),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_390),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_386),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_387),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.C(n_396),
.Y(n_390)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_396),
.B(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_401),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_401),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_408),
.Y(n_409)
);

BUFx4f_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g414 ( 
.A(n_411),
.Y(n_414)
);

INVx13_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);


endmodule