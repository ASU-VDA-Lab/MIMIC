module fake_jpeg_27937_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_21),
.B(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_17),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_13),
.C(n_8),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.C(n_20),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_13),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_18),
.Y(n_39)
);

XNOR2x1_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_15),
.Y(n_36)
);

OAI22x1_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_40),
.B(n_42),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_11),
.C(n_16),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.C(n_26),
.Y(n_50)
);

OAI221xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_25),
.B1(n_22),
.B2(n_2),
.C(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_49),
.B1(n_22),
.B2(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_46),
.C(n_26),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_6),
.B1(n_7),
.B2(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_0),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_0),
.Y(n_56)
);


endmodule