module fake_jpeg_979_n_681 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_681);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_681;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_65),
.B(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_73),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_76),
.B(n_79),
.Y(n_180)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_77),
.Y(n_218)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_8),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

BUFx12f_ASAP7_75t_SL g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2x1_ASAP7_75t_SL g195 ( 
.A(n_86),
.B(n_95),
.Y(n_195)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_90),
.Y(n_206)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_40),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_123),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_45),
.B(n_8),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_102),
.B(n_110),
.Y(n_223)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_103),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_60),
.B(n_8),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_48),
.C(n_25),
.Y(n_167)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_105),
.Y(n_208)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_11),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_44),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_112),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_46),
.B(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_117),
.B(n_124),
.Y(n_216)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_7),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_20),
.B(n_12),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_26),
.Y(n_134)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_24),
.Y(n_127)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_22),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_48),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_24),
.Y(n_133)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_134),
.B(n_142),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_28),
.B1(n_26),
.B2(n_57),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_137),
.A2(n_139),
.B1(n_153),
.B2(n_203),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_61),
.B1(n_24),
.B2(n_52),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_42),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_84),
.B(n_42),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_146),
.B(n_151),
.Y(n_279)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_155),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_95),
.A2(n_61),
.B1(n_24),
.B2(n_52),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_36),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_159),
.B(n_164),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_57),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_166),
.B(n_177),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_167),
.B(n_211),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_87),
.A2(n_21),
.B1(n_30),
.B2(n_59),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_174),
.A2(n_185),
.B1(n_210),
.B2(n_34),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_92),
.A2(n_21),
.B1(n_30),
.B2(n_61),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_176),
.A2(n_183),
.B1(n_189),
.B2(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_181),
.B(n_182),
.Y(n_267)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_118),
.A2(n_30),
.B1(n_61),
.B2(n_55),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_66),
.A2(n_61),
.B1(n_52),
.B2(n_55),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_25),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_188),
.Y(n_269)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_72),
.A2(n_53),
.B1(n_58),
.B2(n_56),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_132),
.B(n_53),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_194),
.B(n_212),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_86),
.A2(n_34),
.B1(n_58),
.B2(n_56),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_80),
.A2(n_129),
.B1(n_128),
.B2(n_120),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_82),
.A2(n_101),
.B1(n_88),
.B2(n_119),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_126),
.B(n_62),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_64),
.B(n_62),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_98),
.A2(n_51),
.B1(n_49),
.B2(n_47),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_219),
.A2(n_123),
.B1(n_107),
.B2(n_2),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_225),
.B(n_262),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_227),
.Y(n_339)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_228),
.Y(n_310)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_230),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_231),
.B(n_261),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_36),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_244),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_99),
.B1(n_100),
.B2(n_115),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_233),
.A2(n_264),
.B1(n_163),
.B2(n_184),
.Y(n_306)
);

AO22x1_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_122),
.B1(n_113),
.B2(n_114),
.Y(n_234)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_236),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_238),
.Y(n_348)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_241),
.Y(n_344)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_32),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_245),
.A2(n_246),
.B1(n_272),
.B2(n_275),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_81),
.B1(n_108),
.B2(n_94),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_247),
.Y(n_346)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_161),
.A2(n_34),
.B1(n_22),
.B2(n_47),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_249),
.A2(n_273),
.B1(n_298),
.B2(n_154),
.Y(n_309)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_250),
.Y(n_354)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_154),
.Y(n_256)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_140),
.B(n_32),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_259),
.B(n_263),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_203),
.A2(n_96),
.B1(n_83),
.B2(n_35),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_260),
.A2(n_299),
.B1(n_5),
.B2(n_6),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_192),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_178),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_35),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_220),
.A2(n_165),
.B1(n_170),
.B2(n_169),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

BUFx2_ASAP7_75t_SL g271 ( 
.A(n_202),
.Y(n_271)
);

INVx13_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_153),
.A2(n_116),
.B1(n_51),
.B2(n_49),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_161),
.A2(n_179),
.B1(n_206),
.B2(n_138),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_162),
.B(n_0),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_283),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_205),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_278),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_204),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_280),
.Y(n_364)
);

AO22x1_ASAP7_75t_SL g281 ( 
.A1(n_139),
.A2(n_121),
.B1(n_2),
.B2(n_3),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_288),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_205),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_286),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_159),
.B(n_1),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_147),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_190),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_206),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_289),
.B(n_290),
.Y(n_356)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_145),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_1),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_291),
.B(n_296),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_152),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_292),
.B(n_301),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_138),
.A2(n_121),
.B1(n_13),
.B2(n_14),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_215),
.B(n_175),
.Y(n_316)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_172),
.B(n_2),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_152),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_297),
.A2(n_5),
.B1(n_6),
.B2(n_19),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_179),
.A2(n_14),
.B1(n_18),
.B2(n_16),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_149),
.A2(n_14),
.B1(n_18),
.B2(n_15),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_141),
.B(n_4),
.Y(n_300)
);

NAND2x1_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_200),
.Y(n_337)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_157),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_148),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_303),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_306),
.B(n_337),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_251),
.A2(n_163),
.B1(n_184),
.B2(n_168),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_307),
.A2(n_315),
.B1(n_319),
.B2(n_331),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

OAI22x1_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_213),
.B1(n_208),
.B2(n_222),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_245),
.A2(n_168),
.B1(n_222),
.B2(n_171),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_316),
.A2(n_336),
.B(n_361),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_294),
.A2(n_215),
.B1(n_175),
.B2(n_171),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_246),
.A2(n_213),
.B1(n_208),
.B2(n_199),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_242),
.A2(n_149),
.B1(n_156),
.B2(n_160),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_283),
.A2(n_199),
.B(n_160),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_200),
.C(n_156),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_262),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_239),
.A2(n_200),
.B1(n_12),
.B2(n_14),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_305),
.B1(n_358),
.B2(n_297),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_347),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_15),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_351),
.B(n_259),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_360),
.B1(n_264),
.B2(n_229),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_272),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_227),
.A2(n_5),
.B1(n_6),
.B2(n_284),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_296),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_372),
.Y(n_417)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_359),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_371),
.A2(n_407),
.B1(n_409),
.B2(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_327),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_312),
.A2(n_285),
.B1(n_244),
.B2(n_232),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_374),
.A2(n_388),
.B1(n_396),
.B2(n_397),
.Y(n_429)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_375),
.Y(n_431)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_314),
.Y(n_376)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_378),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_291),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_387),
.Y(n_425)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_382),
.B(n_411),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_312),
.A2(n_285),
.B(n_234),
.C(n_281),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_385),
.B(n_408),
.Y(n_416)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_311),
.B(n_336),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_386),
.A2(n_340),
.B1(n_354),
.B2(n_344),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_276),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_352),
.A2(n_285),
.B1(n_234),
.B2(n_263),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_304),
.B(n_279),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_389),
.B(n_391),
.Y(n_422)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_348),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_300),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_394),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_300),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_395),
.B(n_398),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_352),
.A2(n_269),
.B1(n_293),
.B2(n_281),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_358),
.A2(n_243),
.B1(n_288),
.B2(n_301),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_322),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_323),
.A2(n_230),
.B1(n_237),
.B2(n_241),
.Y(n_399)
);

AO21x2_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_414),
.B(n_334),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_315),
.A2(n_225),
.B1(n_238),
.B2(n_240),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_400),
.A2(n_365),
.B1(n_335),
.B2(n_345),
.Y(n_424)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_401),
.B(n_403),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_322),
.B(n_270),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_323),
.A2(n_258),
.B1(n_253),
.B2(n_250),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_405),
.A2(n_342),
.B1(n_325),
.B2(n_313),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_226),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_316),
.A2(n_248),
.B(n_289),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_332),
.B(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_364),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_347),
.A2(n_255),
.B1(n_290),
.B2(n_266),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_385),
.A2(n_360),
.B1(n_353),
.B2(n_361),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_421),
.A2(n_436),
.B1(n_442),
.B2(n_371),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_339),
.B(n_337),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_423),
.A2(n_426),
.B(n_427),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_424),
.A2(n_387),
.B1(n_389),
.B2(n_403),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_413),
.A2(n_337),
.B(n_338),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_317),
.B(n_356),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_372),
.B(n_319),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_432),
.C(n_448),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_366),
.B(n_345),
.C(n_267),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_434),
.A2(n_414),
.B1(n_393),
.B2(n_397),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_404),
.A2(n_307),
.B1(n_340),
.B2(n_354),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_396),
.A2(n_344),
.B1(n_328),
.B2(n_346),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_440),
.B(n_451),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_383),
.A2(n_364),
.B(n_328),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_404),
.A2(n_333),
.B1(n_320),
.B2(n_313),
.Y(n_442)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_447),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_257),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_405),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_400),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_386),
.A2(n_346),
.B(n_334),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_388),
.A2(n_333),
.B1(n_325),
.B2(n_342),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_452),
.A2(n_377),
.B1(n_378),
.B2(n_381),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_411),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_369),
.C(n_367),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_430),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g525 ( 
.A(n_457),
.B(n_473),
.C(n_446),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_374),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_458),
.B(n_442),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_459),
.A2(n_484),
.B(n_491),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_460),
.A2(n_463),
.B1(n_464),
.B2(n_466),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_429),
.A2(n_377),
.B1(n_393),
.B2(n_373),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_429),
.A2(n_373),
.B1(n_402),
.B2(n_392),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_423),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_465),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_416),
.A2(n_443),
.B1(n_452),
.B2(n_439),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_470),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_416),
.A2(n_373),
.B1(n_394),
.B2(n_379),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_471),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_430),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_474),
.A2(n_482),
.B1(n_485),
.B2(n_449),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_475),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_447),
.A2(n_428),
.B1(n_450),
.B2(n_425),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_483),
.Y(n_513)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_415),
.Y(n_477)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_417),
.B(n_382),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_480),
.C(n_490),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_376),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_453),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_421),
.A2(n_375),
.B1(n_399),
.B2(n_390),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_422),
.B(n_412),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_R g484 ( 
.A(n_426),
.B(n_409),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_418),
.A2(n_447),
.B1(n_436),
.B2(n_422),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_447),
.A2(n_384),
.B1(n_401),
.B2(n_395),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_492),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_425),
.B(n_407),
.Y(n_487)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_487),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_444),
.Y(n_488)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_489),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_391),
.C(n_280),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_427),
.A2(n_359),
.B(n_362),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_451),
.A2(n_370),
.B(n_362),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_449),
.B(n_410),
.Y(n_493)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_472),
.Y(n_497)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_SL g498 ( 
.A(n_461),
.B(n_455),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_498),
.B(n_515),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_458),
.B(n_445),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_499),
.B(n_503),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_500),
.B(n_507),
.Y(n_550)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_456),
.B(n_448),
.C(n_455),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_510),
.C(n_511),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_456),
.B(n_432),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_491),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_512),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_490),
.C(n_465),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_480),
.B(n_420),
.C(n_446),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_483),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_431),
.Y(n_516)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_516),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_473),
.B(n_431),
.Y(n_517)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_517),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_486),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_518),
.B(n_433),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_460),
.A2(n_485),
.B1(n_488),
.B2(n_461),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_519),
.A2(n_476),
.B1(n_469),
.B2(n_463),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_479),
.B(n_453),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_523),
.C(n_511),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_493),
.Y(n_522)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_522),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_484),
.B(n_437),
.Y(n_523)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_438),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_528),
.B(n_343),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_521),
.A2(n_467),
.B(n_492),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_533),
.B(n_539),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_535),
.A2(n_538),
.B1(n_544),
.B2(n_554),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_524),
.A2(n_513),
.B1(n_496),
.B2(n_527),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_536),
.A2(n_546),
.B1(n_548),
.B2(n_497),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_482),
.B1(n_459),
.B2(n_472),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_516),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_466),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_540),
.B(n_541),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_502),
.B(n_470),
.Y(n_541)
);

MAJx2_ASAP7_75t_L g590 ( 
.A(n_542),
.B(n_256),
.C(n_329),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_519),
.A2(n_501),
.B1(n_527),
.B2(n_513),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_524),
.A2(n_471),
.B1(n_472),
.B2(n_475),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_521),
.A2(n_467),
.B(n_492),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_547),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_514),
.A2(n_447),
.B1(n_464),
.B2(n_477),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_489),
.C(n_478),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_549),
.B(n_552),
.C(n_529),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_523),
.A2(n_506),
.B(n_504),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_557),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_503),
.B(n_435),
.C(n_438),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_495),
.B(n_437),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_499),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_494),
.A2(n_447),
.B1(n_419),
.B2(n_435),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_504),
.A2(n_441),
.B(n_433),
.Y(n_557)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_558),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_494),
.A2(n_441),
.B1(n_410),
.B2(n_333),
.Y(n_560)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_560),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_514),
.A2(n_441),
.B1(n_343),
.B2(n_329),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_562),
.A2(n_509),
.B1(n_529),
.B2(n_505),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_563),
.B(n_509),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_550),
.B(n_526),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_562),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_566),
.A2(n_581),
.B1(n_557),
.B2(n_556),
.Y(n_602)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_568),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_495),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_569),
.B(n_578),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_559),
.B(n_520),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_570),
.B(n_571),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_549),
.B(n_512),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_572),
.B(n_573),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_506),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_545),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_574),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_526),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_576),
.A2(n_584),
.B1(n_563),
.B2(n_548),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_531),
.B(n_517),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_545),
.A2(n_535),
.B1(n_544),
.B2(n_543),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_542),
.B(n_528),
.Y(n_583)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_583),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_540),
.B(n_530),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_532),
.B(n_498),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_585),
.B(n_252),
.C(n_278),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_536),
.A2(n_530),
.B1(n_497),
.B2(n_498),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_586),
.A2(n_321),
.B1(n_310),
.B2(n_357),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_587),
.B(n_589),
.C(n_590),
.Y(n_592)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_588),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_541),
.B(n_505),
.C(n_268),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_577),
.A2(n_533),
.B(n_547),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_593),
.A2(n_597),
.B(n_605),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_568),
.A2(n_543),
.B1(n_561),
.B2(n_555),
.Y(n_594)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_594),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_587),
.B(n_532),
.C(n_534),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_595),
.B(n_598),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_582),
.A2(n_551),
.B(n_555),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_534),
.C(n_546),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_586),
.A2(n_561),
.B1(n_556),
.B2(n_537),
.Y(n_599)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_599),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_600),
.B(n_602),
.Y(n_623)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_601),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_582),
.A2(n_321),
.B(n_310),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_607),
.A2(n_609),
.B1(n_575),
.B2(n_235),
.Y(n_627)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_566),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_608),
.B(n_610),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_574),
.A2(n_357),
.B1(n_274),
.B2(n_287),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_567),
.A2(n_295),
.B1(n_265),
.B2(n_254),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_572),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_578),
.C(n_573),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_614),
.B(n_618),
.Y(n_636)
);

FAx1_ASAP7_75t_L g617 ( 
.A(n_601),
.B(n_564),
.CI(n_581),
.CON(n_617),
.SN(n_617)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_617),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_606),
.B(n_565),
.C(n_589),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_596),
.B(n_579),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_619),
.B(n_622),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_565),
.C(n_585),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_624),
.B(n_631),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_611),
.B(n_580),
.C(n_590),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_625),
.B(n_629),
.Y(n_637)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_627),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_596),
.A2(n_228),
.B(n_236),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_628),
.A2(n_605),
.B(n_604),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_592),
.B(n_355),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_613),
.B(n_355),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_630),
.B(n_604),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_593),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_626),
.A2(n_601),
.B1(n_591),
.B2(n_602),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_633),
.B(n_635),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_620),
.A2(n_591),
.B1(n_594),
.B2(n_599),
.Y(n_634)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_634),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_614),
.B(n_595),
.C(n_598),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_603),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_641),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_623),
.B(n_631),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_632),
.B(n_603),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_643),
.B(n_617),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_617),
.Y(n_644)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_644),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_645),
.B(n_629),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_647),
.B(n_648),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_618),
.B(n_608),
.C(n_597),
.Y(n_648)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_649),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_640),
.A2(n_615),
.B(n_621),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_653),
.A2(n_657),
.B(n_659),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_639),
.B(n_616),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_655),
.B(n_660),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_625),
.Y(n_657)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_658),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_644),
.A2(n_622),
.B(n_612),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_636),
.B(n_624),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_656),
.B(n_646),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_662),
.B(n_666),
.Y(n_670)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_650),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_654),
.B(n_634),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_667),
.B(n_668),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_651),
.B(n_646),
.C(n_648),
.Y(n_668)
);

AO21x1_ASAP7_75t_L g669 ( 
.A1(n_663),
.A2(n_652),
.B(n_653),
.Y(n_669)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_669),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_664),
.B(n_635),
.C(n_657),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_671),
.B(n_672),
.Y(n_674)
);

XOR2xp5_ASAP7_75t_L g672 ( 
.A(n_665),
.B(n_659),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_673),
.B(n_668),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_661),
.C(n_673),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_677),
.A2(n_678),
.B(n_642),
.Y(n_679)
);

A2O1A1O1Ixp25_ASAP7_75t_L g678 ( 
.A1(n_674),
.A2(n_675),
.B(n_670),
.C(n_637),
.D(n_633),
.Y(n_678)
);

OAI31xp33_ASAP7_75t_SL g680 ( 
.A1(n_679),
.A2(n_627),
.A3(n_607),
.B(n_609),
.Y(n_680)
);

BUFx24_ASAP7_75t_SL g681 ( 
.A(n_680),
.Y(n_681)
);


endmodule