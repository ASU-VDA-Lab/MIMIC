module real_jpeg_30128_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_42),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_91)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_4),
.A2(n_18),
.B(n_20),
.C(n_21),
.D(n_29),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_25),
.Y(n_80)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_25),
.B(n_37),
.C(n_80),
.D(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_4),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_57),
.B(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_31),
.B1(n_42),
.B2(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_25),
.B(n_38),
.C(n_41),
.Y(n_37)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_7),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_76),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_75),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_63),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_63),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_47),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_33),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_19),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI32xp33_ASAP7_75t_L g60 ( 
.A1(n_19),
.A2(n_20),
.A3(n_25),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_24),
.B(n_28),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_24),
.A2(n_40),
.A3(n_44),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_41),
.B2(n_45),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_42),
.Y(n_81)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_44),
.B(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_60),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_56),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_53),
.A2(n_91),
.B(n_100),
.Y(n_99)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_98),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.C(n_71),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_69),
.B1(n_70),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_87),
.B(n_107),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B(n_106),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_101),
.B(n_105),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);


endmodule