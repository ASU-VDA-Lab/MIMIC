module real_aes_7340_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_0), .A2(n_176), .B(n_177), .C(n_181), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_1), .B(n_171), .Y(n_182) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_3), .B(n_136), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_4), .A2(n_117), .B(n_452), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_5), .A2(n_122), .B(n_127), .C(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_6), .A2(n_117), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_7), .B(n_171), .Y(n_458) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_8), .A2(n_150), .B(n_200), .Y(n_199) );
AND2x6_ASAP7_75t_L g122 ( .A(n_9), .B(n_123), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_10), .A2(n_122), .B(n_127), .C(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g513 ( .A(n_11), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_12), .B(n_39), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_13), .B(n_180), .Y(n_490) );
INVx1_ASAP7_75t_L g146 ( .A(n_14), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_15), .B(n_136), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_16), .A2(n_137), .B(n_498), .C(n_500), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_17), .B(n_171), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_18), .B(n_164), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_19), .A2(n_127), .B(n_158), .C(n_163), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_20), .A2(n_179), .B(n_194), .C(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_21), .B(n_180), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_22), .A2(n_75), .B1(n_707), .B2(n_708), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_22), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_23), .B(n_180), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_24), .Y(n_439) );
INVx1_ASAP7_75t_L g464 ( .A(n_25), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_26), .A2(n_127), .B(n_163), .C(n_203), .Y(n_202) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_27), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_28), .Y(n_486) );
INVx1_ASAP7_75t_L g540 ( .A(n_29), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_30), .A2(n_117), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g120 ( .A(n_31), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_32), .A2(n_125), .B(n_130), .C(n_140), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_33), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_34), .A2(n_179), .B(n_455), .C(n_457), .Y(n_454) );
INVxp67_ASAP7_75t_L g541 ( .A(n_35), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_36), .B(n_205), .Y(n_204) );
CKINVDCx14_ASAP7_75t_R g453 ( .A(n_37), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_38), .A2(n_127), .B(n_163), .C(n_463), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_40), .A2(n_181), .B(n_511), .C(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_41), .B(n_156), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_42), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_43), .B(n_136), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_44), .B(n_117), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_45), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_46), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_47), .A2(n_125), .B(n_140), .C(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_48), .A2(n_86), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_48), .Y(n_734) );
INVx1_ASAP7_75t_L g178 ( .A(n_49), .Y(n_178) );
INVx1_ASAP7_75t_L g215 ( .A(n_50), .Y(n_215) );
INVx1_ASAP7_75t_L g476 ( .A(n_51), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_52), .B(n_117), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_53), .Y(n_167) );
CKINVDCx14_ASAP7_75t_R g509 ( .A(n_54), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_55), .Y(n_736) );
INVx1_ASAP7_75t_L g123 ( .A(n_56), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_57), .B(n_117), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_58), .B(n_171), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_59), .A2(n_162), .B(n_225), .C(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
INVx1_ASAP7_75t_SL g456 ( .A(n_61), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_62), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_63), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_64), .B(n_171), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_65), .B(n_137), .Y(n_191) );
INVx1_ASAP7_75t_L g442 ( .A(n_66), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_67), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_68), .B(n_133), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_69), .A2(n_127), .B(n_140), .C(n_251), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_70), .Y(n_223) );
INVx1_ASAP7_75t_L g724 ( .A(n_71), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_72), .A2(n_117), .B(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_73), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_74), .A2(n_117), .B(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_75), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_76), .A2(n_156), .B(n_536), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_77), .Y(n_461) );
INVx1_ASAP7_75t_L g496 ( .A(n_78), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_79), .B(n_132), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_80), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_81), .A2(n_117), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g499 ( .A(n_82), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_83), .Y(n_719) );
INVx2_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
INVx1_ASAP7_75t_L g489 ( .A(n_85), .Y(n_489) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_86), .A2(n_101), .B1(n_720), .B2(n_729), .C1(n_737), .C2(n_743), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_86), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_87), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_88), .B(n_180), .Y(n_192) );
OR2x2_ASAP7_75t_L g104 ( .A(n_89), .B(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g429 ( .A(n_89), .Y(n_429) );
OR2x2_ASAP7_75t_L g728 ( .A(n_89), .B(n_718), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_90), .A2(n_127), .B(n_140), .C(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_91), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
INVxp67_ASAP7_75t_L g228 ( .A(n_93), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_94), .B(n_150), .Y(n_514) );
INVx1_ASAP7_75t_L g187 ( .A(n_95), .Y(n_187) );
INVx1_ASAP7_75t_L g252 ( .A(n_96), .Y(n_252) );
INVx2_ASAP7_75t_L g479 ( .A(n_97), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_98), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g217 ( .A(n_99), .B(n_142), .Y(n_217) );
OAI222xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_706), .B1(n_709), .B2(n_715), .C1(n_716), .C2(n_719), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_108), .B1(n_427), .B2(n_430), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g712 ( .A(n_104), .Y(n_712) );
OR2x2_ASAP7_75t_L g428 ( .A(n_105), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g718 ( .A(n_105), .Y(n_718) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_109), .A2(n_710), .B1(n_713), .B2(n_714), .Y(n_709) );
XOR2xp5_ASAP7_75t_L g731 ( .A(n_109), .B(n_732), .Y(n_731) );
OR3x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_341), .C(n_384), .Y(n_109) );
NAND5xp2_ASAP7_75t_L g110 ( .A(n_111), .B(n_268), .C(n_298), .D(n_315), .E(n_330), .Y(n_110) );
AOI221xp5_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_183), .B1(n_230), .B2(n_236), .C(n_240), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_152), .Y(n_112) );
OR2x2_ASAP7_75t_L g245 ( .A(n_113), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g285 ( .A(n_113), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g303 ( .A(n_113), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_113), .B(n_238), .Y(n_320) );
OR2x2_ASAP7_75t_L g332 ( .A(n_113), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_113), .B(n_291), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_113), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_113), .B(n_269), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_113), .B(n_277), .Y(n_383) );
AND2x2_ASAP7_75t_L g415 ( .A(n_113), .B(n_169), .Y(n_415) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_113), .Y(n_423) );
INVx5_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_114), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g242 ( .A(n_114), .B(n_218), .Y(n_242) );
BUFx2_ASAP7_75t_L g265 ( .A(n_114), .Y(n_265) );
AND2x2_ASAP7_75t_L g294 ( .A(n_114), .B(n_153), .Y(n_294) );
AND2x2_ASAP7_75t_L g349 ( .A(n_114), .B(n_246), .Y(n_349) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_147), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_124), .B(n_142), .Y(n_115) );
BUFx2_ASAP7_75t_L g156 ( .A(n_117), .Y(n_156) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_118), .B(n_122), .Y(n_188) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
INVx1_ASAP7_75t_L g195 ( .A(n_120), .Y(n_195) );
INVx1_ASAP7_75t_L g129 ( .A(n_121), .Y(n_129) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
INVx3_ASAP7_75t_L g137 ( .A(n_121), .Y(n_137) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_121), .Y(n_180) );
INVx1_ASAP7_75t_L g205 ( .A(n_121), .Y(n_205) );
INVx4_ASAP7_75t_SL g141 ( .A(n_122), .Y(n_141) );
BUFx3_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_126), .A2(n_141), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_126), .A2(n_141), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_126), .A2(n_141), .B(n_453), .C(n_454), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_126), .A2(n_141), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_126), .A2(n_141), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_126), .A2(n_141), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_126), .A2(n_141), .B(n_537), .C(n_538), .Y(n_536) );
INVx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
BUFx3_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_128), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_135), .C(n_138), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_132), .A2(n_138), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g441 ( .A1(n_132), .A2(n_442), .B(n_443), .C(n_444), .Y(n_441) );
O2A1O1Ixp5_ASAP7_75t_L g488 ( .A1(n_132), .A2(n_444), .B(n_489), .C(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx4_ASAP7_75t_L g226 ( .A(n_134), .Y(n_226) );
INVx2_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_136), .B(n_228), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_136), .A2(n_161), .B(n_464), .C(n_465), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_136), .A2(n_226), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_137), .B(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g500 ( .A(n_139), .Y(n_500) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g165 ( .A(n_142), .Y(n_165) );
INVx1_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_142), .A2(n_212), .B(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_142), .A2(n_188), .B(n_461), .C(n_462), .Y(n_460) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_142), .A2(n_507), .B(n_514), .Y(n_506) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_L g151 ( .A(n_143), .B(n_144), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx3_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_149), .A2(n_186), .B(n_196), .Y(n_185) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_149), .A2(n_249), .B(n_257), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_149), .B(n_258), .Y(n_257) );
AO21x2_ASAP7_75t_L g437 ( .A1(n_149), .A2(n_438), .B(n_445), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_149), .B(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_149), .B(n_492), .Y(n_491) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_150), .A2(n_201), .B(n_202), .Y(n_200) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_152), .B(n_303), .Y(n_312) );
OAI32xp33_ASAP7_75t_L g326 ( .A1(n_152), .A2(n_262), .A3(n_327), .B1(n_328), .B2(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_152), .B(n_328), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_152), .B(n_245), .Y(n_369) );
INVx1_ASAP7_75t_SL g398 ( .A(n_152), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_152), .B(n_185), .C(n_349), .D(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_169), .Y(n_152) );
INVx5_ASAP7_75t_L g239 ( .A(n_153), .Y(n_239) );
AND2x2_ASAP7_75t_L g269 ( .A(n_153), .B(n_170), .Y(n_269) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_153), .Y(n_348) );
AND2x2_ASAP7_75t_L g418 ( .A(n_153), .B(n_365), .Y(n_418) );
OR2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_166), .Y(n_153) );
AOI21xp5_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_157), .B(n_164), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_161), .Y(n_158) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_162), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_165), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_168), .A2(n_485), .B(n_491), .Y(n_484) );
AND2x4_ASAP7_75t_L g291 ( .A(n_169), .B(n_239), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_169), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g325 ( .A(n_169), .B(n_246), .Y(n_325) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g238 ( .A(n_170), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g277 ( .A(n_170), .B(n_248), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_170), .B(n_247), .Y(n_286) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_182), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_179), .B(n_456), .Y(n_455) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g511 ( .A(n_180), .Y(n_511) );
INVx2_ASAP7_75t_L g444 ( .A(n_181), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g354 ( .A1(n_183), .A2(n_355), .B1(n_357), .B2(n_359), .C1(n_362), .C2(n_363), .Y(n_354) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_207), .Y(n_183) );
AND2x2_ASAP7_75t_L g287 ( .A(n_184), .B(n_288), .Y(n_287) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_184), .B(n_265), .C(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_199), .Y(n_184) );
INVx5_ASAP7_75t_SL g235 ( .A(n_185), .Y(n_235) );
OAI322xp33_ASAP7_75t_L g240 ( .A1(n_185), .A2(n_241), .A3(n_243), .B1(n_244), .B2(n_259), .C1(n_262), .C2(n_264), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_185), .B(n_233), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_185), .B(n_219), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_188), .A2(n_439), .B(n_440), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_188), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_193), .A2(n_204), .B(n_206), .Y(n_203) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx2_ASAP7_75t_L g534 ( .A(n_198), .Y(n_534) );
INVx2_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_199), .B(n_209), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_207), .B(n_272), .Y(n_327) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g306 ( .A(n_208), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_218), .Y(n_208) );
OR2x2_ASAP7_75t_L g234 ( .A(n_209), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_209), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g274 ( .A(n_209), .B(n_219), .Y(n_274) );
AND2x2_ASAP7_75t_L g297 ( .A(n_209), .B(n_233), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_209), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g313 ( .A(n_209), .B(n_272), .Y(n_313) );
AND2x2_ASAP7_75t_L g321 ( .A(n_209), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_209), .B(n_281), .Y(n_371) );
INVx5_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g261 ( .A(n_210), .B(n_235), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_210), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g288 ( .A(n_210), .B(n_219), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_210), .B(n_335), .Y(n_376) );
OR2x2_ASAP7_75t_L g392 ( .A(n_210), .B(n_336), .Y(n_392) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_210), .B(n_353), .Y(n_399) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_210), .Y(n_406) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_217), .Y(n_210) );
AND2x2_ASAP7_75t_L g260 ( .A(n_218), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g310 ( .A(n_218), .B(n_233), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_218), .B(n_235), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_218), .B(n_272), .Y(n_394) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_219), .B(n_235), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_219), .B(n_233), .Y(n_282) );
OR2x2_ASAP7_75t_L g336 ( .A(n_219), .B(n_233), .Y(n_336) );
AND2x2_ASAP7_75t_L g353 ( .A(n_219), .B(n_232), .Y(n_353) );
INVxp67_ASAP7_75t_L g375 ( .A(n_219), .Y(n_375) );
AND2x2_ASAP7_75t_L g402 ( .A(n_219), .B(n_272), .Y(n_402) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_219), .Y(n_409) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_220), .A2(n_451), .B(n_458), .Y(n_450) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_220), .A2(n_474), .B(n_480), .Y(n_473) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_220), .A2(n_494), .B(n_501), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_225), .A2(n_252), .B(n_253), .C(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_226), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_226), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_232), .B(n_283), .Y(n_356) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g272 ( .A(n_233), .B(n_235), .Y(n_272) );
OR2x2_ASAP7_75t_L g339 ( .A(n_233), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
OR2x2_ASAP7_75t_L g344 ( .A(n_234), .B(n_336), .Y(n_344) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g243 ( .A(n_238), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_238), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g244 ( .A(n_239), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_239), .B(n_246), .Y(n_279) );
INVx2_ASAP7_75t_L g324 ( .A(n_239), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_239), .B(n_277), .Y(n_337) );
AND2x2_ASAP7_75t_L g362 ( .A(n_239), .B(n_286), .Y(n_362) );
INVx1_ASAP7_75t_L g314 ( .A(n_244), .Y(n_314) );
INVx2_ASAP7_75t_SL g301 ( .A(n_245), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_246), .Y(n_304) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_247), .Y(n_267) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g365 ( .A(n_248), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_256), .Y(n_249) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g457 ( .A(n_255), .Y(n_457) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g334 ( .A(n_261), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g340 ( .A(n_261), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_261), .A2(n_343), .B1(n_345), .B2(n_350), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_261), .B(n_353), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_262), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g296 ( .A(n_263), .Y(n_296) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g278 ( .A(n_265), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_265), .B(n_269), .Y(n_329) );
AND2x2_ASAP7_75t_L g352 ( .A(n_265), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g328 ( .A(n_267), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_275), .C(n_289), .Y(n_268) );
INVx1_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_269), .A2(n_401), .B1(n_403), .B2(n_404), .C(n_407), .Y(n_400) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g419 ( .A(n_272), .Y(n_419) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g368 ( .A(n_274), .B(n_307), .Y(n_368) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_278), .B(n_280), .C(n_284), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OAI32xp33_ASAP7_75t_L g393 ( .A1(n_282), .A2(n_283), .A3(n_346), .B1(n_383), .B2(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
AND2x2_ASAP7_75t_L g425 ( .A(n_285), .B(n_324), .Y(n_425) );
AND2x2_ASAP7_75t_L g372 ( .A(n_286), .B(n_324), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_286), .B(n_294), .Y(n_390) );
AOI31xp33_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .A3(n_293), .B(n_295), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_291), .B(n_303), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_291), .B(n_301), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_291), .A2(n_321), .B1(n_411), .B2(n_414), .C(n_416), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g316 ( .A(n_296), .B(n_317), .Y(n_316) );
AOI222xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_305), .B1(n_308), .B2(n_311), .C1(n_313), .C2(n_314), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g381 ( .A(n_300), .Y(n_381) );
INVx1_ASAP7_75t_L g403 ( .A(n_303), .Y(n_403) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_306), .A2(n_417), .B1(n_419), .B2(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B1(n_321), .B2(n_323), .C(n_326), .Y(n_315) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g412 ( .A(n_318), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g387 ( .A(n_323), .Y(n_387) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g351 ( .A(n_324), .Y(n_351) );
INVx1_ASAP7_75t_L g333 ( .A(n_325), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_328), .B(n_415), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_337), .B2(n_338), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g424 ( .A(n_337), .Y(n_424) );
INVxp33_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_339), .B(n_383), .Y(n_382) );
OAI32xp33_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_374), .A3(n_375), .B1(n_376), .B2(n_377), .Y(n_373) );
NAND4xp25_ASAP7_75t_L g341 ( .A(n_342), .B(n_354), .C(n_366), .D(n_378), .Y(n_341) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_349), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
CKINVDCx16_ASAP7_75t_R g359 ( .A(n_360), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_363), .A2(n_379), .B1(n_396), .B2(n_399), .C(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g414 ( .A(n_365), .B(n_415), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_370), .B2(n_372), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_375), .B(n_406), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND4xp25_ASAP7_75t_L g384 ( .A(n_385), .B(n_395), .C(n_410), .D(n_421), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B(n_391), .C(n_393), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g426 ( .A(n_413), .Y(n_426) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_426), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx6_ASAP7_75t_L g713 ( .A(n_428), .Y(n_713) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_429), .B(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g714 ( .A(n_430), .Y(n_714) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_431), .B(n_661), .Y(n_430) );
NOR4xp25_ASAP7_75t_L g431 ( .A(n_432), .B(n_598), .C(n_632), .D(n_648), .Y(n_431) );
NAND4xp25_ASAP7_75t_SL g432 ( .A(n_433), .B(n_527), .C(n_562), .D(n_578), .Y(n_432) );
AOI222xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_468), .B1(n_502), .B2(n_515), .C1(n_520), .C2(n_526), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI31xp33_ASAP7_75t_L g694 ( .A1(n_435), .A2(n_695), .A3(n_696), .B(n_698), .Y(n_694) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_447), .Y(n_435) );
AND2x2_ASAP7_75t_L g669 ( .A(n_436), .B(n_449), .Y(n_669) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g519 ( .A(n_437), .Y(n_519) );
AND2x2_ASAP7_75t_L g526 ( .A(n_437), .B(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_L g583 ( .A(n_437), .B(n_450), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_447), .B(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_448), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_448), .B(n_530), .Y(n_573) );
AND2x2_ASAP7_75t_L g666 ( .A(n_448), .B(n_606), .Y(n_666) );
OAI321xp33_ASAP7_75t_L g700 ( .A1(n_448), .A2(n_519), .A3(n_673), .B1(n_701), .B2(n_703), .C(n_704), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_448), .B(n_505), .C(n_613), .D(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_459), .Y(n_448) );
AND2x2_ASAP7_75t_L g568 ( .A(n_449), .B(n_517), .Y(n_568) );
AND2x2_ASAP7_75t_L g587 ( .A(n_449), .B(n_519), .Y(n_587) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g518 ( .A(n_450), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g543 ( .A(n_450), .B(n_459), .Y(n_543) );
AND2x2_ASAP7_75t_L g629 ( .A(n_450), .B(n_517), .Y(n_629) );
INVx3_ASAP7_75t_SL g517 ( .A(n_459), .Y(n_517) );
AND2x2_ASAP7_75t_L g561 ( .A(n_459), .B(n_548), .Y(n_561) );
OR2x2_ASAP7_75t_L g594 ( .A(n_459), .B(n_519), .Y(n_594) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_459), .Y(n_601) );
AND2x2_ASAP7_75t_L g630 ( .A(n_459), .B(n_518), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_459), .B(n_603), .Y(n_645) );
AND2x2_ASAP7_75t_L g677 ( .A(n_459), .B(n_669), .Y(n_677) );
AND2x2_ASAP7_75t_L g686 ( .A(n_459), .B(n_531), .Y(n_686) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_466), .Y(n_459) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_481), .Y(n_469) );
INVx1_ASAP7_75t_SL g654 ( .A(n_470), .Y(n_654) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g522 ( .A(n_471), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g504 ( .A(n_472), .B(n_483), .Y(n_504) );
AND2x2_ASAP7_75t_L g590 ( .A(n_472), .B(n_506), .Y(n_590) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g560 ( .A(n_473), .B(n_493), .Y(n_560) );
OR2x2_ASAP7_75t_L g571 ( .A(n_473), .B(n_506), .Y(n_571) );
AND2x2_ASAP7_75t_L g597 ( .A(n_473), .B(n_506), .Y(n_597) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_473), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_481), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_481), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g570 ( .A(n_482), .B(n_571), .Y(n_570) );
AOI322xp5_ASAP7_75t_L g656 ( .A1(n_482), .A2(n_560), .A3(n_566), .B1(n_597), .B2(n_647), .C1(n_657), .C2(n_659), .Y(n_656) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_483), .B(n_505), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_483), .B(n_506), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_483), .B(n_523), .Y(n_577) );
AND2x2_ASAP7_75t_L g631 ( .A(n_483), .B(n_597), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_483), .Y(n_635) );
AND2x2_ASAP7_75t_L g647 ( .A(n_483), .B(n_493), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_483), .B(n_522), .Y(n_679) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g544 ( .A(n_484), .B(n_493), .Y(n_544) );
BUFx3_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
AND3x2_ASAP7_75t_L g640 ( .A(n_484), .B(n_620), .C(n_641), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g503 ( .A(n_493), .B(n_504), .C(n_505), .Y(n_503) );
INVx1_ASAP7_75t_SL g523 ( .A(n_493), .Y(n_523) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_493), .Y(n_625) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g619 ( .A(n_504), .B(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g626 ( .A(n_504), .Y(n_626) );
AND2x2_ASAP7_75t_L g664 ( .A(n_505), .B(n_642), .Y(n_664) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx3_ASAP7_75t_L g545 ( .A(n_506), .Y(n_545) );
AND2x2_ASAP7_75t_L g620 ( .A(n_506), .B(n_523), .Y(n_620) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
OR2x2_ASAP7_75t_L g564 ( .A(n_517), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g683 ( .A(n_517), .B(n_583), .Y(n_683) );
AND2x2_ASAP7_75t_L g697 ( .A(n_517), .B(n_519), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_518), .B(n_531), .Y(n_638) );
AND2x2_ASAP7_75t_L g685 ( .A(n_518), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g548 ( .A(n_519), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g565 ( .A(n_519), .B(n_531), .Y(n_565) );
INVx1_ASAP7_75t_L g575 ( .A(n_519), .Y(n_575) );
AND2x2_ASAP7_75t_L g606 ( .A(n_519), .B(n_531), .Y(n_606) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_521), .A2(n_649), .B1(n_653), .B2(n_655), .C(n_656), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_522), .B(n_524), .Y(n_521) );
AND2x2_ASAP7_75t_L g552 ( .A(n_522), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_525), .B(n_559), .Y(n_702) );
AOI322xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_544), .A3(n_545), .B1(n_546), .B2(n_552), .C1(n_554), .C2(n_561), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_543), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g582 ( .A(n_530), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_530), .B(n_593), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_530), .A2(n_543), .B(n_617), .C(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_530), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_530), .B(n_587), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_530), .B(n_669), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_530), .B(n_697), .Y(n_696) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_531), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_531), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g658 ( .A(n_531), .B(n_545), .Y(n_658) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_535), .B(n_542), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_533), .A2(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g550 ( .A(n_535), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_542), .Y(n_551) );
INVx1_ASAP7_75t_L g633 ( .A(n_543), .Y(n_633) );
OAI31xp33_ASAP7_75t_L g643 ( .A1(n_543), .A2(n_568), .A3(n_644), .B(n_646), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_543), .B(n_549), .Y(n_695) );
INVx1_ASAP7_75t_SL g556 ( .A(n_544), .Y(n_556) );
AND2x2_ASAP7_75t_L g589 ( .A(n_544), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g670 ( .A(n_544), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g555 ( .A(n_545), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g580 ( .A(n_545), .Y(n_580) );
AND2x2_ASAP7_75t_L g607 ( .A(n_545), .B(n_560), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_545), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g699 ( .A(n_545), .B(n_647), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_547), .B(n_617), .Y(n_690) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g586 ( .A(n_549), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_SL g604 ( .A(n_549), .Y(n_604) );
NAND2xp33_ASAP7_75t_SL g554 ( .A(n_555), .B(n_557), .Y(n_554) );
OAI211xp5_ASAP7_75t_SL g598 ( .A1(n_556), .A2(n_599), .B(n_605), .C(n_621), .Y(n_598) );
OR2x2_ASAP7_75t_L g673 ( .A(n_556), .B(n_654), .Y(n_673) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
CKINVDCx16_ASAP7_75t_R g610 ( .A(n_558), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_558), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g579 ( .A(n_560), .B(n_580), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B(n_569), .C(n_572), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_SL g613 ( .A(n_565), .Y(n_613) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_568), .B(n_606), .Y(n_611) );
INVx1_ASAP7_75t_L g617 ( .A(n_568), .Y(n_617) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g576 ( .A(n_571), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g609 ( .A(n_571), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g671 ( .A(n_571), .Y(n_671) );
AOI21xp33_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B(n_576), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_574), .A2(n_585), .B(n_588), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B(n_584), .C(n_591), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_579), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_582), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g595 ( .A(n_583), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_585), .A2(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_590), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g615 ( .A(n_590), .Y(n_615) );
AOI21xp33_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_595), .B(n_596), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g646 ( .A(n_597), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_603), .B(n_629), .Y(n_655) );
AND2x2_ASAP7_75t_L g668 ( .A(n_603), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g682 ( .A(n_603), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g692 ( .A(n_603), .B(n_630), .Y(n_692) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_608), .C(n_616), .Y(n_605) );
INVx1_ASAP7_75t_L g652 ( .A(n_606), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B1(n_612), .B2(n_614), .Y(n_608) );
OR2x2_ASAP7_75t_L g614 ( .A(n_610), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_610), .B(n_671), .Y(n_693) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g687 ( .A(n_620), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_627), .B1(n_630), .B2(n_631), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g705 ( .A(n_625), .Y(n_705) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g651 ( .A(n_629), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_634), .B(n_636), .C(n_643), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_651), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR5xp2_ASAP7_75t_L g661 ( .A(n_662), .B(n_680), .C(n_688), .D(n_694), .E(n_700), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_665), .B(n_667), .C(n_674), .Y(n_662) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_672), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_677), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_687), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g703 ( .A(n_683), .Y(n_703) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_693), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
CKINVDCx16_ASAP7_75t_R g715 ( .A(n_706), .Y(n_715) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_726), .Y(n_721) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_SL g742 ( .A(n_723), .Y(n_742) );
INVx1_ASAP7_75t_L g741 ( .A(n_725), .Y(n_741) );
OA21x2_ASAP7_75t_L g744 ( .A1(n_725), .A2(n_742), .B(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_726), .A2(n_731), .B(n_735), .Y(n_730) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_SL g735 ( .A(n_728), .B(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g745 ( .A(n_728), .Y(n_745) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
CKINVDCx6p67_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
endmodule