module fake_jpeg_14730_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_3),
.B(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_2),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_6),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_33),
.B1(n_29),
.B2(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_36),
.B1(n_17),
.B2(n_20),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_11),
.B(n_16),
.C(n_21),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_10),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_7),
.B(n_8),
.C(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_9),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_22),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_67),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_63),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_75),
.B1(n_72),
.B2(n_59),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_73),
.C(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_23),
.C(n_25),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_26),
.B(n_74),
.Y(n_83)
);


endmodule