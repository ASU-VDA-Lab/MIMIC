module fake_ariane_778_n_1768 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1768);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1768;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_70),
.Y(n_164)
);

BUFx8_ASAP7_75t_SL g165 ( 
.A(n_113),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_34),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_20),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_47),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_99),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_14),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_41),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_20),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_133),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_55),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_46),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_89),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_56),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_11),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_24),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_36),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_65),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_13),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_67),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_72),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_11),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_101),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_49),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_43),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_22),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_124),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_53),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_5),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_68),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_48),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_23),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_82),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_0),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_53),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_22),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_36),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_93),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_61),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_75),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_142),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_40),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_134),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_118),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_64),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_116),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_40),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_96),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_63),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_123),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_84),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_37),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_97),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_112),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_94),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_121),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_1),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_31),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_98),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_106),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_81),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_157),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_2),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_27),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_57),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_48),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_87),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_23),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_144),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_74),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_86),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_27),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_145),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_3),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_154),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_55),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_111),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_95),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_17),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_37),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_14),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_73),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_12),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_109),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_2),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_35),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_110),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_10),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_12),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_69),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_136),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_66),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_19),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_51),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_54),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_52),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_28),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_50),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_148),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_21),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_49),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_51),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_126),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_119),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_62),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_39),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_80),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_5),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_177),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_165),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_1),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_163),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_266),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_220),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_164),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_184),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_176),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_184),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_185),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_185),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_250),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_188),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_188),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_194),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_206),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_190),
.B(n_4),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_256),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_274),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_190),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_196),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_306),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_169),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_250),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_196),
.B(n_4),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_203),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_250),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_170),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_250),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_203),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_173),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_174),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_217),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_217),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_228),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_178),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_215),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_228),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_231),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_232),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_300),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_232),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_235),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_235),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_237),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_237),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_239),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_189),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_238),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_239),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_205),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_207),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_208),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_209),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_300),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_291),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_303),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_211),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_216),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_218),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_221),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_236),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_162),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_300),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_241),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_245),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_318),
.B(n_166),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_241),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_386),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_316),
.A2(n_304),
.B1(n_230),
.B2(n_281),
.Y(n_405)
);

NAND2x1p5_ASAP7_75t_L g406 ( 
.A(n_323),
.B(n_200),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_323),
.B(n_295),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_354),
.A2(n_223),
.B(n_166),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_325),
.B(n_243),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_354),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_327),
.B(n_295),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_327),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_318),
.B(n_223),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_329),
.B(n_309),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_331),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_331),
.B(n_243),
.Y(n_432)
);

INVxp33_ASAP7_75t_SL g433 ( 
.A(n_317),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_332),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_332),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_338),
.B(n_167),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_339),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_344),
.B(n_309),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_344),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_348),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_321),
.B(n_240),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_341),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_353),
.B(n_249),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_321),
.B(n_240),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_350),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_360),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_457),
.Y(n_462)
);

AND3x2_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_343),
.C(n_335),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_398),
.B(n_334),
.Y(n_465)
);

INVx6_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_427),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_394),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_405),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_433),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_427),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_420),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_420),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g477 ( 
.A(n_437),
.B(n_249),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_427),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_445),
.B(n_356),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_403),
.B(n_364),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_403),
.B(n_330),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_452),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_405),
.A2(n_263),
.B1(n_253),
.B2(n_257),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_405),
.B(n_357),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_427),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_369),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_445),
.B(n_454),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_392),
.A2(n_428),
.B1(n_437),
.B2(n_406),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_392),
.A2(n_389),
.B1(n_385),
.B2(n_384),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_427),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_403),
.B(n_345),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_454),
.B(n_370),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_441),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_396),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_441),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_412),
.B(n_316),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_441),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_447),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_447),
.B(n_373),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_394),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_374),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_437),
.A2(n_388),
.B1(n_368),
.B2(n_372),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_433),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_441),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_362),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_396),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_415),
.B(n_377),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_441),
.B(n_375),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_402),
.B(n_337),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_437),
.A2(n_388),
.B1(n_372),
.B2(n_368),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_416),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_SL g527 ( 
.A1(n_393),
.A2(n_365),
.B(n_364),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_451),
.B(n_376),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_441),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_441),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_406),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_444),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_397),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_460),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_451),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_397),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_444),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_416),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_435),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_444),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_460),
.B(n_387),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_397),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_397),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_444),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_437),
.A2(n_406),
.B1(n_460),
.B2(n_421),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_460),
.B(n_366),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_444),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_437),
.A2(n_406),
.B1(n_421),
.B2(n_412),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_435),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_406),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_435),
.B(n_380),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_412),
.Y(n_560)
);

AO22x2_ASAP7_75t_L g561 ( 
.A1(n_393),
.A2(n_367),
.B1(n_167),
.B2(n_281),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_412),
.B(n_381),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_393),
.B(n_340),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_421),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_435),
.B(n_382),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_421),
.B(n_301),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_429),
.B(n_161),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_435),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_446),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_423),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_426),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_423),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

BUFx6f_ASAP7_75t_SL g574 ( 
.A(n_426),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_446),
.B(n_260),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_429),
.B(n_301),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_423),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_446),
.B(n_262),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_453),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_423),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_424),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_424),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_453),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_453),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_453),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_453),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_426),
.B(n_268),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_456),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_456),
.B(n_314),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_430),
.B(n_324),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_SL g593 ( 
.A1(n_419),
.A2(n_181),
.B(n_177),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_430),
.B(n_326),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_456),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g596 ( 
.A(n_419),
.B(n_265),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_430),
.B(n_268),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_456),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_429),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_461),
.B(n_333),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_429),
.B(n_181),
.Y(n_601)
);

OAI21xp33_ASAP7_75t_SL g602 ( 
.A1(n_419),
.A2(n_186),
.B(n_183),
.Y(n_602)
);

XOR2x2_ASAP7_75t_L g603 ( 
.A(n_432),
.B(n_359),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_595),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_531),
.B(n_431),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_526),
.B(n_440),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_477),
.A2(n_461),
.B1(n_431),
.B2(n_434),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_569),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_487),
.B(n_456),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_469),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_514),
.B(n_458),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_528),
.B(n_458),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_478),
.Y(n_615)
);

BUFx6f_ASAP7_75t_SL g616 ( 
.A(n_511),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_494),
.B(n_336),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_477),
.B(n_458),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_477),
.A2(n_440),
.B1(n_461),
.B2(n_455),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_508),
.B(n_458),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_595),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_569),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_470),
.A2(n_561),
.B1(n_556),
.B2(n_552),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_579),
.Y(n_626)
);

CKINVDCx11_ASAP7_75t_R g627 ( 
.A(n_462),
.Y(n_627)
);

BUFx12f_ASAP7_75t_SL g628 ( 
.A(n_470),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_508),
.B(n_458),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_571),
.B(n_568),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_531),
.B(n_431),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_584),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_564),
.B(n_458),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_503),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_564),
.B(n_599),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_L g636 ( 
.A(n_471),
.B(n_432),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_599),
.B(n_434),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_473),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_473),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_491),
.B(n_371),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_R g641 ( 
.A(n_471),
.B(n_378),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_474),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_563),
.B(n_379),
.Y(n_644)
);

BUFx8_ASAP7_75t_L g645 ( 
.A(n_574),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_466),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_474),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_601),
.B(n_440),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_571),
.B(n_436),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_571),
.B(n_436),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_584),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_568),
.B(n_436),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_568),
.B(n_439),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_560),
.B(n_439),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_585),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_475),
.Y(n_656)
);

CKINVDCx16_ASAP7_75t_R g657 ( 
.A(n_542),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_494),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_497),
.B(n_440),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_567),
.B(n_515),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_585),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_470),
.A2(n_442),
.B1(n_449),
.B2(n_448),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_543),
.B(n_442),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_497),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_542),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_475),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_543),
.B(n_448),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_567),
.B(n_525),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_470),
.A2(n_561),
.B1(n_601),
.B2(n_597),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_563),
.B(n_449),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_516),
.B(n_450),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_480),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_492),
.B(n_449),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_513),
.B(n_562),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_516),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_480),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_587),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_570),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_590),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_498),
.B(n_450),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_601),
.B(n_425),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_604),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_543),
.B(n_425),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_557),
.B(n_425),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_557),
.B(n_425),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_465),
.B(n_244),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_604),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_601),
.B(n_438),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_565),
.B(n_438),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_536),
.A2(n_459),
.B(n_438),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_465),
.Y(n_692)
);

NOR2x2_ASAP7_75t_L g693 ( 
.A(n_566),
.B(n_459),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_590),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_570),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_562),
.B(n_459),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_566),
.A2(n_259),
.B1(n_459),
.B2(n_222),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_496),
.B(n_424),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_583),
.B(n_424),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_557),
.B(n_424),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_589),
.A2(n_311),
.B1(n_278),
.B2(n_279),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_561),
.A2(n_226),
.B1(n_247),
.B2(n_187),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_561),
.A2(n_226),
.B1(n_247),
.B2(n_187),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_583),
.B(n_573),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_572),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_573),
.B(n_278),
.Y(n_706)
);

BUFx5_ASAP7_75t_L g707 ( 
.A(n_598),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_592),
.B(n_161),
.Y(n_708)
);

INVxp33_ASAP7_75t_L g709 ( 
.A(n_594),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_589),
.A2(n_279),
.B1(n_286),
.B2(n_312),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_558),
.B(n_269),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_588),
.B(n_422),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_572),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_511),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_588),
.B(n_286),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_509),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_588),
.B(n_422),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_581),
.B(n_422),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_598),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_597),
.A2(n_247),
.B1(n_226),
.B2(n_280),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_468),
.B(n_290),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_600),
.B(n_272),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_581),
.B(n_422),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_509),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_481),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_559),
.B(n_273),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_582),
.B(n_422),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_481),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_558),
.B(n_275),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_483),
.Y(n_731)
);

INVx3_ASAP7_75t_R g732 ( 
.A(n_524),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_540),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_577),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_566),
.A2(n_161),
.B1(n_280),
.B2(n_187),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_566),
.A2(n_576),
.B1(n_488),
.B2(n_540),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_483),
.B(n_276),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_576),
.A2(n_283),
.B1(n_315),
.B2(n_186),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_586),
.B(n_422),
.Y(n_739)
);

NAND2x1_ASAP7_75t_L g740 ( 
.A(n_466),
.B(n_468),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_524),
.B(n_282),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_486),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_468),
.B(n_290),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_482),
.B(n_287),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_591),
.B(n_391),
.Y(n_745)
);

INVxp33_ASAP7_75t_L g746 ( 
.A(n_489),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_580),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_486),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_493),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_484),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_553),
.B(n_391),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_493),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_504),
.B(n_288),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_580),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_SL g755 ( 
.A(n_512),
.B(n_294),
.C(n_289),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_502),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_483),
.B(n_395),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_485),
.B(n_395),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_502),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_506),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_484),
.B(n_299),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_484),
.B(n_302),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_506),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_519),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_511),
.B(n_280),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_501),
.B(n_395),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_519),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_522),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_679),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_641),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_634),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_645),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_671),
.B(n_576),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_722),
.B(n_576),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_704),
.A2(n_613),
.B(n_612),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_682),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_690),
.A2(n_523),
.B(n_537),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_609),
.Y(n_778)
);

AOI21x1_ASAP7_75t_L g779 ( 
.A1(n_652),
.A2(n_467),
.B(n_464),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_623),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_696),
.B(n_463),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_646),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_614),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_665),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_624),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_681),
.B(n_527),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_657),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_741),
.A2(n_593),
.B(n_602),
.C(n_596),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_709),
.B(n_537),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_707),
.B(n_522),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_649),
.A2(n_578),
.B(n_575),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_675),
.B(n_603),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_674),
.B(n_518),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_650),
.A2(n_476),
.B(n_472),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_635),
.B(n_521),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_648),
.B(n_535),
.Y(n_796)
);

NOR2x2_ASAP7_75t_L g797 ( 
.A(n_627),
.B(n_489),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_626),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_614),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_646),
.Y(n_800)
);

OAI321xp33_ASAP7_75t_L g801 ( 
.A1(n_708),
.A2(n_212),
.A3(n_315),
.B1(n_214),
.B2(n_222),
.C(n_225),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_650),
.A2(n_495),
.B(n_479),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_545),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_709),
.B(n_603),
.Y(n_804)
);

OAI321xp33_ASAP7_75t_L g805 ( 
.A1(n_670),
.A2(n_283),
.A3(n_308),
.B1(n_197),
.B2(n_195),
.C(n_193),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_692),
.B(n_466),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_676),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_632),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_712),
.A2(n_495),
.B(n_479),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_629),
.B(n_593),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_618),
.A2(n_466),
.B1(n_546),
.B2(n_535),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_717),
.A2(n_610),
.B(n_684),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_707),
.B(n_538),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_654),
.B(n_636),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_645),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_695),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_634),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_672),
.B(n_538),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_660),
.B(n_546),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_685),
.A2(n_500),
.B(n_499),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_628),
.B(n_547),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_611),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_685),
.A2(n_500),
.B(n_499),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_662),
.A2(n_547),
.B1(n_548),
.B2(n_490),
.Y(n_825)
);

OAI21xp33_ASAP7_75t_L g826 ( 
.A1(n_761),
.A2(n_307),
.B(n_305),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_686),
.A2(n_507),
.B(n_505),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_652),
.A2(n_517),
.B(n_510),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_615),
.B(n_548),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_658),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_663),
.A2(n_517),
.B(n_510),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_669),
.B(n_490),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_620),
.B(n_490),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_651),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_625),
.A2(n_541),
.B1(n_549),
.B2(n_551),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_640),
.A2(n_313),
.B1(n_192),
.B2(n_183),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_617),
.Y(n_837)
);

OAI21xp33_ASAP7_75t_L g838 ( 
.A1(n_762),
.A2(n_726),
.B(n_744),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_695),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_711),
.A2(n_555),
.B1(n_520),
.B2(n_551),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_663),
.A2(n_529),
.B(n_520),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_668),
.A2(n_555),
.B(n_529),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_659),
.B(n_541),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_705),
.Y(n_844)
);

AOI21x1_ASAP7_75t_L g845 ( 
.A1(n_653),
.A2(n_530),
.B(n_550),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_668),
.A2(n_533),
.B(n_550),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_628),
.B(n_541),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_707),
.B(n_549),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_707),
.B(n_731),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_627),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_700),
.A2(n_631),
.B(n_606),
.Y(n_851)
);

AO21x2_ASAP7_75t_L g852 ( 
.A1(n_691),
.A2(n_413),
.B(n_534),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_750),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_699),
.A2(n_661),
.B(n_655),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_666),
.Y(n_855)
);

AND2x2_ASAP7_75t_SL g856 ( 
.A(n_737),
.B(n_296),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_633),
.A2(n_637),
.B(n_743),
.C(n_721),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_606),
.A2(n_532),
.B(n_530),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_664),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_619),
.B(n_549),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_648),
.B(n_532),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_676),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_705),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_608),
.A2(n_413),
.B(n_192),
.C(n_193),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_SL g865 ( 
.A(n_714),
.B(n_195),
.C(n_197),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_707),
.B(n_554),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_634),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_678),
.A2(n_533),
.B(n_544),
.Y(n_868)
);

NOR2x1p5_ASAP7_75t_L g869 ( 
.A(n_714),
.B(n_212),
.Y(n_869)
);

AO21x1_ASAP7_75t_L g870 ( 
.A1(n_631),
.A2(n_312),
.B(n_311),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_721),
.A2(n_202),
.B(n_308),
.C(n_252),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_680),
.A2(n_544),
.B(n_539),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_648),
.B(n_534),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_SL g874 ( 
.A(n_644),
.B(n_214),
.C(n_225),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_713),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_718),
.A2(n_728),
.B(n_723),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_607),
.B(n_687),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_694),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_739),
.A2(n_539),
.B(n_554),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_630),
.A2(n_413),
.B(n_404),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_682),
.B(n_252),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_682),
.B(n_261),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_630),
.A2(n_390),
.B(n_404),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_713),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_719),
.A2(n_390),
.B(n_404),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_740),
.A2(n_390),
.B(n_410),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_727),
.A2(n_296),
.B(n_410),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_746),
.B(n_261),
.Y(n_888)
);

OR2x6_ASAP7_75t_L g889 ( 
.A(n_619),
.B(n_285),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_751),
.A2(n_763),
.B(n_756),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_689),
.B(n_285),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_756),
.A2(n_390),
.B(n_410),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_725),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_727),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_763),
.A2(n_160),
.B(n_168),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_634),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_764),
.A2(n_251),
.B(n_172),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_698),
.A2(n_418),
.B(n_417),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_764),
.A2(n_254),
.B(n_179),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_689),
.B(n_293),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_689),
.B(n_750),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_707),
.B(n_201),
.Y(n_903)
);

AND2x2_ASAP7_75t_SL g904 ( 
.A(n_737),
.B(n_293),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_734),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_743),
.A2(n_418),
.B(n_417),
.C(n_411),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_706),
.A2(n_418),
.B(n_399),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_716),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_765),
.B(n_399),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_707),
.B(n_408),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_715),
.A2(n_399),
.B(n_411),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_767),
.A2(n_246),
.B(n_182),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_767),
.A2(n_248),
.B(n_191),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_729),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_732),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_753),
.B(n_401),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_605),
.A2(n_200),
.B1(n_409),
.B2(n_401),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_616),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_716),
.B(n_408),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_736),
.B(n_407),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_711),
.B(n_730),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_768),
.A2(n_255),
.B(n_198),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_730),
.B(n_407),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_768),
.A2(n_258),
.B(n_199),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_716),
.B(n_408),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_701),
.A2(n_171),
.B(n_310),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_720),
.B(n_409),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_755),
.B(n_204),
.C(n_210),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_746),
.B(n_6),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_745),
.A2(n_264),
.B(n_213),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_742),
.A2(n_267),
.B(n_219),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_605),
.B(n_224),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_748),
.A2(n_277),
.B(n_227),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_605),
.B(n_229),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_619),
.B(n_284),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_749),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_643),
.B(n_622),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_622),
.B(n_233),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_734),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_616),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_757),
.A2(n_752),
.B(n_760),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_758),
.A2(n_400),
.B(n_414),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_747),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_738),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_622),
.B(n_234),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_747),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_645),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_759),
.A2(n_297),
.B(n_242),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_735),
.B(n_8),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_775),
.A2(n_851),
.B(n_813),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_838),
.A2(n_697),
.B(n_688),
.C(n_683),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_776),
.B(n_643),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_778),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_876),
.A2(n_683),
.B(n_688),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_776),
.B(n_643),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_780),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_SL g957 ( 
.A1(n_789),
.A2(n_688),
.B(n_683),
.C(n_638),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_776),
.B(n_716),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_856),
.A2(n_710),
.B1(n_703),
.B2(n_702),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_803),
.B(n_638),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_784),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_792),
.B(n_639),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_772),
.B(n_724),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_796),
.B(n_724),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_770),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_785),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_837),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_771),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_910),
.A2(n_766),
.B(n_724),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_774),
.A2(n_656),
.B(n_639),
.C(n_677),
.Y(n_970)
);

NOR2xp67_ASAP7_75t_SL g971 ( 
.A(n_807),
.B(n_733),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_910),
.A2(n_733),
.B(n_724),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_777),
.A2(n_733),
.B(n_647),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_798),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_770),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_904),
.A2(n_667),
.B(n_642),
.C(n_677),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_773),
.A2(n_673),
.B(n_754),
.C(n_693),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_904),
.A2(n_673),
.B(n_754),
.C(n_271),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_771),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_804),
.B(n_616),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_807),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_866),
.A2(n_298),
.B(n_292),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_866),
.A2(n_414),
.B(n_408),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_SL g984 ( 
.A1(n_789),
.A2(n_9),
.B(n_10),
.C(n_16),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_808),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_830),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_SL g987 ( 
.A1(n_836),
.A2(n_175),
.B1(n_18),
.B2(n_19),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_862),
.B(n_17),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_769),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_858),
.A2(n_848),
.B(n_814),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_817),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_862),
.B(n_18),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_859),
.B(n_21),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_787),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_856),
.B(n_806),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_806),
.B(n_414),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_788),
.A2(n_921),
.B(n_786),
.C(n_857),
.Y(n_997)
);

OAI21xp33_ASAP7_75t_SL g998 ( 
.A1(n_902),
.A2(n_25),
.B(n_26),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_834),
.Y(n_999)
);

INVx3_ASAP7_75t_SL g1000 ( 
.A(n_797),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_848),
.A2(n_414),
.B(n_408),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_877),
.B(n_25),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_788),
.A2(n_874),
.B(n_815),
.C(n_826),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_944),
.B(n_29),
.C(n_32),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_781),
.B(n_29),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_801),
.B(n_935),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_855),
.Y(n_1007)
);

OAI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_865),
.A2(n_175),
.B(n_33),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_823),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_888),
.B(n_32),
.Y(n_1010)
);

BUFx12f_ASAP7_75t_L g1011 ( 
.A(n_823),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_796),
.B(n_33),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_772),
.Y(n_1013)
);

BUFx8_ASAP7_75t_SL g1014 ( 
.A(n_816),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_811),
.A2(n_175),
.B1(n_35),
.B2(n_38),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_878),
.A2(n_175),
.B1(n_38),
.B2(n_39),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_949),
.A2(n_400),
.B1(n_414),
.B2(n_408),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_790),
.A2(n_414),
.B(n_408),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_790),
.A2(n_414),
.B(n_408),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_843),
.A2(n_34),
.B(n_42),
.C(n_43),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_854),
.A2(n_414),
.B(n_44),
.C(n_45),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_929),
.A2(n_400),
.B1(n_45),
.B2(n_46),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_892),
.B(n_42),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_889),
.B(n_50),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_928),
.A2(n_54),
.B(n_56),
.C(n_59),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_800),
.B(n_117),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_816),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_791),
.A2(n_59),
.B(n_400),
.C(n_79),
.Y(n_1028)
);

INVx6_ASAP7_75t_SL g1029 ( 
.A(n_889),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_915),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_947),
.B(n_78),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_800),
.B(n_400),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_894),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_914),
.Y(n_1034)
);

O2A1O1Ixp5_ASAP7_75t_L g1035 ( 
.A1(n_903),
.A2(n_400),
.B(n_85),
.C(n_92),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_800),
.B(n_400),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_936),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_869),
.B(n_400),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_947),
.B(n_83),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_796),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_793),
.B(n_100),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_881),
.B(n_103),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_839),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_797),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_SL g1045 ( 
.A1(n_919),
.A2(n_925),
.B(n_903),
.C(n_849),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_814),
.A2(n_104),
.B(n_108),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_822),
.B(n_847),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_871),
.A2(n_937),
.B(n_822),
.C(n_916),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_833),
.A2(n_114),
.B1(n_120),
.B2(n_129),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_861),
.A2(n_130),
.B1(n_135),
.B2(n_138),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_873),
.A2(n_141),
.B1(n_147),
.B2(n_149),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_850),
.Y(n_1052)
);

AND2x6_ASAP7_75t_L g1053 ( 
.A(n_782),
.B(n_155),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_795),
.A2(n_159),
.B1(n_864),
.B2(n_901),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_771),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_882),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_844),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_891),
.B(n_918),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_819),
.A2(n_812),
.B(n_945),
.C(n_938),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_937),
.A2(n_941),
.B(n_847),
.C(n_868),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_863),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_820),
.B(n_863),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_SL g1063 ( 
.A1(n_849),
.A2(n_872),
.B(n_934),
.C(n_932),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_SL g1064 ( 
.A(n_800),
.B(n_782),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_840),
.A2(n_805),
.B(n_832),
.C(n_890),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_783),
.B(n_799),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_783),
.B(n_799),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_829),
.B(n_771),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_923),
.A2(n_926),
.B(n_906),
.C(n_930),
.Y(n_1069)
);

CKINVDCx14_ASAP7_75t_R g1070 ( 
.A(n_940),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_864),
.A2(n_853),
.B1(n_782),
.B2(n_809),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_875),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_SL g1073 ( 
.A1(n_842),
.A2(n_846),
.B(n_824),
.C(n_821),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_875),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_810),
.A2(n_879),
.B(n_827),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_818),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_884),
.B(n_939),
.Y(n_1077)
);

AND3x1_ASAP7_75t_SL g1078 ( 
.A(n_931),
.B(n_948),
.C(n_933),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_909),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_896),
.B(n_913),
.C(n_900),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_897),
.A2(n_870),
.B1(n_835),
.B2(n_853),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_897),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_884),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_818),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_794),
.A2(n_802),
.B(n_831),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_841),
.A2(n_880),
.B(n_809),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_L g1087 ( 
.A(n_920),
.B(n_927),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_853),
.A2(n_919),
.B(n_925),
.C(n_825),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_895),
.A2(n_946),
.B1(n_943),
.B2(n_939),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_905),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_905),
.B(n_943),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1086),
.A2(n_942),
.B(n_887),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_950),
.A2(n_887),
.B(n_899),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_997),
.A2(n_809),
.B(n_885),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_963),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_SL g1096 ( 
.A1(n_1015),
.A2(n_1016),
.B(n_1066),
.C(n_1049),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_SL g1097 ( 
.A1(n_1015),
.A2(n_1016),
.B(n_1049),
.C(n_1054),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_1089),
.A2(n_917),
.A3(n_883),
.B(n_893),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_964),
.B(n_867),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_994),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1029),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1029),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1041),
.A2(n_886),
.B(n_852),
.Y(n_1103)
);

OAI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1000),
.A2(n_779),
.B1(n_845),
.B2(n_828),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_959),
.A2(n_818),
.B1(n_908),
.B2(n_867),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_1011),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_964),
.B(n_818),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_1054),
.A2(n_924),
.A3(n_922),
.B(n_912),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_961),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_975),
.Y(n_1110)
);

AO22x1_ASAP7_75t_L g1111 ( 
.A1(n_959),
.A2(n_908),
.B1(n_867),
.B2(n_911),
.Y(n_1111)
);

OAI22x1_ASAP7_75t_L g1112 ( 
.A1(n_1024),
.A2(n_860),
.B1(n_867),
.B2(n_908),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_962),
.B(n_980),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1060),
.A2(n_907),
.B(n_898),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1045),
.A2(n_852),
.B(n_1065),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1010),
.B(n_988),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1041),
.A2(n_1063),
.B(n_1088),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1047),
.B(n_967),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1003),
.A2(n_1008),
.B(n_978),
.C(n_1005),
.Y(n_1119)
);

AO32x2_ASAP7_75t_L g1120 ( 
.A1(n_987),
.A2(n_1071),
.A3(n_1050),
.B1(n_1051),
.B2(n_984),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_963),
.B(n_1013),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1056),
.B(n_986),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1048),
.A2(n_1069),
.B(n_969),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1004),
.A2(n_1025),
.B(n_1021),
.C(n_992),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_954),
.A2(n_1085),
.B(n_973),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_995),
.A2(n_1006),
.B1(n_1012),
.B2(n_993),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_1052),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1059),
.A2(n_990),
.B(n_1073),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1012),
.A2(n_1002),
.B1(n_1022),
.B2(n_1079),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1071),
.A2(n_960),
.B(n_972),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_960),
.A2(n_957),
.B(n_996),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1009),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_983),
.A2(n_1018),
.B(n_1019),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_963),
.B(n_1013),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_968),
.B(n_979),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1027),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1076),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_951),
.A2(n_1081),
.B(n_976),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1080),
.A2(n_1042),
.B(n_1062),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_977),
.A2(n_1020),
.B(n_1087),
.C(n_970),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1044),
.B(n_1023),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_956),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1062),
.A2(n_1028),
.B(n_1046),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1001),
.A2(n_1051),
.B(n_1050),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_966),
.A2(n_1007),
.B1(n_999),
.B2(n_985),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1014),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1032),
.A2(n_1036),
.B(n_1084),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1058),
.A2(n_981),
.B1(n_1030),
.B2(n_974),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1017),
.A2(n_998),
.B(n_1037),
.C(n_1035),
.Y(n_1150)
);

OAI22x1_ASAP7_75t_L g1151 ( 
.A1(n_1038),
.A2(n_1067),
.B1(n_965),
.B2(n_1068),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_952),
.A2(n_955),
.B(n_1082),
.C(n_982),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1067),
.A2(n_1070),
.B(n_1026),
.C(n_958),
.Y(n_1153)
);

AO32x2_ASAP7_75t_L g1154 ( 
.A1(n_965),
.A2(n_1078),
.A3(n_1090),
.B1(n_1083),
.B2(n_1072),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1026),
.A2(n_1091),
.B(n_1077),
.Y(n_1155)
);

CKINVDCx6p67_ASAP7_75t_R g1156 ( 
.A(n_1053),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_968),
.A2(n_1055),
.B(n_979),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_968),
.A2(n_1055),
.B(n_979),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_971),
.A2(n_1064),
.B(n_989),
.C(n_991),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1055),
.B(n_1043),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_R g1161 ( 
.A(n_1031),
.B(n_1039),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_958),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1057),
.A2(n_1074),
.B(n_1061),
.C(n_1053),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1053),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1053),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1053),
.A2(n_838),
.B(n_950),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1012),
.A2(n_904),
.B1(n_856),
.B2(n_773),
.Y(n_1167)
);

INVxp67_ASAP7_75t_SL g1168 ( 
.A(n_1040),
.Y(n_1168)
);

OAI22x1_ASAP7_75t_L g1169 ( 
.A1(n_1000),
.A2(n_489),
.B1(n_640),
.B2(n_1024),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1086),
.A2(n_950),
.B(n_1075),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1003),
.A2(n_838),
.B(n_722),
.C(n_856),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1086),
.A2(n_950),
.B(n_1075),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_958),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_961),
.B(n_792),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_981),
.B(n_709),
.Y(n_1175)
);

BUFx8_ASAP7_75t_L g1176 ( 
.A(n_975),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_975),
.Y(n_1177)
);

INVxp67_ASAP7_75t_SL g1178 ( 
.A(n_1040),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1089),
.A2(n_997),
.A3(n_1054),
.B(n_1065),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_967),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1047),
.B(n_904),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1011),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_962),
.B(n_792),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1024),
.A2(n_722),
.B(n_988),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1003),
.A2(n_838),
.B(n_722),
.C(n_856),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1003),
.A2(n_838),
.B(n_722),
.C(n_856),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_961),
.B(n_792),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_967),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_1003),
.A2(n_722),
.B(n_838),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1086),
.A2(n_950),
.B(n_1075),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1015),
.A2(n_722),
.B(n_838),
.C(n_709),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_SL g1197 ( 
.A1(n_997),
.A2(n_921),
.B(n_838),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_962),
.B(n_877),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_959),
.A2(n_470),
.B1(n_709),
.B2(n_765),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1003),
.A2(n_838),
.B(n_722),
.C(n_856),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_994),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_963),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1086),
.A2(n_950),
.B(n_1075),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1086),
.A2(n_950),
.B(n_1075),
.Y(n_1204)
);

CKINVDCx11_ASAP7_75t_R g1205 ( 
.A(n_994),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_962),
.B(n_877),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_1003),
.B(n_838),
.C(n_722),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1089),
.A2(n_997),
.A3(n_1054),
.B(n_1065),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_950),
.B(n_1075),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1003),
.A2(n_838),
.B(n_722),
.C(n_856),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1089),
.A2(n_997),
.A3(n_1054),
.B(n_1065),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_1060),
.B(n_838),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1003),
.A2(n_838),
.B(n_722),
.C(n_856),
.Y(n_1215)
);

NOR4xp25_ASAP7_75t_L g1216 ( 
.A(n_959),
.B(n_838),
.C(n_1016),
.D(n_1015),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_953),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_962),
.B(n_877),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_950),
.A2(n_838),
.B(n_997),
.Y(n_1219)
);

NOR2xp67_ASAP7_75t_SL g1220 ( 
.A(n_975),
.B(n_542),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_962),
.B(n_877),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_994),
.Y(n_1222)
);

AO32x2_ASAP7_75t_L g1223 ( 
.A1(n_1015),
.A2(n_1016),
.A3(n_959),
.B1(n_1054),
.B2(n_987),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_962),
.B(n_792),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_950),
.A2(n_1086),
.B(n_1075),
.Y(n_1225)
);

BUFx10_ASAP7_75t_L g1226 ( 
.A(n_981),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_1003),
.B(n_838),
.C(n_722),
.Y(n_1227)
);

AOI221xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1015),
.A2(n_1016),
.B1(n_1008),
.B2(n_944),
.C(n_788),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_1054),
.A2(n_1015),
.B(n_1003),
.Y(n_1229)
);

NOR4xp25_ASAP7_75t_L g1230 ( 
.A(n_959),
.B(n_838),
.C(n_1016),
.D(n_1015),
.Y(n_1230)
);

NOR2x1_ASAP7_75t_SL g1231 ( 
.A(n_963),
.B(n_968),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_997),
.A2(n_1060),
.B(n_1045),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1073),
.A2(n_630),
.B(n_838),
.C(n_1060),
.Y(n_1233)
);

BUFx2_ASAP7_75t_SL g1234 ( 
.A(n_994),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_962),
.B(n_877),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1137),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1165),
.B(n_1095),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1205),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1167),
.A2(n_1116),
.B1(n_1227),
.B2(n_1207),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1149),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1167),
.A2(n_1207),
.B1(n_1227),
.B2(n_1129),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1109),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1222),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1169),
.A2(n_1199),
.B1(n_1229),
.B2(n_1182),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1095),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1226),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1187),
.B(n_1118),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_SL g1248 ( 
.A(n_1146),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1226),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1171),
.A2(n_1190),
.B(n_1188),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1145),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1186),
.A2(n_1224),
.B1(n_1193),
.B2(n_1213),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1187),
.A2(n_1215),
.B1(n_1200),
.B2(n_1211),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1126),
.A2(n_1191),
.B1(n_1174),
.B2(n_1141),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1175),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1121),
.Y(n_1256)
);

INVx6_ASAP7_75t_L g1257 ( 
.A(n_1095),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1126),
.A2(n_1196),
.B1(n_1124),
.B2(n_1119),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1113),
.A2(n_1235),
.B1(n_1198),
.B2(n_1206),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1218),
.A2(n_1221),
.B1(n_1138),
.B2(n_1223),
.Y(n_1260)
);

CKINVDCx11_ASAP7_75t_R g1261 ( 
.A(n_1201),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1180),
.B(n_1192),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1138),
.A2(n_1223),
.B1(n_1165),
.B2(n_1156),
.Y(n_1263)
);

CKINVDCx8_ASAP7_75t_R g1264 ( 
.A(n_1234),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_SL g1265 ( 
.A(n_1127),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1100),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1105),
.A2(n_1165),
.B1(n_1148),
.B2(n_1122),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1181),
.A2(n_1189),
.B(n_1209),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1121),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1145),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1106),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1155),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1223),
.A2(n_1164),
.B1(n_1216),
.B2(n_1230),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1142),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1176),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1217),
.Y(n_1276)
);

INVx5_ASAP7_75t_L g1277 ( 
.A(n_1164),
.Y(n_1277)
);

BUFx10_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1134),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1099),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_L g1281 ( 
.A(n_1134),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1144),
.A2(n_1195),
.B(n_1214),
.Y(n_1282)
);

BUFx2_ASAP7_75t_SL g1283 ( 
.A(n_1110),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1232),
.A2(n_1105),
.B1(n_1230),
.B2(n_1216),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1154),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1232),
.A2(n_1192),
.B1(n_1180),
.B2(n_1168),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1178),
.A2(n_1228),
.B1(n_1114),
.B2(n_1123),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1099),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1132),
.B(n_1161),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1202),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1228),
.A2(n_1114),
.B1(n_1123),
.B2(n_1219),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1154),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1184),
.A2(n_1185),
.B1(n_1197),
.B2(n_1150),
.Y(n_1293)
);

BUFx2_ASAP7_75t_R g1294 ( 
.A(n_1183),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1107),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1177),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1202),
.B(n_1173),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1166),
.A2(n_1117),
.B(n_1153),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1101),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1154),
.Y(n_1300)
);

INVx8_ASAP7_75t_L g1301 ( 
.A(n_1160),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1115),
.A2(n_1102),
.B1(n_1220),
.B2(n_1112),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1176),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1177),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1231),
.A2(n_1202),
.B1(n_1097),
.B2(n_1096),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1140),
.A2(n_1094),
.B1(n_1128),
.B2(n_1131),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1115),
.A2(n_1151),
.B1(n_1139),
.B2(n_1104),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1162),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1162),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1162),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1159),
.A2(n_1143),
.B1(n_1152),
.B2(n_1130),
.Y(n_1311)
);

INVx8_ASAP7_75t_L g1312 ( 
.A(n_1173),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1107),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1111),
.A2(n_1120),
.B1(n_1212),
.B2(n_1179),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1120),
.A2(n_1163),
.B(n_1233),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1135),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1135),
.B(n_1120),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1179),
.Y(n_1318)
);

BUFx4f_ASAP7_75t_SL g1319 ( 
.A(n_1157),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1147),
.A2(n_1179),
.B1(n_1208),
.B2(n_1212),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1208),
.A2(n_1212),
.B1(n_1103),
.B2(n_1225),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1208),
.A2(n_1108),
.B1(n_1225),
.B2(n_1158),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1108),
.A2(n_1172),
.B1(n_1204),
.B2(n_1203),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1093),
.A2(n_1125),
.B1(n_1133),
.B2(n_1092),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1170),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1108),
.A2(n_1194),
.B1(n_1210),
.B2(n_1098),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1098),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1098),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1205),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1226),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1149),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1149),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1118),
.B(n_1116),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1149),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1127),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1167),
.A2(n_804),
.B1(n_904),
.B2(n_489),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1169),
.A2(n_470),
.B1(n_462),
.B2(n_836),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1167),
.A2(n_804),
.B1(n_904),
.B2(n_489),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1137),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1187),
.A2(n_1116),
.B1(n_904),
.B2(n_856),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1137),
.Y(n_1341)
);

AO22x1_ASAP7_75t_L g1342 ( 
.A1(n_1116),
.A2(n_640),
.B1(n_1024),
.B2(n_959),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1095),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1167),
.A2(n_856),
.B1(n_904),
.B2(n_640),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1167),
.A2(n_804),
.B1(n_904),
.B2(n_489),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1118),
.B(n_1116),
.Y(n_1346)
);

BUFx8_ASAP7_75t_SL g1347 ( 
.A(n_1146),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1109),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1149),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1187),
.A2(n_1116),
.B1(n_904),
.B2(n_856),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1187),
.A2(n_1116),
.B1(n_640),
.B2(n_1199),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1167),
.A2(n_804),
.B1(n_904),
.B2(n_489),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1118),
.B(n_1116),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1187),
.A2(n_1116),
.B1(n_904),
.B2(n_856),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1205),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1137),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1167),
.A2(n_804),
.B1(n_904),
.B2(n_489),
.Y(n_1357)
);

BUFx4_ASAP7_75t_SL g1358 ( 
.A(n_1146),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1149),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1187),
.A2(n_1116),
.B1(n_640),
.B2(n_1199),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1167),
.A2(n_856),
.B1(n_904),
.B2(n_640),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1205),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1167),
.A2(n_804),
.B1(n_904),
.B2(n_489),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1167),
.A2(n_856),
.B1(n_904),
.B2(n_640),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1251),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1270),
.B(n_1285),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1260),
.B(n_1273),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1282),
.A2(n_1326),
.B(n_1311),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1274),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1261),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1274),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1324),
.A2(n_1306),
.B(n_1293),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1285),
.B(n_1292),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1292),
.B(n_1300),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1320),
.A2(n_1268),
.B(n_1328),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1276),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1300),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1318),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1318),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1340),
.A2(n_1350),
.B1(n_1354),
.B2(n_1360),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1348),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1327),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1347),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1317),
.B(n_1284),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1272),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1325),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1255),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1258),
.A2(n_1351),
.B(n_1344),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1291),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1260),
.B(n_1287),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1284),
.B(n_1247),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1247),
.B(n_1314),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1361),
.A2(n_1364),
.B(n_1291),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1240),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1287),
.B(n_1263),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1339),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1324),
.A2(n_1321),
.B(n_1298),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1277),
.B(n_1256),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1256),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1336),
.A2(n_1363),
.B1(n_1338),
.B2(n_1357),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1331),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1332),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1336),
.A2(n_1363),
.B(n_1345),
.C(n_1357),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1277),
.B(n_1279),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1334),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1349),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1359),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1250),
.A2(n_1253),
.B(n_1315),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1263),
.B(n_1321),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1262),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1277),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1322),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1239),
.B(n_1307),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1313),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1356),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1319),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1319),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1255),
.B(n_1289),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1241),
.A2(n_1244),
.B(n_1352),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1323),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1356),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1286),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1286),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1269),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1316),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1305),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1252),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1236),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1252),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1341),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1338),
.A2(n_1352),
.B1(n_1345),
.B2(n_1342),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1267),
.A2(n_1244),
.B(n_1302),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1302),
.A2(n_1254),
.B(n_1259),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1254),
.B(n_1259),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1299),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1398),
.B(n_1288),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1398),
.B(n_1278),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1390),
.A2(n_1246),
.B(n_1249),
.C(n_1330),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1393),
.B(n_1290),
.Y(n_1441)
);

OAI211xp5_ASAP7_75t_L g1442 ( 
.A1(n_1410),
.A2(n_1264),
.B(n_1266),
.C(n_1296),
.Y(n_1442)
);

OAI211xp5_ASAP7_75t_L g1443 ( 
.A1(n_1390),
.A2(n_1421),
.B(n_1393),
.C(n_1415),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1370),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1421),
.A2(n_1337),
.B1(n_1271),
.B2(n_1283),
.C(n_1335),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1433),
.A2(n_1280),
.B1(n_1281),
.B2(n_1303),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1380),
.A2(n_1275),
.B(n_1358),
.C(n_1248),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1405),
.A2(n_1335),
.B1(n_1304),
.B2(n_1296),
.C(n_1355),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_L g1449 ( 
.A(n_1418),
.B(n_1362),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1433),
.A2(n_1281),
.B1(n_1294),
.B2(n_1243),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1395),
.A2(n_1237),
.B(n_1297),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1391),
.B(n_1290),
.Y(n_1452)
);

OAI211xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1381),
.A2(n_1382),
.B(n_1430),
.C(n_1417),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_SL g1454 ( 
.A1(n_1384),
.A2(n_1423),
.B(n_1395),
.C(n_1437),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1386),
.B(n_1238),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1386),
.B(n_1329),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1309),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1391),
.B(n_1295),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1366),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1426),
.B(n_1295),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1412),
.B(n_1301),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1401),
.B(n_1265),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1366),
.B(n_1308),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1415),
.A2(n_1237),
.B(n_1312),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1392),
.A2(n_1312),
.B(n_1265),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_L g1466 ( 
.A(n_1420),
.B(n_1248),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1399),
.A2(n_1368),
.B(n_1372),
.Y(n_1467)
);

NAND4xp25_ASAP7_75t_L g1468 ( 
.A(n_1394),
.B(n_1310),
.C(n_1312),
.D(n_1245),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1365),
.B(n_1308),
.Y(n_1469)
);

AO32x2_ASAP7_75t_L g1470 ( 
.A1(n_1373),
.A2(n_1257),
.A3(n_1308),
.B1(n_1343),
.B2(n_1374),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1396),
.B(n_1257),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1367),
.A2(n_1343),
.B1(n_1435),
.B2(n_1394),
.Y(n_1472)
);

AO32x2_ASAP7_75t_L g1473 ( 
.A1(n_1373),
.A2(n_1343),
.A3(n_1374),
.B1(n_1425),
.B2(n_1424),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1396),
.B(n_1403),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1432),
.B(n_1389),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1401),
.B(n_1400),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1432),
.B(n_1404),
.Y(n_1477)
);

BUFx8_ASAP7_75t_SL g1478 ( 
.A(n_1370),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1418),
.A2(n_1419),
.B(n_1388),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1402),
.A2(n_1367),
.B1(n_1435),
.B2(n_1397),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1428),
.A2(n_1431),
.B(n_1429),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1434),
.A2(n_1436),
.B1(n_1431),
.B2(n_1429),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1365),
.B(n_1376),
.Y(n_1483)
);

OAI21xp33_ASAP7_75t_L g1484 ( 
.A1(n_1422),
.A2(n_1428),
.B(n_1424),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1369),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1422),
.A2(n_1414),
.B(n_1425),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1370),
.B(n_1385),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1436),
.A2(n_1411),
.B(n_1414),
.C(n_1418),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1408),
.B(n_1409),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_SL g1490 ( 
.A(n_1413),
.B(n_1434),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1467),
.B(n_1375),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1485),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1470),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_1375),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1483),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1483),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1459),
.Y(n_1497)
);

AND2x2_ASAP7_75t_SL g1498 ( 
.A(n_1476),
.B(n_1411),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1479),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1375),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1444),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1474),
.Y(n_1502)
);

AND2x2_ASAP7_75t_SL g1503 ( 
.A(n_1476),
.B(n_1406),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1477),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1489),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1470),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1470),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1480),
.A2(n_1434),
.B1(n_1427),
.B2(n_1407),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1469),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1473),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1490),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1458),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1458),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1452),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1463),
.B(n_1377),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1480),
.A2(n_1427),
.B1(n_1407),
.B2(n_1383),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1463),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1482),
.B(n_1383),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1452),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1445),
.A2(n_1379),
.B1(n_1378),
.B2(n_1416),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1496),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1508),
.A2(n_1443),
.B(n_1488),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1492),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1493),
.B(n_1438),
.Y(n_1526)
);

OAI322xp33_ASAP7_75t_L g1527 ( 
.A1(n_1519),
.A2(n_1472),
.A3(n_1450),
.B1(n_1440),
.B2(n_1487),
.C1(n_1441),
.C2(n_1446),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1491),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1499),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1493),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1493),
.B(n_1507),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1513),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1514),
.Y(n_1534)
);

INVx5_ASAP7_75t_L g1535 ( 
.A(n_1491),
.Y(n_1535)
);

AND2x2_ASAP7_75t_SL g1536 ( 
.A(n_1498),
.B(n_1486),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1508),
.A2(n_1448),
.B1(n_1450),
.B2(n_1445),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1492),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1517),
.A2(n_1448),
.B1(n_1484),
.B2(n_1481),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1491),
.A2(n_1481),
.B(n_1379),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1517),
.A2(n_1500),
.B1(n_1511),
.B2(n_1519),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1494),
.B(n_1454),
.C(n_1447),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1507),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1503),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1441),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1455),
.Y(n_1547)
);

OAI33xp33_ASAP7_75t_L g1548 ( 
.A1(n_1514),
.A2(n_1453),
.A3(n_1471),
.B1(n_1461),
.B2(n_1468),
.B3(n_1371),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1501),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1495),
.B(n_1460),
.Y(n_1550)
);

OAI321xp33_ASAP7_75t_L g1551 ( 
.A1(n_1521),
.A2(n_1451),
.A3(n_1465),
.B1(n_1464),
.B2(n_1442),
.C(n_1456),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1495),
.B(n_1439),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1503),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1498),
.A2(n_1521),
.B1(n_1504),
.B2(n_1503),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1494),
.A2(n_1378),
.B(n_1387),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1499),
.Y(n_1556)
);

INVx5_ASAP7_75t_L g1557 ( 
.A(n_1494),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1510),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1523),
.B(n_1515),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1547),
.Y(n_1561)
);

OR2x6_ASAP7_75t_SL g1562 ( 
.A(n_1542),
.B(n_1512),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1525),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1538),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1553),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1546),
.B(n_1497),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1546),
.B(n_1550),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_1537),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

OAI33xp33_ASAP7_75t_L g1571 ( 
.A1(n_1537),
.A2(n_1506),
.A3(n_1520),
.B1(n_1495),
.B2(n_1505),
.B3(n_1502),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1533),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1555),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1546),
.B(n_1497),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1553),
.B(n_1503),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1504),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1544),
.B(n_1518),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1544),
.B(n_1518),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1531),
.B(n_1478),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1550),
.B(n_1516),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1547),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1520),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1522),
.B(n_1516),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1555),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1555),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1552),
.B(n_1520),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1569),
.A2(n_1524),
.B1(n_1551),
.B2(n_1542),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1569),
.A2(n_1541),
.B(n_1529),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1572),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1573),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1534),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1559),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1573),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1568),
.B(n_1530),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1571),
.A2(n_1524),
.B1(n_1536),
.B2(n_1541),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1535),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1559),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1590),
.B(n_1535),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1590),
.B(n_1535),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1575),
.B(n_1535),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1564),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1566),
.B(n_1535),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1564),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1565),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1561),
.B(n_1522),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1581),
.B(n_1554),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_1531),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1562),
.B(n_1535),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1535),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1543),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1563),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_1543),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1563),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1573),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1535),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1577),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1570),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1576),
.B(n_1535),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1582),
.B(n_1557),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1570),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1577),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1563),
.B(n_1557),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1585),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1578),
.B(n_1557),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1572),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1580),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1587),
.B(n_1567),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1592),
.A2(n_1593),
.B1(n_1600),
.B2(n_1539),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1594),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.B(n_1578),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1597),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1634),
.B(n_1587),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1602),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1595),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1614),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1584),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1614),
.B(n_1579),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1602),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1630),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1630),
.B(n_1579),
.Y(n_1649)
);

AND2x2_ASAP7_75t_SL g1650 ( 
.A(n_1613),
.B(n_1531),
.Y(n_1650)
);

NAND3xp33_ASAP7_75t_L g1651 ( 
.A(n_1593),
.B(n_1539),
.C(n_1529),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1531),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1531),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1634),
.B(n_1558),
.Y(n_1654)
);

NOR3xp33_ASAP7_75t_L g1655 ( 
.A(n_1633),
.B(n_1551),
.C(n_1527),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1606),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1606),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1634),
.B(n_1586),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1596),
.B(n_1567),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1608),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1608),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1609),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1629),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1596),
.B(n_1591),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1560),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1609),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1603),
.B(n_1549),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1612),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1632),
.B(n_1545),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1670)
);

OAI31xp33_ASAP7_75t_L g1671 ( 
.A1(n_1651),
.A2(n_1611),
.A3(n_1554),
.B(n_1556),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1648),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1635),
.A2(n_1655),
.B1(n_1645),
.B2(n_1536),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1665),
.A2(n_1633),
.B(n_1527),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_SL g1675 ( 
.A(n_1636),
.B(n_1637),
.C(n_1654),
.Y(n_1675)
);

OAI21xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1650),
.A2(n_1616),
.B(n_1626),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1649),
.B(n_1632),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1649),
.A2(n_1536),
.B1(n_1540),
.B2(n_1548),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1641),
.B(n_1532),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1667),
.A2(n_1626),
.B(n_1616),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1650),
.A2(n_1616),
.B(n_1626),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1643),
.A2(n_1598),
.B(n_1595),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1641),
.A2(n_1557),
.B1(n_1549),
.B2(n_1536),
.Y(n_1683)
);

NOR4xp25_ASAP7_75t_L g1684 ( 
.A(n_1639),
.B(n_1620),
.C(n_1618),
.D(n_1627),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1659),
.B(n_1610),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1639),
.Y(n_1686)
);

XNOR2xp5_ASAP7_75t_L g1687 ( 
.A(n_1638),
.B(n_1501),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1658),
.B(n_1532),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1644),
.A2(n_1511),
.B(n_1557),
.C(n_1532),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1638),
.B(n_1549),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1659),
.B(n_1532),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1644),
.A2(n_1557),
.B1(n_1549),
.B2(n_1556),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1652),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

AOI31xp33_ASAP7_75t_L g1695 ( 
.A1(n_1652),
.A2(n_1466),
.A3(n_1620),
.B(n_1631),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1664),
.B(n_1532),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1674),
.A2(n_1653),
.B(n_1644),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_L g1698 ( 
.A(n_1675),
.B(n_1653),
.C(n_1660),
.Y(n_1698)
);

AOI32xp33_ASAP7_75t_L g1699 ( 
.A1(n_1683),
.A2(n_1646),
.A3(n_1669),
.B1(n_1556),
.B2(n_1670),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1672),
.B(n_1646),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1685),
.B(n_1670),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1677),
.B(n_1662),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1684),
.B(n_1666),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1687),
.Y(n_1704)
);

INVxp33_ASAP7_75t_L g1705 ( 
.A(n_1690),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_SL g1706 ( 
.A1(n_1671),
.A2(n_1695),
.B(n_1673),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1678),
.A2(n_1588),
.B1(n_1577),
.B2(n_1620),
.C(n_1599),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1686),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1682),
.Y(n_1710)
);

AOI32xp33_ASAP7_75t_L g1711 ( 
.A1(n_1683),
.A2(n_1691),
.A3(n_1679),
.B1(n_1696),
.B2(n_1688),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1693),
.A2(n_1557),
.B1(n_1549),
.B2(n_1663),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1682),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1692),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1680),
.B(n_1667),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1705),
.B(n_1676),
.Y(n_1716)
);

NAND2x1_ASAP7_75t_L g1717 ( 
.A(n_1700),
.B(n_1663),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1701),
.B(n_1610),
.Y(n_1718)
);

AOI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1703),
.A2(n_1643),
.B(n_1642),
.Y(n_1719)
);

AOI222xp33_ASAP7_75t_L g1720 ( 
.A1(n_1697),
.A2(n_1598),
.B1(n_1588),
.B2(n_1589),
.C1(n_1681),
.C2(n_1668),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1713),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1697),
.A2(n_1692),
.B(n_1642),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1703),
.A2(n_1647),
.B(n_1640),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1704),
.A2(n_1501),
.B1(n_1663),
.B2(n_1457),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1706),
.B(n_1699),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1707),
.A2(n_1588),
.B1(n_1589),
.B2(n_1628),
.Y(n_1726)
);

NOR3xp33_ASAP7_75t_SL g1727 ( 
.A(n_1725),
.B(n_1698),
.C(n_1712),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1720),
.A2(n_1710),
.B1(n_1714),
.B2(n_1715),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_L g1729 ( 
.A(n_1719),
.B(n_1709),
.C(n_1708),
.Y(n_1729)
);

AOI222xp33_ASAP7_75t_L g1730 ( 
.A1(n_1721),
.A2(n_1628),
.B1(n_1595),
.B2(n_1621),
.C1(n_1623),
.C2(n_1647),
.Y(n_1730)
);

OAI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1718),
.A2(n_1723),
.B1(n_1722),
.B2(n_1557),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1726),
.A2(n_1623),
.B1(n_1621),
.B2(n_1628),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1716),
.B(n_1702),
.C(n_1711),
.Y(n_1733)
);

NAND4xp25_ASAP7_75t_L g1734 ( 
.A(n_1724),
.B(n_1712),
.C(n_1689),
.D(n_1668),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_SL g1735 ( 
.A(n_1717),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_SL g1736 ( 
.A1(n_1725),
.A2(n_1607),
.B(n_1629),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1733),
.B(n_1661),
.C(n_1657),
.D(n_1656),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1734),
.B(n_1656),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1731),
.A2(n_1661),
.B(n_1657),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1736),
.A2(n_1624),
.B(n_1612),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1728),
.A2(n_1543),
.B1(n_1604),
.B2(n_1603),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1741),
.A2(n_1729),
.B1(n_1730),
.B2(n_1727),
.C(n_1732),
.Y(n_1742)
);

OAI321xp33_ASAP7_75t_L g1743 ( 
.A1(n_1737),
.A2(n_1735),
.A3(n_1621),
.B1(n_1623),
.B2(n_1599),
.C(n_1605),
.Y(n_1743)
);

NAND2x1_ASAP7_75t_SL g1744 ( 
.A(n_1738),
.B(n_1607),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1739),
.A2(n_1627),
.B(n_1624),
.Y(n_1745)
);

NAND4xp25_ASAP7_75t_L g1746 ( 
.A(n_1740),
.B(n_1607),
.C(n_1605),
.D(n_1601),
.Y(n_1746)
);

OAI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1618),
.B(n_1605),
.C(n_1631),
.Y(n_1747)
);

NOR3xp33_ASAP7_75t_L g1748 ( 
.A(n_1742),
.B(n_1618),
.C(n_1548),
.Y(n_1748)
);

NAND4xp75_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1631),
.C(n_1604),
.D(n_1603),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1747),
.A2(n_1601),
.B1(n_1629),
.B2(n_1604),
.Y(n_1750)
);

AO22x1_ASAP7_75t_L g1751 ( 
.A1(n_1744),
.A2(n_1607),
.B1(n_1629),
.B2(n_1618),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1743),
.A2(n_1607),
.B(n_1629),
.Y(n_1752)
);

AOI222xp33_ASAP7_75t_L g1753 ( 
.A1(n_1751),
.A2(n_1543),
.B1(n_1746),
.B2(n_1530),
.C1(n_1511),
.C2(n_1528),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1752),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1750),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1754),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1756),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1757),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1757),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_1758),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1759),
.B(n_1755),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1760),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_L g1763 ( 
.A(n_1761),
.B(n_1748),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1762),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1764),
.B(n_1763),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1753),
.B1(n_1749),
.B2(n_1619),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_R g1767 ( 
.A1(n_1766),
.A2(n_1601),
.B1(n_1625),
.B2(n_1622),
.C(n_1580),
.Y(n_1767)
);

AOI211xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1449),
.B(n_1462),
.C(n_1617),
.Y(n_1768)
);


endmodule