module fake_jpeg_31265_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_55),
.Y(n_139)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_26),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_72),
.Y(n_103)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_82),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_28),
.Y(n_121)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_24),
.B(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_14),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_41),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_21),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_38),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_104),
.B(n_106),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_28),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_111),
.B(n_50),
.Y(n_226)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_101),
.Y(n_115)
);

CKINVDCx9p33_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_43),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_121),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_40),
.C(n_43),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_154),
.Y(n_172)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_123),
.B(n_124),
.Y(n_187)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_55),
.B(n_40),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g212 ( 
.A(n_131),
.B(n_118),
.C(n_148),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_71),
.B1(n_78),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_135),
.A2(n_153),
.B1(n_131),
.B2(n_98),
.Y(n_224)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_66),
.B(n_36),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_150),
.B(n_165),
.Y(n_219)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_54),
.A2(n_38),
.B1(n_23),
.B2(n_36),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_74),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_61),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_61),
.B(n_19),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_166),
.Y(n_262)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_167),
.Y(n_267)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_103),
.B(n_87),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_178),
.C(n_211),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_62),
.B1(n_64),
.B2(n_58),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_195),
.B1(n_153),
.B2(n_129),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_103),
.B(n_92),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_186),
.Y(n_231)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_95),
.B1(n_53),
.B2(n_38),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_205),
.B1(n_215),
.B2(n_135),
.Y(n_236)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_193),
.B(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_113),
.A2(n_68),
.B1(n_67),
.B2(n_89),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_91),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_196),
.B(n_218),
.Y(n_273)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

BUFx16f_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_204),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_119),
.A2(n_23),
.B1(n_38),
.B2(n_69),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_207),
.Y(n_247)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_213),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_117),
.B(n_88),
.C(n_90),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_209),
.B(n_3),
.C(n_5),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_111),
.A2(n_65),
.B1(n_39),
.B2(n_14),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_134),
.B(n_12),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_144),
.A2(n_23),
.B1(n_69),
.B2(n_50),
.Y(n_215)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_221),
.B(n_226),
.Y(n_248)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_217),
.B(n_223),
.Y(n_253)
);

CKINVDCx12_ASAP7_75t_R g218 ( 
.A(n_138),
.Y(n_218)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_220),
.A2(n_222),
.B1(n_2),
.B2(n_3),
.Y(n_270)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_136),
.B(n_39),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_215),
.B1(n_188),
.B2(n_205),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_161),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_235),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_136),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_234),
.B(n_245),
.C(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_110),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_236),
.B(n_240),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_122),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_244),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_177),
.A2(n_163),
.B1(n_128),
.B2(n_120),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_241),
.A2(n_256),
.B1(n_263),
.B2(n_274),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_172),
.A2(n_165),
.B1(n_156),
.B2(n_77),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_243),
.A2(n_261),
.B1(n_271),
.B2(n_242),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_138),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_175),
.B(n_1),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_187),
.B(n_139),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_258),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_168),
.B(n_139),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_195),
.A2(n_52),
.B1(n_60),
.B2(n_14),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_184),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_183),
.B(n_1),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_5),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_222),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_167),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_7),
.Y(n_320)
);

INVx4_ASAP7_75t_SL g279 ( 
.A(n_252),
.Y(n_279)
);

INVx11_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

CKINVDCx12_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_190),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_295),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_166),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_284),
.B(n_288),
.Y(n_355)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_286),
.A2(n_293),
.B1(n_294),
.B2(n_308),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_233),
.B(n_198),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_206),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_250),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_291),
.B(n_292),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_216),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_256),
.A2(n_225),
.B1(n_185),
.B2(n_199),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_201),
.B1(n_213),
.B2(n_203),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_228),
.B(n_216),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_242),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_300),
.Y(n_339)
);

FAx1_ASAP7_75t_L g297 ( 
.A(n_238),
.B(n_180),
.CI(n_204),
.CON(n_297),
.SN(n_297)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_297),
.A2(n_251),
.B(n_252),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_232),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_207),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_303),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_221),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_244),
.A2(n_220),
.B(n_6),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_237),
.B(n_320),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_238),
.B(n_234),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_305),
.B(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_316),
.Y(n_347)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_227),
.Y(n_307)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_254),
.A2(n_170),
.B1(n_173),
.B2(n_181),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_6),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_240),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_324),
.B1(n_263),
.B2(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_278),
.B(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_315),
.B(n_262),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_7),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_260),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_317),
.Y(n_326)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_318),
.Y(n_361)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_319),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_322),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_245),
.B(n_8),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_277),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_248),
.B(n_232),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_257),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_323),
.B(n_325),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_247),
.B(n_246),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_330),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_301),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_326),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_281),
.A2(n_238),
.A3(n_241),
.B1(n_245),
.B2(n_270),
.Y(n_336)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_265),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_282),
.B(n_246),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_298),
.A2(n_314),
.B1(n_311),
.B2(n_289),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_342),
.A2(n_346),
.B1(n_341),
.B2(n_353),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_299),
.A2(n_262),
.B(n_251),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_343),
.A2(n_359),
.B(n_296),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_322),
.B(n_297),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_298),
.A2(n_255),
.B1(n_269),
.B2(n_272),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_283),
.A2(n_255),
.B(n_269),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_348),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_349),
.B(n_354),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_272),
.B1(n_275),
.B2(n_277),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_358),
.B1(n_360),
.B2(n_308),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_282),
.B(n_275),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_290),
.A2(n_229),
.B1(n_237),
.B2(n_286),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_290),
.A2(n_293),
.B1(n_287),
.B2(n_310),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_289),
.B(n_316),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_365),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_287),
.B(n_305),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_361),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_370),
.B(n_396),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_344),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_371),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_372),
.A2(n_378),
.B1(n_381),
.B2(n_384),
.Y(n_421)
);

CKINVDCx12_ASAP7_75t_R g373 ( 
.A(n_327),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_375),
.B(n_342),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_344),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_379),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_339),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_330),
.A2(n_297),
.B1(n_304),
.B2(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_383),
.A2(n_386),
.B(n_387),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_360),
.A2(n_312),
.B1(n_306),
.B2(n_294),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_329),
.A2(n_313),
.B1(n_285),
.B2(n_307),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_388),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_315),
.B(n_279),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_329),
.A2(n_279),
.B1(n_319),
.B2(n_358),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_331),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_393),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_328),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_395),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_392),
.B(n_327),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_341),
.A2(n_353),
.B1(n_352),
.B2(n_364),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_326),
.B(n_335),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_399),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_362),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_398),
.B(n_400),
.Y(n_413)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_355),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_359),
.A2(n_348),
.B1(n_338),
.B2(n_336),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_367),
.A2(n_348),
.B1(n_366),
.B2(n_345),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_403),
.A2(n_405),
.B1(n_407),
.B2(n_415),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_334),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_414),
.C(n_377),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_367),
.A2(n_348),
.B1(n_363),
.B2(n_343),
.Y(n_407)
);

A2O1A1O1Ixp25_ASAP7_75t_L g409 ( 
.A1(n_389),
.A2(n_333),
.B(n_347),
.C(n_349),
.D(n_337),
.Y(n_409)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_369),
.B(n_333),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_371),
.B(n_347),
.Y(n_415)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_415),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_417),
.A2(n_431),
.B1(n_411),
.B2(n_405),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_376),
.B(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_383),
.A2(n_332),
.B(n_350),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_419),
.A2(n_390),
.B(n_374),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_356),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_427),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_423),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_356),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_380),
.B(n_350),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_431),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_351),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_389),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_441),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_403),
.A2(n_401),
.B1(n_378),
.B2(n_407),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_433),
.A2(n_457),
.B1(n_411),
.B2(n_410),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_434),
.B(n_406),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_377),
.C(n_387),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_438),
.C(n_440),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_386),
.B(n_368),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_453),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_375),
.C(n_391),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_379),
.C(n_384),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_394),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_395),
.Y(n_442)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_421),
.A2(n_400),
.B1(n_398),
.B2(n_368),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_425),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_388),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_448),
.C(n_454),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_382),
.C(n_385),
.Y(n_448)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_450),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_416),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_451),
.B(n_452),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_351),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_427),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_390),
.C(n_420),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_445),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_459),
.B(n_460),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_436),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_439),
.B(n_413),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_465),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_456),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_469),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_409),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_428),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_408),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_477),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_456),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_474),
.B(n_476),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_446),
.A2(n_430),
.B1(n_423),
.B2(n_429),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_433),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g481 ( 
.A(n_464),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_491),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_495),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_458),
.A2(n_437),
.B(n_410),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_466),
.B(n_458),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_484),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_477),
.A2(n_438),
.B1(n_454),
.B2(n_457),
.Y(n_487)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_440),
.C(n_441),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_490),
.B(n_494),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_475),
.B(n_412),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_447),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_460),
.B(n_455),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_497),
.A2(n_501),
.B(n_489),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_480),
.A2(n_465),
.B1(n_448),
.B2(n_467),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_499),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_419),
.B(n_475),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_471),
.C(n_459),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_506),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_472),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_472),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_493),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_429),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_423),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_506),
.B(n_484),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_510),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_513),
.C(n_516),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_504),
.A2(n_483),
.B(n_488),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_512),
.A2(n_517),
.B(n_497),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_479),
.C(n_482),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_470),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_502),
.Y(n_518)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_498),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_520),
.C(n_499),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_473),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_521),
.A2(n_501),
.B(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_525),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_522),
.C(n_523),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_524),
.A3(n_508),
.B1(n_485),
.B2(n_505),
.C1(n_424),
.C2(n_412),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_507),
.B(n_450),
.C(n_527),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_496),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_531),
.B(n_496),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_430),
.C(n_424),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_478),
.Y(n_534)
);


endmodule