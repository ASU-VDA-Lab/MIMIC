module fake_jpeg_13392_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_1),
.A2(n_3),
.B(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_24),
.B(n_17),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_6),
.Y(n_23)
);

OR2x4_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_9),
.B(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_12),
.B1(n_17),
.B2(n_13),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_29),
.B(n_34),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_4),
.B1(n_13),
.B2(n_37),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_35),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_36),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_28),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_28),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_42),
.C(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_41),
.Y(n_53)
);

OA21x2_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_39),
.B(n_49),
.Y(n_52)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_41),
.C(n_47),
.D(n_48),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_39),
.B(n_52),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_44),
.Y(n_56)
);


endmodule