module fake_jpeg_30435_n_379 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_379);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_60),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_14),
.Y(n_97)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_18),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_17),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_1),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_65),
.Y(n_96)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_42),
.B1(n_38),
.B2(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_22),
.B1(n_47),
.B2(n_32),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_42),
.B1(n_38),
.B2(n_33),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_83),
.B1(n_85),
.B2(n_29),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_42),
.B1(n_38),
.B2(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_78),
.B1(n_28),
.B2(n_37),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_25),
.B1(n_35),
.B2(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_29),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_34),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_25),
.C(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_21),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_113),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_110),
.B1(n_116),
.B2(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_108),
.A2(n_132),
.B1(n_62),
.B2(n_37),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_33),
.B(n_22),
.C(n_32),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_118),
.B(n_75),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_63),
.B1(n_66),
.B2(n_64),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_127),
.Y(n_147)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_32),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_124),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_56),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_86),
.C(n_77),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_52),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_59),
.B1(n_35),
.B2(n_24),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_24),
.B(n_37),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_52),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_130),
.Y(n_161)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_133),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_95),
.B1(n_94),
.B2(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_66),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_35),
.B1(n_45),
.B2(n_28),
.Y(n_132)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_71),
.B1(n_85),
.B2(n_92),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_137),
.B(n_100),
.Y(n_189)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_93),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_92),
.B1(n_79),
.B2(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_117),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_96),
.B1(n_91),
.B2(n_79),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_157),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_96),
.B1(n_91),
.B2(n_79),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_89),
.B(n_96),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_158),
.B(n_110),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_156),
.C(n_123),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_112),
.B(n_120),
.C(n_122),
.Y(n_154)
);

INVx5_ASAP7_75t_SL g170 ( 
.A(n_154),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_81),
.C(n_77),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_81),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_64),
.B1(n_62),
.B2(n_99),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_162),
.B1(n_107),
.B2(n_103),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_100),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_102),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_189),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_116),
.B1(n_118),
.B2(n_123),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_185),
.B1(n_192),
.B2(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_177),
.B(n_153),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_187),
.B1(n_160),
.B2(n_151),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_183),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_109),
.B1(n_119),
.B2(n_107),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_190),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_101),
.B1(n_114),
.B2(n_117),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_128),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_152),
.C(n_158),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_137),
.A2(n_131),
.B(n_103),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_212),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_156),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_211),
.C(n_188),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_200),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_204),
.B1(n_207),
.B2(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_162),
.B1(n_163),
.B2(n_145),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_210),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_135),
.B1(n_138),
.B2(n_154),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_205),
.A2(n_207),
.B1(n_206),
.B2(n_195),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_160),
.B1(n_165),
.B2(n_152),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_187),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_135),
.B1(n_151),
.B2(n_158),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_161),
.C(n_159),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_171),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_161),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_219),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_190),
.B(n_176),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_220),
.A2(n_236),
.B(n_131),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_229),
.C(n_230),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_180),
.B(n_183),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_234),
.B(n_245),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_205),
.B1(n_202),
.B2(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_231),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_188),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_173),
.C(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_168),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_232),
.B(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_159),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_208),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_184),
.B(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_173),
.C(n_174),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_239),
.C(n_143),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_209),
.B(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_218),
.B1(n_146),
.B2(n_182),
.Y(n_267)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_248),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_209),
.A2(n_170),
.B(n_135),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_198),
.A2(n_170),
.B(n_135),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_204),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_203),
.A2(n_164),
.B(n_172),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_201),
.B(n_172),
.Y(n_253)
);

INVxp33_ASAP7_75t_SL g248 ( 
.A(n_206),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_266),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_252),
.A2(n_256),
.B1(n_264),
.B2(n_242),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_212),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_260),
.B(n_275),
.Y(n_281)
);

XOR2x2_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_138),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_37),
.Y(n_298)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_245),
.B1(n_236),
.B2(n_234),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_141),
.C(n_201),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_265),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_218),
.B1(n_216),
.B2(n_138),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_267),
.B1(n_270),
.B2(n_227),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_218),
.B1(n_182),
.B2(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_155),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_221),
.A2(n_139),
.B1(n_138),
.B2(n_155),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_147),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_138),
.C(n_146),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_191),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_273),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_221),
.A2(n_136),
.B1(n_191),
.B2(n_149),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_133),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_233),
.B(n_143),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_239),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_282),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_235),
.C(n_230),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_285),
.C(n_287),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_280),
.A2(n_294),
.B1(n_264),
.B2(n_271),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_225),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_221),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_247),
.C(n_244),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_269),
.B1(n_263),
.B2(n_11),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_238),
.C(n_231),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_228),
.C(n_226),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_292),
.C(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_226),
.C(n_136),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_251),
.B(n_12),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_293),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_127),
.B1(n_115),
.B2(n_51),
.Y(n_294)
);

NAND4xp25_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_133),
.C(n_11),
.D(n_12),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_275),
.B(n_274),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_305),
.B(n_308),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_267),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_251),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_303),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_256),
.B(n_274),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_253),
.B(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_252),
.C(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_287),
.C(n_280),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_313),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_271),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_285),
.B(n_263),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_294),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_321),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_295),
.C(n_283),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_327),
.C(n_330),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_278),
.Y(n_321)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_283),
.C(n_290),
.Y(n_327)
);

AOI221xp5_ASAP7_75t_L g329 ( 
.A1(n_305),
.A2(n_269),
.B1(n_284),
.B2(n_277),
.C(n_292),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_304),
.B(n_315),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_298),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_17),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_331),
.B(n_333),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_15),
.B(n_14),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_28),
.B(n_3),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_299),
.B(n_312),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_334),
.B(n_335),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_325),
.A2(n_307),
.B(n_306),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_4),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_323),
.A2(n_313),
.B1(n_304),
.B2(n_317),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_343),
.B1(n_333),
.B2(n_326),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_310),
.C(n_37),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_330),
.C(n_320),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_28),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_347),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_1),
.B(n_2),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_1),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_345),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_328),
.A2(n_2),
.B(n_3),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_350),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_324),
.C(n_327),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_354),
.Y(n_363)
);

AOI322xp5_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_321),
.A3(n_28),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_3),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_352),
.A2(n_356),
.B(n_348),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_340),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_357),
.Y(n_365)
);

AO221x1_ASAP7_75t_L g356 ( 
.A1(n_339),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_28),
.C(n_20),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_353),
.A2(n_336),
.B(n_341),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_360),
.B(n_362),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_350),
.A2(n_347),
.B(n_345),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_364),
.A2(n_366),
.B(n_4),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_358),
.B(n_5),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_358),
.C(n_20),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_367),
.A2(n_370),
.B(n_371),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_20),
.C(n_6),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_372),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_7),
.B(n_8),
.Y(n_375)
);

AOI322xp5_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_20),
.C1(n_241),
.C2(n_307),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_369),
.B1(n_9),
.B2(n_10),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_SL g378 ( 
.A1(n_376),
.A2(n_377),
.B(n_9),
.C(n_10),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_378),
.B(n_374),
.Y(n_379)
);


endmodule