module fake_aes_9657_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
OR2x6_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
AO31x2_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_4), .A3(n_1), .B(n_2), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_2), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_5), .B(n_0), .Y(n_8) );
NAND3xp33_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .C(n_0), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
XNOR2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_7), .Y(n_11) );
OAI22x1_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_10), .B1(n_8), .B2(n_1), .Y(n_12) );
AOI22xp33_ASAP7_75t_SL g13 ( .A1(n_12), .A2(n_11), .B1(n_0), .B2(n_1), .Y(n_13) );
endmodule