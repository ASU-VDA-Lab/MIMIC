module fake_jpeg_7534_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx8_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_11),
.B2(n_19),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_11),
.B1(n_16),
.B2(n_13),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_38),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_19),
.B1(n_17),
.B2(n_10),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_21),
.B1(n_11),
.B2(n_20),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_19),
.C(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_23),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_23),
.B1(n_15),
.B2(n_12),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_52),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_23),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_35),
.C(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_57),
.B(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_37),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_43),
.C(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_42),
.Y(n_65)
);

A2O1A1O1Ixp25_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_69),
.B(n_49),
.C(n_15),
.D(n_12),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_59),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_24),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_58),
.B(n_57),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_32),
.B(n_30),
.Y(n_84)
);

AOI221xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_78),
.B1(n_70),
.B2(n_75),
.C(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_59),
.B1(n_31),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_31),
.B1(n_60),
.B2(n_69),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_30),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_86),
.B1(n_1),
.B2(n_3),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_81),
.B1(n_85),
.B2(n_83),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_32),
.C(n_30),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_15),
.B(n_12),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_76),
.B1(n_78),
.B2(n_15),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_4),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_5),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_79),
.B(n_4),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_97),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_3),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_87),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI21x1_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_6),
.B(n_7),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_101),
.B(n_7),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_8),
.C(n_103),
.Y(n_106)
);


endmodule