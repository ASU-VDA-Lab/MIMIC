module real_aes_1361_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_0), .B(n_136), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_1), .A2(n_118), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_2), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_3), .B(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g123 ( .A(n_4), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_5), .B(n_126), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_6), .B(n_113), .Y(n_463) );
INVx1_ASAP7_75t_L g491 ( .A(n_7), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g810 ( .A(n_8), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_9), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_10), .A2(n_105), .B1(n_774), .B2(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_10), .Y(n_801) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_11), .B(n_130), .Y(n_163) );
INVx2_ASAP7_75t_L g115 ( .A(n_12), .Y(n_115) );
AOI221x1_ASAP7_75t_L g205 ( .A1(n_13), .A2(n_25), .B1(n_118), .B2(n_136), .C(n_206), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_14), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_15), .B(n_136), .Y(n_159) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_16), .A2(n_157), .B(n_158), .Y(n_156) );
INVx1_ASAP7_75t_L g472 ( .A(n_17), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_18), .B(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_19), .B(n_126), .Y(n_125) );
AO21x1_ASAP7_75t_L g177 ( .A1(n_20), .A2(n_136), .B(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g429 ( .A(n_21), .Y(n_429) );
INVx1_ASAP7_75t_L g470 ( .A(n_22), .Y(n_470) );
INVx1_ASAP7_75t_SL g456 ( .A(n_23), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_24), .B(n_137), .Y(n_550) );
NAND2x1_ASAP7_75t_L g191 ( .A(n_26), .B(n_126), .Y(n_191) );
AOI33xp33_ASAP7_75t_L g518 ( .A1(n_27), .A2(n_53), .A3(n_446), .B1(n_453), .B2(n_519), .B3(n_520), .Y(n_518) );
NAND2x1_ASAP7_75t_L g145 ( .A(n_28), .B(n_130), .Y(n_145) );
INVx1_ASAP7_75t_L g500 ( .A(n_29), .Y(n_500) );
OR2x2_ASAP7_75t_L g114 ( .A(n_30), .B(n_85), .Y(n_114) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_30), .A2(n_85), .B(n_115), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_31), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_32), .B(n_130), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_33), .B(n_126), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_34), .B(n_130), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_35), .A2(n_118), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g119 ( .A(n_36), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g134 ( .A(n_36), .B(n_123), .Y(n_134) );
INVx1_ASAP7_75t_L g452 ( .A(n_36), .Y(n_452) );
OR2x6_ASAP7_75t_L g427 ( .A(n_37), .B(n_428), .Y(n_427) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_37), .B(n_809), .C(n_811), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_38), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_39), .B(n_136), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_40), .B(n_444), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_41), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_42), .A2(n_113), .B1(n_153), .B2(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_43), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_44), .B(n_137), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_45), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_46), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_47), .B(n_130), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_48), .B(n_157), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_49), .B(n_137), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_50), .A2(n_118), .B(n_144), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_51), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_52), .B(n_130), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_54), .B(n_137), .Y(n_530) );
INVx1_ASAP7_75t_L g122 ( .A(n_55), .Y(n_122) );
INVx1_ASAP7_75t_L g132 ( .A(n_55), .Y(n_132) );
AND2x2_ASAP7_75t_L g531 ( .A(n_56), .B(n_149), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_57), .A2(n_73), .B1(n_444), .B2(n_450), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_58), .B(n_444), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_59), .B(n_126), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_60), .B(n_153), .Y(n_508) );
AOI21xp5_ASAP7_75t_SL g480 ( .A1(n_61), .A2(n_450), .B(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_62), .A2(n_118), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g466 ( .A(n_63), .Y(n_466) );
AO21x1_ASAP7_75t_L g179 ( .A1(n_64), .A2(n_118), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_65), .B(n_136), .Y(n_167) );
INVx1_ASAP7_75t_L g529 ( .A(n_66), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_67), .B(n_136), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_68), .A2(n_450), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g228 ( .A(n_69), .B(n_150), .Y(n_228) );
INVx1_ASAP7_75t_L g120 ( .A(n_70), .Y(n_120) );
INVx1_ASAP7_75t_L g128 ( .A(n_70), .Y(n_128) );
AND2x2_ASAP7_75t_L g151 ( .A(n_71), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_72), .B(n_444), .Y(n_521) );
AND2x2_ASAP7_75t_L g459 ( .A(n_74), .B(n_152), .Y(n_459) );
INVx1_ASAP7_75t_L g467 ( .A(n_75), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_76), .A2(n_450), .B(n_455), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_77), .A2(n_450), .B(n_513), .C(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_SL g772 ( .A1(n_78), .A2(n_102), .B1(n_773), .B2(n_777), .Y(n_772) );
INVx1_ASAP7_75t_L g430 ( .A(n_79), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_79), .B(n_429), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_80), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g165 ( .A(n_81), .B(n_152), .Y(n_165) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_82), .B(n_152), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_83), .A2(n_450), .B1(n_516), .B2(n_517), .Y(n_515) );
AND2x2_ASAP7_75t_L g178 ( .A(n_84), .B(n_113), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_86), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g195 ( .A(n_87), .B(n_152), .Y(n_195) );
INVx1_ASAP7_75t_L g482 ( .A(n_88), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_89), .B(n_126), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_90), .A2(n_118), .B(n_124), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_91), .B(n_130), .Y(n_207) );
AND2x2_ASAP7_75t_L g522 ( .A(n_92), .B(n_152), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_93), .B(n_126), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_94), .A2(n_498), .B(n_499), .C(n_501), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_95), .Y(n_102) );
BUFx2_ASAP7_75t_L g785 ( .A(n_96), .Y(n_785) );
BUFx2_ASAP7_75t_SL g798 ( .A(n_96), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_97), .A2(n_118), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_98), .B(n_137), .Y(n_483) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_804), .B(n_813), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_781), .B(n_794), .Y(n_100) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_103), .B(n_772), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_422), .B1(n_431), .B2(n_435), .Y(n_104) );
INVx2_ASAP7_75t_L g774 ( .A(n_105), .Y(n_774) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_320), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_232), .C(n_287), .Y(n_106) );
AOI221xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_172), .B1(n_196), .B2(n_200), .C(n_210), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_155), .Y(n_108) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_109), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g231 ( .A(n_109), .Y(n_231) );
AND2x2_ASAP7_75t_L g276 ( .A(n_109), .B(n_213), .Y(n_276) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_140), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g264 ( .A(n_111), .Y(n_264) );
INVx1_ASAP7_75t_L g274 ( .A(n_111), .Y(n_274) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_138), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_112), .B(n_139), .Y(n_138) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_112), .A2(n_116), .B(n_138), .Y(n_238) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_113), .A2(n_159), .B(n_160), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_113), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_113), .B(n_133), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_113), .A2(n_480), .B(n_484), .Y(n_479) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_114), .B(n_115), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_135), .Y(n_116) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx3_ASAP7_75t_L g448 ( .A(n_119), .Y(n_448) );
AND2x6_ASAP7_75t_L g130 ( .A(n_120), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g454 ( .A(n_120), .Y(n_454) );
AND2x4_ASAP7_75t_L g450 ( .A(n_121), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x4_ASAP7_75t_L g126 ( .A(n_122), .B(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g446 ( .A(n_122), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_123), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_133), .Y(n_124) );
INVxp67_ASAP7_75t_L g473 ( .A(n_126), .Y(n_473) );
AND2x4_ASAP7_75t_L g137 ( .A(n_127), .B(n_131), .Y(n_137) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVxp67_ASAP7_75t_L g471 ( .A(n_130), .Y(n_471) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_133), .A2(n_145), .B(n_146), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_133), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_133), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_133), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_133), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_133), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_133), .A2(n_225), .B(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g455 ( .A1(n_133), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_133), .A2(n_457), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_133), .A2(n_457), .B(n_491), .C(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g516 ( .A(n_133), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_133), .A2(n_457), .B(n_529), .C(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_133), .A2(n_550), .B(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g136 ( .A(n_134), .B(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_134), .Y(n_501) );
INVx1_ASAP7_75t_L g468 ( .A(n_137), .Y(n_468) );
OR2x2_ASAP7_75t_L g253 ( .A(n_140), .B(n_156), .Y(n_253) );
NAND2x1p5_ASAP7_75t_L g284 ( .A(n_140), .B(n_199), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_140), .B(n_164), .Y(n_297) );
INVx2_ASAP7_75t_L g306 ( .A(n_140), .Y(n_306) );
AND2x2_ASAP7_75t_L g327 ( .A(n_140), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g411 ( .A(n_140), .B(n_230), .Y(n_411) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g239 ( .A(n_141), .B(n_164), .Y(n_239) );
AND2x2_ASAP7_75t_L g372 ( .A(n_141), .B(n_199), .Y(n_372) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_141), .Y(n_398) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B(n_151), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_148), .A2(n_442), .B(n_459), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_149), .A2(n_167), .B(n_168), .Y(n_166) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_149), .A2(n_205), .B(n_209), .Y(n_204) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_149), .A2(n_205), .B(n_209), .Y(n_216) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_152), .A2(n_194), .B1(n_497), .B2(n_502), .Y(n_496) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_153), .B(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx4f_ASAP7_75t_L g157 ( .A(n_154), .Y(n_157) );
AND2x4_ASAP7_75t_L g326 ( .A(n_155), .B(n_327), .Y(n_326) );
AOI321xp33_ASAP7_75t_L g340 ( .A1(n_155), .A2(n_269), .A3(n_270), .B1(n_302), .B2(n_341), .C(n_344), .Y(n_340) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_164), .Y(n_155) );
BUFx3_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
INVx2_ASAP7_75t_L g230 ( .A(n_156), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_156), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g263 ( .A(n_156), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g296 ( .A(n_156), .Y(n_296) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_157), .A2(n_489), .B(n_493), .Y(n_488) );
INVx2_ASAP7_75t_SL g513 ( .A(n_157), .Y(n_513) );
INVx5_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
NOR2x1_ASAP7_75t_SL g248 ( .A(n_164), .B(n_238), .Y(n_248) );
BUFx2_ASAP7_75t_L g343 ( .A(n_164), .Y(n_343) );
OR2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVxp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_185), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_174), .B(n_242), .Y(n_241) );
NOR4xp25_ASAP7_75t_L g344 ( .A(n_174), .B(n_338), .C(n_342), .D(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g382 ( .A(n_174), .Y(n_382) );
AND2x2_ASAP7_75t_L g416 ( .A(n_174), .B(n_356), .Y(n_416) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g271 ( .A(n_176), .Y(n_271) );
OAI21x1_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_179), .B(n_183), .Y(n_176) );
INVx1_ASAP7_75t_L g184 ( .A(n_178), .Y(n_184) );
AOI33xp33_ASAP7_75t_L g412 ( .A1(n_185), .A2(n_214), .A3(n_245), .B1(n_261), .B2(n_367), .B3(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g202 ( .A(n_186), .B(n_203), .Y(n_202) );
AND2x4_ASAP7_75t_L g212 ( .A(n_186), .B(n_213), .Y(n_212) );
BUFx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g219 ( .A(n_187), .Y(n_219) );
INVxp67_ASAP7_75t_L g300 ( .A(n_187), .Y(n_300) );
AND2x2_ASAP7_75t_L g356 ( .A(n_187), .B(n_221), .Y(n_356) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_194), .B(n_195), .Y(n_187) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_188), .A2(n_194), .B(n_195), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_193), .Y(n_188) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_194), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_194), .A2(n_222), .B(n_228), .Y(n_257) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_194), .A2(n_525), .B(n_531), .Y(n_524) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_194), .A2(n_525), .B(n_531), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_196), .A2(n_378), .B(n_379), .Y(n_377) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
AND2x2_ASAP7_75t_L g365 ( .A(n_197), .B(n_239), .Y(n_365) );
AND3x2_ASAP7_75t_L g367 ( .A(n_197), .B(n_251), .C(n_306), .Y(n_367) );
INVx3_ASAP7_75t_SL g319 ( .A(n_198), .Y(n_319) );
INVx4_ASAP7_75t_L g213 ( .A(n_199), .Y(n_213) );
AND2x2_ASAP7_75t_L g251 ( .A(n_199), .B(n_238), .Y(n_251) );
INVxp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g245 ( .A(n_203), .Y(n_245) );
AND2x4_ASAP7_75t_L g270 ( .A(n_203), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g333 ( .A(n_203), .B(n_221), .Y(n_333) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g303 ( .A(n_204), .Y(n_303) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_204), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_R g210 ( .A1(n_211), .A2(n_214), .B(n_218), .C(n_229), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g262 ( .A(n_213), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_213), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_213), .B(n_230), .Y(n_391) );
INVx1_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g373 ( .A(n_215), .B(n_363), .Y(n_373) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g220 ( .A(n_216), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g242 ( .A(n_216), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g258 ( .A(n_216), .B(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g291 ( .A(n_216), .B(n_271), .Y(n_291) );
AND2x4_ASAP7_75t_L g256 ( .A(n_217), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g280 ( .A(n_217), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g318 ( .A(n_217), .B(n_243), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g246 ( .A(n_219), .B(n_243), .Y(n_246) );
AND2x2_ASAP7_75t_L g261 ( .A(n_219), .B(n_221), .Y(n_261) );
BUFx2_ASAP7_75t_L g317 ( .A(n_219), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_219), .B(n_242), .Y(n_331) );
INVx2_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_227), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g279 ( .A1(n_229), .A2(n_280), .B1(n_282), .B2(n_286), .Y(n_279) );
INVx2_ASAP7_75t_SL g310 ( .A(n_229), .Y(n_310) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x2_ASAP7_75t_L g285 ( .A(n_230), .B(n_238), .Y(n_285) );
INVx1_ASAP7_75t_L g392 ( .A(n_231), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_265), .C(n_279), .Y(n_232) );
OAI221xp5_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_240), .B1(n_244), .B2(n_247), .C(n_249), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_239), .Y(n_235) );
INVxp67_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g293 ( .A(n_237), .Y(n_293) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_237), .Y(n_421) );
INVx1_ASAP7_75t_L g384 ( .A(n_239), .Y(n_384) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_239), .B(n_263), .Y(n_394) );
INVxp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_243), .B(n_271), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
OR2x2_ASAP7_75t_L g277 ( .A(n_245), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g355 ( .A(n_245), .Y(n_355) );
AND2x2_ASAP7_75t_L g290 ( .A(n_246), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g336 ( .A(n_248), .B(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g413 ( .A(n_248), .B(n_411), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B1(n_261), .B2(n_262), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g272 ( .A(n_253), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx2_ASAP7_75t_L g278 ( .A(n_256), .Y(n_278) );
AND2x4_ASAP7_75t_L g302 ( .A(n_256), .B(n_303), .Y(n_302) );
OAI21xp33_ASAP7_75t_SL g332 ( .A1(n_256), .A2(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g359 ( .A(n_256), .B(n_317), .Y(n_359) );
INVx2_ASAP7_75t_L g281 ( .A(n_257), .Y(n_281) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_257), .Y(n_314) );
INVx1_ASAP7_75t_SL g338 ( .A(n_258), .Y(n_338) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g269 ( .A(n_260), .Y(n_269) );
AND2x4_ASAP7_75t_SL g363 ( .A(n_260), .B(n_281), .Y(n_363) );
AND2x2_ASAP7_75t_L g360 ( .A(n_263), .B(n_306), .Y(n_360) );
AND2x2_ASAP7_75t_L g386 ( .A(n_263), .B(n_372), .Y(n_386) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
INVx1_ASAP7_75t_L g328 ( .A(n_264), .Y(n_328) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_272), .B1(n_275), .B2(n_277), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_270), .B(n_281), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_270), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g409 ( .A(n_270), .Y(n_409) );
INVx2_ASAP7_75t_SL g334 ( .A(n_272), .Y(n_334) );
AND2x2_ASAP7_75t_L g346 ( .A(n_274), .B(n_306), .Y(n_346) );
INVx2_ASAP7_75t_L g352 ( .A(n_274), .Y(n_352) );
INVxp33_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_280), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g402 ( .A(n_280), .Y(n_402) );
INVx1_ASAP7_75t_L g330 ( .A(n_282), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_283), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g341 ( .A(n_285), .B(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_285), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_414) );
NOR3xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_309), .C(n_312), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .B1(n_294), .B2(n_298), .C(n_301), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_SL g407 ( .A(n_292), .Y(n_407) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g376 ( .A(n_293), .B(n_342), .Y(n_376) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g307 ( .A(n_296), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g378 ( .A(n_298), .Y(n_378) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g375 ( .A(n_299), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_300), .Y(n_381) );
OR2x2_ASAP7_75t_L g404 ( .A(n_300), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g313 ( .A(n_303), .Y(n_313) );
AND2x2_ASAP7_75t_L g383 ( .A(n_303), .B(n_363), .Y(n_383) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_303), .B(n_316), .Y(n_415) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g420 ( .A(n_306), .Y(n_420) );
INVx1_ASAP7_75t_L g370 ( .A(n_308), .Y(n_370) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_315), .C(n_319), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_313), .B(n_363), .Y(n_387) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_316), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g324 ( .A(n_318), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g405 ( .A(n_318), .Y(n_405) );
NAND4xp75_ASAP7_75t_L g320 ( .A(n_321), .B(n_377), .C(n_393), .D(n_414), .Y(n_320) );
NOR3x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_339), .C(n_361), .Y(n_321) );
NAND4xp75_ASAP7_75t_L g322 ( .A(n_323), .B(n_329), .C(n_332), .D(n_335), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_324), .B(n_326), .Y(n_323) );
AND2x2_ASAP7_75t_L g374 ( .A(n_325), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g399 ( .A(n_326), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_SL g388 ( .A(n_331), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_347), .Y(n_339) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_343), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_353), .B(n_357), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI322xp33_ASAP7_75t_L g379 ( .A1(n_351), .A2(n_380), .A3(n_384), .B1(n_385), .B2(n_387), .C1(n_388), .C2(n_389), .Y(n_379) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_352), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_355), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_356), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
OAI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B(n_366), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_373), .B1(n_374), .B2(n_376), .Y(n_368) );
NOR2xp33_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .Y(n_380) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_386), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g396 ( .A(n_391), .B(n_397), .Y(n_396) );
O2A1O1Ixp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_400), .C(n_403), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_406), .B1(n_408), .B2(n_410), .C(n_412), .Y(n_403) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
CKINVDCx6p67_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
INVx4_ASAP7_75t_SL g775 ( .A(n_423), .Y(n_775) );
INVx3_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
AND2x6_ASAP7_75t_SL g425 ( .A(n_426), .B(n_427), .Y(n_425) );
OR2x6_ASAP7_75t_SL g433 ( .A(n_426), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g780 ( .A(n_426), .B(n_427), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_426), .B(n_434), .Y(n_792) );
CKINVDCx16_ASAP7_75t_R g811 ( .A(n_426), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_427), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
OAI22x1_ASAP7_75t_L g773 ( .A1(n_433), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_435), .Y(n_776) );
OR3x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_637), .C(n_708), .Y(n_435) );
NAND3x1_ASAP7_75t_SL g436 ( .A(n_437), .B(n_564), .C(n_586), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_554), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_485), .B1(n_532), .B2(n_536), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_439), .A2(n_740), .B1(n_741), .B2(n_743), .Y(n_739) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_460), .Y(n_439) );
AND2x2_ASAP7_75t_L g555 ( .A(n_440), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_440), .B(n_602), .Y(n_621) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g539 ( .A(n_441), .Y(n_539) );
AND2x2_ASAP7_75t_L g589 ( .A(n_441), .B(n_462), .Y(n_589) );
INVx1_ASAP7_75t_L g628 ( .A(n_441), .Y(n_628) );
OR2x2_ASAP7_75t_L g665 ( .A(n_441), .B(n_477), .Y(n_665) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_441), .Y(n_677) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_441), .Y(n_701) );
AND2x2_ASAP7_75t_L g758 ( .A(n_441), .B(n_585), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g509 ( .A(n_444), .Y(n_509) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g545 ( .A(n_445), .Y(n_545) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
OR2x6_ASAP7_75t_L g457 ( .A(n_446), .B(n_454), .Y(n_457) );
INVxp33_ASAP7_75t_L g519 ( .A(n_446), .Y(n_519) );
INVx1_ASAP7_75t_L g546 ( .A(n_448), .Y(n_546) );
INVxp67_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
NOR2x1p5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g520 ( .A(n_453), .Y(n_520) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_457), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_465) );
INVxp67_ASAP7_75t_L g498 ( .A(n_457), .Y(n_498) );
INVx2_ASAP7_75t_L g552 ( .A(n_457), .Y(n_552) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_475), .Y(n_460) );
INVx1_ASAP7_75t_L g633 ( .A(n_461), .Y(n_633) );
AND2x2_ASAP7_75t_L g659 ( .A(n_461), .B(n_477), .Y(n_659) );
NAND2x1_ASAP7_75t_L g675 ( .A(n_461), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g556 ( .A(n_462), .B(n_542), .Y(n_556) );
INVx3_ASAP7_75t_L g585 ( .A(n_462), .Y(n_585) );
NOR2x1_ASAP7_75t_SL g704 ( .A(n_462), .B(n_477), .Y(n_704) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_469), .B(n_474), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_468), .B(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_469) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_475), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g583 ( .A(n_476), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g553 ( .A(n_477), .Y(n_553) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_477), .Y(n_598) );
AND2x2_ASAP7_75t_L g670 ( .A(n_477), .B(n_542), .Y(n_670) );
AND2x4_ASAP7_75t_L g687 ( .A(n_477), .B(n_631), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_477), .B(n_629), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_477), .B(n_538), .Y(n_763) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_485), .A2(n_580), .B1(n_651), .B2(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_510), .Y(n_485) );
INVx2_ASAP7_75t_L g653 ( .A(n_486), .Y(n_653) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_494), .Y(n_486) );
BUFx3_ASAP7_75t_L g643 ( .A(n_487), .Y(n_643) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_488), .B(n_512), .Y(n_535) );
INVx2_ASAP7_75t_L g559 ( .A(n_488), .Y(n_559) );
INVx1_ASAP7_75t_L g571 ( .A(n_488), .Y(n_571) );
AND2x4_ASAP7_75t_L g578 ( .A(n_488), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g595 ( .A(n_488), .B(n_495), .Y(n_595) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_488), .Y(n_609) );
INVxp67_ASAP7_75t_L g617 ( .A(n_488), .Y(n_617) );
AND2x2_ASAP7_75t_L g646 ( .A(n_494), .B(n_562), .Y(n_646) );
AND2x2_ASAP7_75t_L g662 ( .A(n_494), .B(n_563), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g749 ( .A(n_494), .B(n_562), .Y(n_749) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g558 ( .A(n_495), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
INVx1_ASAP7_75t_L g582 ( .A(n_495), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_495), .B(n_524), .Y(n_619) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g742 ( .A(n_510), .Y(n_742) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_523), .Y(n_510) );
AND2x2_ASAP7_75t_L g616 ( .A(n_511), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g645 ( .A(n_511), .Y(n_645) );
AND2x2_ASAP7_75t_L g747 ( .A(n_511), .B(n_562), .Y(n_747) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_512), .B(n_524), .Y(n_607) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_522), .Y(n_512) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_513), .A2(n_514), .B(n_522), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_515), .B(n_521), .Y(n_514) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g533 ( .A(n_523), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g722 ( .A(n_523), .B(n_643), .Y(n_722) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_524), .Y(n_636) );
AND2x2_ASAP7_75t_L g663 ( .A(n_524), .B(n_609), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_L g577 ( .A(n_533), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
AND2x2_ASAP7_75t_L g681 ( .A(n_533), .B(n_558), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_533), .B(n_701), .Y(n_706) );
AND2x2_ASAP7_75t_L g716 ( .A(n_533), .B(n_595), .Y(n_716) );
OR2x2_ASAP7_75t_L g753 ( .A(n_533), .B(n_653), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_534), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g713 ( .A(n_534), .B(n_569), .Y(n_713) );
AND2x2_ASAP7_75t_L g729 ( .A(n_534), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g723 ( .A(n_535), .B(n_619), .Y(n_723) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g605 ( .A(n_537), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_537), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g703 ( .A(n_537), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_537), .B(n_584), .Y(n_728) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_538), .Y(n_575) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_539), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_540), .A2(n_573), .B1(n_591), .B2(n_594), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_540), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g707 ( .A(n_540), .Y(n_707) );
AND2x4_ASAP7_75t_SL g540 ( .A(n_541), .B(n_553), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g584 ( .A(n_542), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g604 ( .A(n_542), .Y(n_604) );
INVx1_ASAP7_75t_L g631 ( .A(n_542), .Y(n_631) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .C(n_547), .Y(n_544) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_553), .Y(n_573) );
AND2x4_ASAP7_75t_L g630 ( .A(n_553), .B(n_631), .Y(n_630) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_553), .B(n_660), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
AND2x2_ASAP7_75t_L g655 ( .A(n_555), .B(n_598), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g735 ( .A1(n_555), .A2(n_736), .B(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g613 ( .A(n_556), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_557), .A2(n_667), .B1(n_671), .B2(n_674), .Y(n_666) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_558), .Y(n_624) );
AND2x2_ASAP7_75t_L g634 ( .A(n_558), .B(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g673 ( .A(n_558), .Y(n_673) );
NAND2x1_ASAP7_75t_SL g698 ( .A(n_558), .B(n_567), .Y(n_698) );
AND2x2_ASAP7_75t_L g594 ( .A(n_560), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_562), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g567 ( .A(n_563), .Y(n_567) );
INVx2_ASAP7_75t_L g579 ( .A(n_563), .Y(n_579) );
AOI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_572), .B(n_576), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_567), .B(n_761), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_568), .A2(n_657), .B1(n_661), .B2(n_664), .Y(n_656) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
BUFx2_ASAP7_75t_L g761 ( .A(n_569), .Y(n_761) );
INVx1_ASAP7_75t_SL g768 ( .A(n_569), .Y(n_768) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_570), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OA21x2_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B(n_583), .Y(n_576) );
AND2x2_ASAP7_75t_L g580 ( .A(n_578), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g622 ( .A(n_578), .B(n_618), .Y(n_622) );
AND2x2_ASAP7_75t_L g737 ( .A(n_578), .B(n_635), .Y(n_737) );
AND2x2_ASAP7_75t_L g740 ( .A(n_578), .B(n_646), .Y(n_740) );
AND2x4_ASAP7_75t_L g748 ( .A(n_578), .B(n_749), .Y(n_748) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_580), .A2(n_703), .B(n_705), .Y(n_702) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g730 ( .A(n_582), .Y(n_730) );
AND2x2_ASAP7_75t_L g746 ( .A(n_582), .B(n_747), .Y(n_746) );
INVx4_ASAP7_75t_L g660 ( .A(n_584), .Y(n_660) );
INVx1_ASAP7_75t_L g629 ( .A(n_585), .Y(n_629) );
AND2x2_ASAP7_75t_L g651 ( .A(n_585), .B(n_604), .Y(n_651) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_610), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_590), .B(n_596), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g597 ( .A(n_589), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_SL g750 ( .A(n_589), .B(n_602), .Y(n_750) );
AND2x2_ASAP7_75t_L g771 ( .A(n_589), .B(n_687), .Y(n_771) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g697 ( .A(n_594), .Y(n_697) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_606), .Y(n_596) );
OR2x6_ASAP7_75t_L g649 ( .A(n_598), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g672 ( .A(n_607), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g769 ( .A(n_607), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_608), .B(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_623), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B1(n_620), .B2(n_622), .Y(n_611) );
OR2x2_ASAP7_75t_L g683 ( .A(n_613), .B(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_615), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g689 ( .A(n_618), .Y(n_689) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_632), .B2(n_634), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
AND2x4_ASAP7_75t_SL g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g632 ( .A(n_630), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g693 ( .A(n_633), .B(n_687), .Y(n_693) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_678), .Y(n_637) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_639), .B(n_652), .Y(n_638) );
AOI21xp33_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_641), .B(n_647), .Y(n_639) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp33_ASAP7_75t_SL g717 ( .A1(n_649), .A2(n_718), .B1(n_720), .B2(n_723), .Y(n_717) );
NOR2x1_ASAP7_75t_L g664 ( .A(n_650), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g700 ( .A(n_651), .B(n_701), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_666), .Y(n_652) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVxp33_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g669 ( .A(n_660), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_661), .A2(n_681), .B1(n_682), .B2(n_685), .C(n_688), .Y(n_680) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g721 ( .A(n_662), .Y(n_721) );
INVx2_ASAP7_75t_SL g719 ( .A(n_665), .Y(n_719) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND2x1_ASAP7_75t_L g718 ( .A(n_669), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g715 ( .A(n_675), .Y(n_715) );
INVx1_ASAP7_75t_L g744 ( .A(n_676), .Y(n_744) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_694), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_692), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g733 ( .A(n_684), .Y(n_733) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g754 ( .A(n_687), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g759 ( .A(n_687), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVxp33_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g712 ( .A(n_691), .Y(n_712) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_699), .B(n_702), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g755 ( .A(n_701), .Y(n_755) );
AND2x2_ASAP7_75t_L g743 ( .A(n_704), .B(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_R g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_724), .C(n_751), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_717), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_714), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_738), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_726), .B(n_735), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_734), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_739), .B(n_745), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_748), .B(n_750), .Y(n_745) );
INVx1_ASAP7_75t_L g764 ( .A(n_748), .Y(n_764) );
AOI211xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B(n_756), .C(n_765), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_760), .B1(n_762), .B2(n_764), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_770), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVxp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_786), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_787), .A2(n_800), .B(n_802), .Y(n_799) );
NOR2xp33_ASAP7_75t_SL g787 ( .A(n_788), .B(n_793), .Y(n_787) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
BUFx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
BUFx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g803 ( .A(n_792), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_799), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
CKINVDCx8_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
BUFx4f_ASAP7_75t_SL g816 ( .A(n_807), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g807 ( .A(n_808), .B(n_812), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
endmodule