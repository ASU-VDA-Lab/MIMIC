module real_aes_7991_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_88), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g444 ( .A(n_0), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_1), .A2(n_149), .B(n_154), .C(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_2), .A2(n_144), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g464 ( .A(n_3), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_4), .B(n_168), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_5), .A2(n_16), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_5), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_6), .A2(n_144), .B(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_L g149 ( .A(n_7), .B(n_150), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_8), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_8), .Y(n_726) );
INVx1_ASAP7_75t_L g178 ( .A(n_9), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_10), .B(n_45), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_11), .A2(n_256), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_12), .B(n_159), .Y(n_195) );
INVx1_ASAP7_75t_L g486 ( .A(n_13), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_14), .B(n_158), .Y(n_534) );
INVx1_ASAP7_75t_L g142 ( .A(n_15), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_16), .Y(n_731) );
INVx1_ASAP7_75t_L g546 ( .A(n_17), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_18), .A2(n_179), .B(n_204), .C(n_206), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_19), .B(n_168), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_20), .B(n_475), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_21), .B(n_144), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_22), .B(n_264), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_23), .A2(n_158), .B(n_160), .C(n_164), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_24), .A2(n_49), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_24), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_24), .B(n_168), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_25), .B(n_159), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_26), .A2(n_162), .B(n_206), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_27), .B(n_159), .Y(n_240) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_28), .Y(n_224) );
INVx1_ASAP7_75t_L g238 ( .A(n_29), .Y(n_238) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_31), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_32), .B(n_159), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_33), .A2(n_449), .B1(n_724), .B2(n_725), .C1(n_734), .C2(n_735), .Y(n_448) );
INVx1_ASAP7_75t_L g261 ( .A(n_34), .Y(n_261) );
INVx1_ASAP7_75t_L g499 ( .A(n_35), .Y(n_499) );
INVx2_ASAP7_75t_L g147 ( .A(n_36), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_37), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_38), .A2(n_158), .B(n_217), .C(n_219), .Y(n_216) );
INVxp67_ASAP7_75t_L g262 ( .A(n_39), .Y(n_262) );
CKINVDCx14_ASAP7_75t_R g215 ( .A(n_40), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_41), .A2(n_154), .B(n_237), .C(n_243), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_42), .A2(n_149), .B(n_154), .C(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_43), .A2(n_93), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_43), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_44), .A2(n_105), .B1(n_114), .B2(n_739), .Y(n_104) );
INVx1_ASAP7_75t_L g498 ( .A(n_46), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_47), .A2(n_176), .B(n_177), .C(n_180), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_48), .B(n_159), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_49), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_50), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_51), .Y(n_258) );
INVx1_ASAP7_75t_L g152 ( .A(n_52), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_53), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_54), .B(n_144), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_55), .A2(n_154), .B1(n_164), .B2(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_56), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_57), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_58), .Y(n_461) );
CKINVDCx14_ASAP7_75t_R g174 ( .A(n_59), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_60), .A2(n_176), .B(n_219), .C(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_61), .Y(n_527) );
INVx1_ASAP7_75t_L g483 ( .A(n_62), .Y(n_483) );
INVx1_ASAP7_75t_L g150 ( .A(n_63), .Y(n_150) );
INVx1_ASAP7_75t_L g141 ( .A(n_64), .Y(n_141) );
INVx1_ASAP7_75t_SL g218 ( .A(n_65), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_67), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g227 ( .A(n_68), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_SL g474 ( .A1(n_69), .A2(n_219), .B(n_475), .C(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g477 ( .A(n_70), .Y(n_477) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_72), .A2(n_144), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_73), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_74), .A2(n_144), .B(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_75), .Y(n_502) );
INVx1_ASAP7_75t_L g521 ( .A(n_76), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_77), .A2(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g202 ( .A(n_78), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_79), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_80), .A2(n_149), .B(n_154), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_81), .A2(n_144), .B(n_151), .Y(n_143) );
INVx1_ASAP7_75t_L g205 ( .A(n_82), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_83), .B(n_239), .Y(n_515) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
INVx1_ASAP7_75t_L g192 ( .A(n_85), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_86), .B(n_475), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_87), .A2(n_149), .B(n_154), .C(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g441 ( .A(n_88), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g451 ( .A(n_88), .Y(n_451) );
OR2x2_ASAP7_75t_L g723 ( .A(n_88), .B(n_443), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_89), .A2(n_154), .B(n_226), .C(n_229), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_90), .A2(n_729), .B1(n_730), .B2(n_733), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_90), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_91), .B(n_171), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_92), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_93), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_94), .A2(n_149), .B(n_154), .C(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_95), .Y(n_538) );
INVx1_ASAP7_75t_L g473 ( .A(n_96), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_97), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_98), .B(n_239), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_99), .B(n_137), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_100), .B(n_137), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_101), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g161 ( .A(n_102), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_103), .A2(n_144), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g739 ( .A(n_107), .Y(n_739) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g443 ( .A(n_108), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_447), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g738 ( .A(n_117), .Y(n_738) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_439), .B(n_445), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_437), .B2(n_438), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_122), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_125), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_435), .B2(n_436), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_126), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_129), .A2(n_450), .B1(n_452), .B2(n_721), .Y(n_449) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g436 ( .A(n_130), .Y(n_436) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_361), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_303), .C(n_333), .D(n_343), .Y(n_131) );
OAI211xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_208), .B(n_266), .C(n_293), .Y(n_132) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_133), .A2(n_308), .B1(n_389), .B2(n_390), .C1(n_391), .C2(n_392), .Y(n_388) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_183), .Y(n_133) );
AOI33xp33_ASAP7_75t_L g314 ( .A1(n_134), .A2(n_301), .A3(n_302), .B1(n_315), .B2(n_320), .B3(n_322), .Y(n_314) );
OAI211xp5_ASAP7_75t_SL g371 ( .A1(n_134), .A2(n_372), .B(n_374), .C(n_376), .Y(n_371) );
OR2x2_ASAP7_75t_L g387 ( .A(n_134), .B(n_373), .Y(n_387) );
INVx1_ASAP7_75t_L g420 ( .A(n_134), .Y(n_420) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_170), .Y(n_134) );
INVx2_ASAP7_75t_L g297 ( .A(n_135), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_135), .B(n_199), .Y(n_313) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_135), .Y(n_348) );
AND2x2_ASAP7_75t_L g377 ( .A(n_135), .B(n_170), .Y(n_377) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_167), .Y(n_135) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_136), .A2(n_200), .B(n_207), .Y(n_199) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_136), .A2(n_213), .B(n_221), .Y(n_212) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx4_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_137), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g254 ( .A(n_138), .Y(n_254) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_139), .B(n_140), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx2_ASAP7_75t_L g256 ( .A(n_144), .Y(n_256) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_145), .B(n_149), .Y(n_189) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g242 ( .A(n_146), .Y(n_242) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
INVx1_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx3_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx1_ASAP7_75t_L g475 ( .A(n_148), .Y(n_475) );
INVx4_ASAP7_75t_SL g166 ( .A(n_149), .Y(n_166) );
BUFx3_ASAP7_75t_L g243 ( .A(n_149), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_153), .B(n_157), .C(n_166), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_153), .A2(n_166), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_153), .A2(n_166), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_153), .A2(n_166), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_153), .A2(n_166), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_153), .A2(n_166), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_153), .A2(n_166), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_153), .A2(n_166), .B(n_543), .C(n_544), .Y(n_542) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_158), .B(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_162), .B(n_205), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_162), .A2(n_239), .B1(n_261), .B2(n_262), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_162), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_163), .A2(n_194), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g466 ( .A(n_164), .Y(n_466) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_166), .A2(n_189), .B1(n_496), .B2(n_500), .Y(n_495) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_168), .A2(n_481), .B(n_487), .Y(n_480) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_169), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_169), .A2(n_223), .B(n_230), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_169), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_SL g517 ( .A(n_169), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g277 ( .A(n_170), .Y(n_277) );
BUFx3_ASAP7_75t_L g285 ( .A(n_170), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_170), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g296 ( .A(n_170), .B(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_170), .B(n_184), .Y(n_325) );
AND2x2_ASAP7_75t_L g394 ( .A(n_170), .B(n_328), .Y(n_394) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_182), .Y(n_170) );
INVx1_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx2_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_171), .A2(n_189), .B(n_235), .C(n_236), .Y(n_234) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_171), .A2(n_541), .B(n_547), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx5_ASAP7_75t_L g239 ( .A(n_179), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_179), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_179), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g196 ( .A(n_180), .Y(n_196) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g206 ( .A(n_181), .Y(n_206) );
INVx2_ASAP7_75t_SL g288 ( .A(n_183), .Y(n_288) );
OR2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_184), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g330 ( .A(n_184), .Y(n_330) );
AND2x2_ASAP7_75t_L g341 ( .A(n_184), .B(n_297), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_184), .B(n_326), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_184), .B(n_328), .Y(n_373) );
AND2x2_ASAP7_75t_L g432 ( .A(n_184), .B(n_377), .Y(n_432) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g302 ( .A(n_185), .B(n_199), .Y(n_302) );
AND2x2_ASAP7_75t_L g312 ( .A(n_185), .B(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g334 ( .A(n_185), .Y(n_334) );
AND3x2_ASAP7_75t_L g393 ( .A(n_185), .B(n_394), .C(n_395), .Y(n_393) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_186), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_186), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_186), .B(n_538), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_189), .A2(n_224), .B(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_189), .A2(n_461), .B(n_462), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_189), .A2(n_521), .B(n_522), .Y(n_520) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_193), .A2(n_196), .B(n_227), .C(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_196), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_196), .A2(n_524), .B(n_525), .Y(n_523) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
INVx1_ASAP7_75t_SL g328 ( .A(n_199), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_199), .B(n_277), .C(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_246), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_209), .A2(n_312), .B(n_364), .C(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_211), .B(n_233), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_211), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g380 ( .A(n_211), .Y(n_380) );
AND2x2_ASAP7_75t_L g401 ( .A(n_211), .B(n_248), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_211), .B(n_310), .Y(n_429) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AND2x2_ASAP7_75t_L g274 ( .A(n_212), .B(n_265), .Y(n_274) );
INVx2_ASAP7_75t_L g281 ( .A(n_212), .Y(n_281) );
AND2x2_ASAP7_75t_L g301 ( .A(n_212), .B(n_248), .Y(n_301) );
AND2x2_ASAP7_75t_L g351 ( .A(n_212), .B(n_233), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_212), .Y(n_355) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_220), .Y(n_535) );
INVx2_ASAP7_75t_SL g265 ( .A(n_222), .Y(n_265) );
BUFx2_ASAP7_75t_L g291 ( .A(n_222), .Y(n_291) );
AND2x2_ASAP7_75t_L g418 ( .A(n_222), .B(n_233), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g264 ( .A(n_232), .Y(n_264) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_232), .A2(n_530), .B(n_537), .Y(n_529) );
INVx3_ASAP7_75t_SL g248 ( .A(n_233), .Y(n_248) );
AND2x2_ASAP7_75t_L g273 ( .A(n_233), .B(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g280 ( .A(n_233), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g310 ( .A(n_233), .B(n_270), .Y(n_310) );
OR2x2_ASAP7_75t_L g319 ( .A(n_233), .B(n_265), .Y(n_319) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
AND2x2_ASAP7_75t_L g342 ( .A(n_233), .B(n_295), .Y(n_342) );
AND2x2_ASAP7_75t_L g370 ( .A(n_233), .B(n_250), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_233), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g408 ( .A(n_233), .B(n_249), .Y(n_408) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_244), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .C(n_241), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_239), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_242), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g332 ( .A(n_248), .B(n_281), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_248), .B(n_274), .Y(n_360) );
AND2x2_ASAP7_75t_L g378 ( .A(n_248), .B(n_295), .Y(n_378) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_265), .Y(n_249) );
AND2x2_ASAP7_75t_L g279 ( .A(n_250), .B(n_265), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_250), .B(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g317 ( .A(n_250), .Y(n_317) );
OR2x2_ASAP7_75t_L g365 ( .A(n_250), .B(n_285), .Y(n_365) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_255), .B(n_263), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_252), .A2(n_271), .B(n_272), .Y(n_270) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_252), .A2(n_520), .B(n_526), .Y(n_519) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI21xp5_ASAP7_75t_SL g511 ( .A1(n_253), .A2(n_512), .B(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_254), .A2(n_460), .B(n_467), .Y(n_459) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_254), .A2(n_495), .B(n_501), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_254), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
AND2x2_ASAP7_75t_L g300 ( .A(n_265), .B(n_270), .Y(n_300) );
INVx1_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_265), .B(n_281), .Y(n_403) );
AOI222xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_275), .B1(n_278), .B2(n_282), .C1(n_286), .C2(n_289), .Y(n_266) );
INVx1_ASAP7_75t_L g398 ( .A(n_267), .Y(n_398) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_273), .Y(n_267) );
AND2x2_ASAP7_75t_L g294 ( .A(n_268), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g305 ( .A(n_268), .B(n_274), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_268), .B(n_296), .Y(n_321) );
OAI222xp33_ASAP7_75t_L g343 ( .A1(n_268), .A2(n_344), .B1(n_349), .B2(n_350), .C1(n_358), .C2(n_360), .Y(n_343) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g331 ( .A(n_270), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_270), .B(n_351), .Y(n_391) );
AND2x2_ASAP7_75t_L g402 ( .A(n_270), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g410 ( .A(n_273), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_275), .B(n_326), .Y(n_389) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_277), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g347 ( .A(n_277), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx3_ASAP7_75t_L g292 ( .A(n_280), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_280), .A2(n_383), .B(n_386), .C(n_388), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_280), .B(n_317), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_280), .B(n_300), .Y(n_422) );
AND2x2_ASAP7_75t_L g295 ( .A(n_281), .B(n_291), .Y(n_295) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_285), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g374 ( .A(n_285), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g413 ( .A(n_285), .B(n_313), .Y(n_413) );
INVx1_ASAP7_75t_L g425 ( .A(n_285), .Y(n_425) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_288), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g406 ( .A(n_291), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_298), .C(n_302), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_294), .A2(n_324), .B1(n_339), .B2(n_342), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_295), .B(n_309), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_295), .B(n_317), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_296), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g359 ( .A(n_296), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_296), .B(n_346), .Y(n_366) );
INVx2_ASAP7_75t_L g327 ( .A(n_297), .Y(n_327) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NOR4xp25_ASAP7_75t_L g304 ( .A(n_301), .B(n_305), .C(n_306), .D(n_309), .Y(n_304) );
INVx1_ASAP7_75t_SL g375 ( .A(n_302), .Y(n_375) );
AND2x2_ASAP7_75t_L g419 ( .A(n_302), .B(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_311), .B(n_314), .C(n_323), .Y(n_303) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_310), .B(n_380), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_312), .A2(n_431), .B1(n_432), .B2(n_433), .Y(n_430) );
INVx1_ASAP7_75t_SL g385 ( .A(n_313), .Y(n_385) );
AND2x2_ASAP7_75t_L g424 ( .A(n_313), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_317), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_321), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_322), .B(n_347), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_329), .B(n_331), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g399 ( .A(n_326), .Y(n_399) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g427 ( .A(n_327), .Y(n_427) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_328), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B(n_338), .Y(n_333) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_334), .Y(n_346) );
OR2x2_ASAP7_75t_L g384 ( .A(n_334), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI21xp33_ASAP7_75t_SL g379 ( .A1(n_337), .A2(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_341), .A2(n_368), .B1(n_371), .B2(n_378), .C(n_379), .Y(n_367) );
INVx1_ASAP7_75t_SL g411 ( .A(n_342), .Y(n_411) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OR2x2_ASAP7_75t_L g358 ( .A(n_346), .B(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_355), .B2(n_356), .Y(n_350) );
INVx1_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_354), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_396), .C(n_409), .D(n_421), .Y(n_361) );
NAND3xp33_ASAP7_75t_SL g362 ( .A(n_363), .B(n_367), .C(n_382), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_365), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_372), .B(n_377), .Y(n_381) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_384), .A2(n_410), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_409) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_386), .A2(n_401), .B(n_402), .C(n_404), .Y(n_400) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_387), .A2(n_405), .B1(n_407), .B2(n_408), .Y(n_404) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_399), .C(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g415 ( .A(n_408), .Y(n_415) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_423), .B1(n_426), .B2(n_428), .C(n_430), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_436), .A2(n_450), .B1(n_453), .B2(n_723), .Y(n_734) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g446 ( .A(n_440), .Y(n_446) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_442), .B(n_451), .Y(n_737) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g450 ( .A(n_443), .B(n_451), .Y(n_450) );
AOI21xp33_ASAP7_75t_SL g447 ( .A1(n_445), .A2(n_448), .B(n_738), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_637), .Y(n_453) );
NOR5xp2_ASAP7_75t_L g454 ( .A(n_455), .B(n_560), .C(n_592), .D(n_607), .E(n_624), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_488), .B(n_507), .C(n_548), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_469), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_457), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_457), .B(n_612), .Y(n_675) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_458), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_458), .B(n_504), .Y(n_561) );
AND2x2_ASAP7_75t_L g602 ( .A(n_458), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_458), .B(n_571), .Y(n_606) );
OR2x2_ASAP7_75t_L g643 ( .A(n_458), .B(n_494), .Y(n_643) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g493 ( .A(n_459), .B(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g551 ( .A(n_459), .Y(n_551) );
OR2x2_ASAP7_75t_L g714 ( .A(n_459), .B(n_554), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_469), .A2(n_617), .B1(n_618), .B2(n_621), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_469), .B(n_551), .Y(n_700) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
AND2x2_ASAP7_75t_L g506 ( .A(n_470), .B(n_494), .Y(n_506) );
AND2x2_ASAP7_75t_L g553 ( .A(n_470), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g558 ( .A(n_470), .Y(n_558) );
INVx3_ASAP7_75t_L g571 ( .A(n_470), .Y(n_571) );
OR2x2_ASAP7_75t_L g591 ( .A(n_470), .B(n_554), .Y(n_591) );
AND2x2_ASAP7_75t_L g610 ( .A(n_470), .B(n_480), .Y(n_610) );
BUFx2_ASAP7_75t_L g642 ( .A(n_470), .Y(n_642) );
AND2x4_ASAP7_75t_L g557 ( .A(n_479), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g492 ( .A(n_480), .Y(n_492) );
INVx2_ASAP7_75t_L g505 ( .A(n_480), .Y(n_505) );
OR2x2_ASAP7_75t_L g573 ( .A(n_480), .B(n_554), .Y(n_573) );
AND2x2_ASAP7_75t_L g603 ( .A(n_480), .B(n_494), .Y(n_603) );
AND2x2_ASAP7_75t_L g620 ( .A(n_480), .B(n_551), .Y(n_620) );
AND2x2_ASAP7_75t_L g660 ( .A(n_480), .B(n_571), .Y(n_660) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_480), .B(n_506), .Y(n_696) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp33_ASAP7_75t_SL g489 ( .A(n_490), .B(n_503), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_491), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_492), .A2(n_506), .B(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_492), .B(n_494), .Y(n_690) );
AND2x2_ASAP7_75t_L g626 ( .A(n_493), .B(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g554 ( .A(n_494), .Y(n_554) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_494), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_503), .B(n_551), .Y(n_719) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_504), .A2(n_662), .B1(n_663), .B2(n_668), .Y(n_661) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g552 ( .A(n_505), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g590 ( .A(n_505), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g627 ( .A(n_505), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_506), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g681 ( .A(n_506), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_528), .Y(n_508) );
INVx4_ASAP7_75t_L g567 ( .A(n_509), .Y(n_567) );
AND2x2_ASAP7_75t_L g645 ( .A(n_509), .B(n_612), .Y(n_645) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
INVx3_ASAP7_75t_L g564 ( .A(n_510), .Y(n_564) );
AND2x2_ASAP7_75t_L g578 ( .A(n_510), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
INVx2_ASAP7_75t_L g596 ( .A(n_510), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_510), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g653 ( .A(n_510), .B(n_648), .Y(n_653) );
AND2x2_ASAP7_75t_L g718 ( .A(n_510), .B(n_688), .Y(n_718) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_517), .Y(n_510) );
AND2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_540), .Y(n_559) );
INVx2_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g630 ( .A(n_528), .B(n_578), .Y(n_630) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
INVx2_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
INVx1_ASAP7_75t_L g577 ( .A(n_529), .Y(n_577) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_529), .B(n_579), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g612 ( .A(n_539), .B(n_569), .Y(n_612) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
AND2x2_ASAP7_75t_L g648 ( .A(n_540), .B(n_579), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_555), .B(n_559), .Y(n_548) );
INVx1_ASAP7_75t_SL g593 ( .A(n_549), .Y(n_593) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_550), .B(n_557), .Y(n_650) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g599 ( .A(n_551), .B(n_554), .Y(n_599) );
AND2x2_ASAP7_75t_L g628 ( .A(n_551), .B(n_572), .Y(n_628) );
OR2x2_ASAP7_75t_L g631 ( .A(n_551), .B(n_591), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_552), .A2(n_644), .B1(n_696), .B2(n_697), .C1(n_699), .C2(n_701), .Y(n_695) );
BUFx2_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g598 ( .A(n_557), .B(n_599), .Y(n_598) );
INVx3_ASAP7_75t_SL g615 ( .A(n_557), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_557), .B(n_609), .Y(n_669) );
AND2x2_ASAP7_75t_L g604 ( .A(n_559), .B(n_564), .Y(n_604) );
INVx1_ASAP7_75t_L g623 ( .A(n_559), .Y(n_623) );
OAI221xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_562), .B1(n_566), .B2(n_570), .C(n_574), .Y(n_560) );
OR2x2_ASAP7_75t_L g632 ( .A(n_562), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_587), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_564), .B(n_577), .Y(n_657) );
AND2x2_ASAP7_75t_L g662 ( .A(n_564), .B(n_612), .Y(n_662) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_564), .Y(n_672) );
NAND2x1_ASAP7_75t_SL g683 ( .A(n_564), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g568 ( .A(n_565), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g588 ( .A(n_565), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_565), .B(n_583), .Y(n_614) );
INVx1_ASAP7_75t_L g680 ( .A(n_565), .Y(n_680) );
INVx1_ASAP7_75t_L g655 ( .A(n_566), .Y(n_655) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g667 ( .A(n_567), .Y(n_667) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_567), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g684 ( .A(n_568), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_568), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g587 ( .A(n_569), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_569), .B(n_579), .Y(n_600) );
INVx1_ASAP7_75t_L g666 ( .A(n_569), .Y(n_666) );
INVx1_ASAP7_75t_L g687 ( .A(n_570), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_580), .B(n_589), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
AND2x2_ASAP7_75t_L g720 ( .A(n_576), .B(n_653), .Y(n_720) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g688 ( .A(n_577), .B(n_648), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g601 ( .A1(n_578), .A2(n_584), .A3(n_602), .B1(n_604), .B2(n_605), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g703 ( .A1(n_578), .A2(n_610), .A3(n_693), .B1(n_704), .B2(n_705), .C1(n_706), .C2(n_708), .Y(n_703) );
INVx2_ASAP7_75t_L g583 ( .A(n_579), .Y(n_583) );
INVx1_ASAP7_75t_L g693 ( .A(n_579), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_581), .B(n_587), .Y(n_636) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_582), .B(n_648), .Y(n_698) );
INVx1_ASAP7_75t_L g585 ( .A(n_583), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_583), .B(n_612), .Y(n_702) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_591), .B(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_597), .B2(n_600), .C(n_601), .Y(n_592) );
OR2x2_ASAP7_75t_L g613 ( .A(n_594), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g622 ( .A(n_594), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g647 ( .A(n_595), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g651 ( .A(n_605), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B1(n_613), .B2(n_615), .C(n_616), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_609), .A2(n_640), .B1(n_644), .B2(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_610), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g715 ( .A(n_610), .Y(n_715) );
INVx1_ASAP7_75t_L g709 ( .A(n_612), .Y(n_709) );
INVx1_ASAP7_75t_SL g644 ( .A(n_613), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_615), .B(n_643), .Y(n_705) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_620), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g686 ( .A(n_620), .Y(n_686) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_629), .B1(n_631), .B2(n_632), .C(n_634), .Y(n_624) );
NOR2xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_628), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_626), .A2(n_644), .B1(n_690), .B2(n_691), .Y(n_689) );
CKINVDCx14_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_631), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR3xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_670), .C(n_694), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_639), .B(n_646), .C(n_654), .D(n_661), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g717 ( .A(n_642), .Y(n_717) );
INVx3_ASAP7_75t_SL g711 ( .A(n_643), .Y(n_711) );
OR2x2_ASAP7_75t_L g716 ( .A(n_643), .B(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_651), .B2(n_653), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_648), .B(n_666), .Y(n_707) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_656), .B(n_658), .Y(n_654) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_676), .C(n_689), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g704 ( .A(n_675), .Y(n_704) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_681), .B1(n_682), .B2(n_685), .C1(n_687), .C2(n_688), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND4xp25_ASAP7_75t_SL g713 ( .A(n_686), .B(n_714), .C(n_715), .D(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND3xp33_ASAP7_75t_SL g694 ( .A(n_695), .B(n_703), .C(n_712), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_712) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
endmodule