module real_aes_16769_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_842, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_842;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_0), .Y(n_159) );
AND2x4_ASAP7_75t_L g837 ( .A(n_1), .B(n_838), .Y(n_837) );
BUFx3_ASAP7_75t_L g210 ( .A(n_2), .Y(n_210) );
INVx1_ASAP7_75t_L g838 ( .A(n_3), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_4), .A2(n_130), .B1(n_827), .B2(n_828), .Y(n_826) );
INVxp67_ASAP7_75t_SL g827 ( .A(n_4), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_5), .B(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g111 ( .A(n_6), .B(n_23), .Y(n_111) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_7), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_8), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_9), .A2(n_122), .B1(n_123), .B2(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_9), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_10), .B(n_180), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_11), .B(n_180), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_12), .B(n_140), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_13), .A2(n_80), .B1(n_177), .B2(n_180), .Y(n_179) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_14), .A2(n_36), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_15), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_16), .B(n_149), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_17), .Y(n_552) );
AO32x1_ASAP7_75t_L g171 ( .A1(n_18), .A2(n_172), .A3(n_173), .B1(n_182), .B2(n_184), .Y(n_171) );
AO32x2_ASAP7_75t_L g288 ( .A1(n_18), .A2(n_172), .A3(n_173), .B1(n_182), .B2(n_184), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_19), .B(n_512), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_20), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_21), .B(n_184), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_22), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_24), .A2(n_42), .B1(n_149), .B2(n_151), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_25), .A2(n_88), .B1(n_177), .B2(n_178), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_26), .B(n_220), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_27), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_28), .B(n_245), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_29), .A2(n_61), .B1(n_178), .B2(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_30), .B(n_180), .Y(n_498) );
INVx2_ASAP7_75t_L g117 ( .A(n_31), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_32), .B(n_181), .Y(n_508) );
INVx1_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
BUFx3_ASAP7_75t_L g120 ( .A(n_33), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_34), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_35), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g557 ( .A(n_37), .B(n_517), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_38), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_39), .B(n_160), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_40), .B(n_512), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_41), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_43), .B(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_44), .A2(n_75), .B1(n_160), .B2(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_45), .B(n_189), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_46), .A2(n_157), .B(n_174), .C(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_47), .A2(n_77), .B1(n_177), .B2(n_180), .Y(n_206) );
INVx1_ASAP7_75t_L g144 ( .A(n_48), .Y(n_144) );
AND2x4_ASAP7_75t_L g164 ( .A(n_49), .B(n_165), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_50), .A2(n_51), .B1(n_151), .B2(n_178), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_52), .B(n_184), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_53), .B(n_517), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_54), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_55), .B(n_178), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_56), .B(n_177), .Y(n_216) );
INVx1_ASAP7_75t_L g165 ( .A(n_57), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_58), .B(n_184), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_59), .A2(n_157), .B(n_158), .C(n_161), .Y(n_156) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_60), .B(n_177), .C(n_222), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_62), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_63), .B(n_184), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_64), .B(n_501), .Y(n_539) );
AND2x2_ASAP7_75t_L g166 ( .A(n_65), .B(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_66), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_67), .B(n_149), .C(n_181), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_68), .A2(n_100), .B1(n_830), .B2(n_839), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_69), .A2(n_91), .B1(n_160), .B2(n_180), .Y(n_247) );
INVx2_ASAP7_75t_L g155 ( .A(n_70), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_71), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_72), .B(n_501), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_73), .B(n_154), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_74), .B(n_180), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_76), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_78), .B(n_237), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_79), .A2(n_87), .B1(n_512), .B2(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_81), .B(n_180), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_82), .B(n_222), .Y(n_221) );
NAND2xp33_ASAP7_75t_SL g580 ( .A(n_83), .B(n_218), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_84), .B(n_233), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_85), .A2(n_98), .B1(n_151), .B2(n_178), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_86), .B(n_245), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_89), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_90), .B(n_140), .Y(n_269) );
NAND2xp33_ASAP7_75t_L g565 ( .A(n_92), .B(n_218), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_93), .B(n_517), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_94), .B(n_154), .C(n_218), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_95), .B(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_96), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_97), .B(n_512), .Y(n_542) );
OR2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_112), .Y(n_100) );
INVxp67_ASAP7_75t_L g829 ( .A(n_101), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
INVx4_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx8_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x6_ASAP7_75t_SL g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_109), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_110), .B(n_119), .Y(n_118) );
AND3x2_ASAP7_75t_L g822 ( .A(n_110), .B(n_823), .C(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_111), .B(n_120), .Y(n_814) );
BUFx2_ASAP7_75t_L g834 ( .A(n_111), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_815), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B(n_807), .Y(n_113) );
BUFx12f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x6_ASAP7_75t_SL g115 ( .A(n_116), .B(n_118), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_117), .B(n_812), .Y(n_811) );
INVx3_ASAP7_75t_L g818 ( .A(n_117), .Y(n_818) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_485), .B2(n_487), .Y(n_126) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_127), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g813 ( .A(n_128), .B(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx2_ASAP7_75t_L g824 ( .A(n_129), .Y(n_824) );
INVx1_ASAP7_75t_L g828 ( .A(n_130), .Y(n_828) );
NAND4xp75_ASAP7_75t_L g130 ( .A(n_131), .B(n_359), .C(n_413), .D(n_457), .Y(n_130) );
NOR2x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_312), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_278), .Y(n_132) );
O2A1O1Ixp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_195), .B(n_199), .C(n_251), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
AND2x2_ASAP7_75t_L g329 ( .A(n_135), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g318 ( .A(n_136), .B(n_254), .Y(n_318) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_137), .Y(n_284) );
AND2x2_ASAP7_75t_L g333 ( .A(n_137), .B(n_185), .Y(n_333) );
INVx1_ASAP7_75t_L g345 ( .A(n_137), .Y(n_345) );
INVx1_ASAP7_75t_L g443 ( .A(n_137), .Y(n_443) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
AOI21x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_166), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp67_ASAP7_75t_SL g547 ( .A(n_140), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AO31x2_ASAP7_75t_L g518 ( .A1(n_141), .A2(n_519), .A3(n_524), .B(n_525), .Y(n_518) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx2_ASAP7_75t_L g213 ( .A(n_142), .Y(n_213) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_156), .B(n_163), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_147), .B(n_153), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B1(n_151), .B2(n_152), .Y(n_147) );
INVx2_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_150), .Y(n_151) );
INVx1_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx1_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
INVx2_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
INVx1_ASAP7_75t_L g233 ( .A(n_150), .Y(n_233) );
INVx3_ASAP7_75t_L g501 ( .A(n_150), .Y(n_501) );
INVx1_ASAP7_75t_L g513 ( .A(n_150), .Y(n_513) );
INVx1_ASAP7_75t_L g239 ( .A(n_151), .Y(n_239) );
AOI21x1_ASAP7_75t_L g510 ( .A1(n_153), .A2(n_511), .B(n_514), .Y(n_510) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g246 ( .A(n_154), .Y(n_246) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
INVx1_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
BUFx8_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
INVx1_ASAP7_75t_L g568 ( .A(n_157), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx2_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
INVx2_ASAP7_75t_L g523 ( .A(n_161), .Y(n_523) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g238 ( .A(n_162), .Y(n_238) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
AO31x2_ASAP7_75t_L g185 ( .A1(n_164), .A2(n_186), .A3(n_187), .B(n_193), .Y(n_185) );
BUFx10_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
BUFx10_ASAP7_75t_L g524 ( .A(n_164), .Y(n_524) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_168), .B(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_168), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g271 ( .A(n_170), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_185), .Y(n_170) );
AND2x2_ASAP7_75t_L g198 ( .A(n_171), .B(n_185), .Y(n_198) );
INVx1_ASAP7_75t_L g311 ( .A(n_171), .Y(n_311) );
INVx1_ASAP7_75t_L g422 ( .A(n_171), .Y(n_422) );
INVx4_ASAP7_75t_L g184 ( .A(n_172), .Y(n_184) );
BUFx3_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_172), .B(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_172), .B(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g228 ( .A(n_172), .Y(n_228) );
INVx2_ASAP7_75t_SL g260 ( .A(n_172), .Y(n_260) );
AND2x4_ASAP7_75t_SL g570 ( .A(n_172), .B(n_204), .Y(n_570) );
INVx1_ASAP7_75t_SL g573 ( .A(n_172), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B1(n_179), .B2(n_181), .Y(n_173) );
O2A1O1Ixp5_ASAP7_75t_L g230 ( .A1(n_174), .A2(n_231), .B(n_232), .C(n_234), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_174), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_174), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_174), .A2(n_564), .B(n_565), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_174), .A2(n_579), .B(n_580), .Y(n_578) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
INVx2_ASAP7_75t_SL g245 ( .A(n_177), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_177), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_178), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g521 ( .A(n_178), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_178), .A2(n_501), .B1(n_555), .B2(n_556), .Y(n_554) );
INVx3_ASAP7_75t_L g268 ( .A(n_180), .Y(n_268) );
INVx1_ASAP7_75t_L g515 ( .A(n_180), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_180), .A2(n_576), .B(n_577), .Y(n_575) );
INVx6_ASAP7_75t_L g190 ( .A(n_181), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_181), .A2(n_190), .B1(n_206), .B2(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_181), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_181), .A2(n_500), .B(n_502), .Y(n_499) );
O2A1O1Ixp5_ASAP7_75t_L g626 ( .A1(n_181), .A2(n_232), .B(n_627), .C(n_628), .Y(n_626) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_182), .A2(n_262), .B(n_265), .Y(n_261) );
INVx2_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_SL g248 ( .A(n_183), .Y(n_248) );
INVx2_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
INVx3_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_185), .B(n_258), .Y(n_309) );
AND2x2_ASAP7_75t_L g344 ( .A(n_185), .B(n_345), .Y(n_344) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_186), .A2(n_243), .A3(n_248), .B(n_249), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_190), .A2(n_244), .B1(n_246), .B2(n_247), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_190), .A2(n_266), .B(n_267), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_190), .A2(n_520), .B1(n_522), .B2(n_523), .Y(n_519) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_192), .A2(n_263), .B(n_264), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_192), .A2(n_542), .B(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_198), .Y(n_195) );
INVx1_ASAP7_75t_L g384 ( .A(n_196), .Y(n_384) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g253 ( .A(n_197), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_197), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g286 ( .A(n_197), .Y(n_286) );
OR2x2_ASAP7_75t_L g350 ( .A(n_197), .B(n_258), .Y(n_350) );
OR2x2_ASAP7_75t_L g421 ( .A(n_197), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g358 ( .A(n_198), .Y(n_358) );
AND2x2_ASAP7_75t_L g410 ( .A(n_198), .B(n_273), .Y(n_410) );
AND2x2_ASAP7_75t_L g467 ( .A(n_198), .B(n_384), .Y(n_467) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_225), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_200), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g476 ( .A(n_200), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
INVx2_ASAP7_75t_L g277 ( .A(n_201), .Y(n_277) );
AND2x2_ASAP7_75t_L g302 ( .A(n_201), .B(n_281), .Y(n_302) );
AND2x2_ASAP7_75t_L g372 ( .A(n_201), .B(n_242), .Y(n_372) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g326 ( .A(n_202), .Y(n_326) );
AOI31xp67_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .A3(n_205), .B(n_208), .Y(n_202) );
OAI21x1_ASAP7_75t_L g214 ( .A1(n_204), .A2(n_215), .B(n_219), .Y(n_214) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_204), .A2(n_230), .B(n_235), .Y(n_229) );
OAI21x1_ASAP7_75t_L g495 ( .A1(n_204), .A2(n_496), .B(n_499), .Y(n_495) );
OAI21x1_ASAP7_75t_L g506 ( .A1(n_204), .A2(n_507), .B(n_510), .Y(n_506) );
OAI21x1_ASAP7_75t_L g537 ( .A1(n_204), .A2(n_538), .B(n_541), .Y(n_537) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_204), .A2(n_575), .B(n_578), .Y(n_574) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_204), .A2(n_626), .B(n_629), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g280 ( .A(n_211), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g341 ( .A(n_211), .B(n_227), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_214), .B(n_224), .Y(n_211) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_212), .A2(n_214), .B(n_224), .Y(n_297) );
OAI21xp33_ASAP7_75t_SL g536 ( .A1(n_212), .A2(n_537), .B(n_544), .Y(n_536) );
OAI21x1_ASAP7_75t_L g606 ( .A1(n_212), .A2(n_537), .B(n_544), .Y(n_606) );
OAI21x1_ASAP7_75t_L g624 ( .A1(n_212), .A2(n_625), .B(n_633), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_212), .A2(n_625), .B(n_633), .Y(n_656) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g517 ( .A(n_213), .Y(n_517) );
INVx2_ASAP7_75t_L g632 ( .A(n_218), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_223), .Y(n_219) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g348 ( .A(n_226), .B(n_325), .Y(n_348) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_242), .Y(n_226) );
INVx2_ASAP7_75t_SL g270 ( .A(n_227), .Y(n_270) );
BUFx2_ASAP7_75t_L g323 ( .A(n_227), .Y(n_323) );
INVx1_ASAP7_75t_L g395 ( .A(n_227), .Y(n_395) );
AND2x2_ASAP7_75t_L g428 ( .A(n_227), .B(n_276), .Y(n_428) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_241), .Y(n_227) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_228), .A2(n_229), .B(n_241), .Y(n_281) );
OAI21x1_ASAP7_75t_L g494 ( .A1(n_228), .A2(n_495), .B(n_503), .Y(n_494) );
OAI21x1_ASAP7_75t_L g505 ( .A1(n_228), .A2(n_506), .B(n_516), .Y(n_505) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_228), .A2(n_495), .B(n_503), .Y(n_586) );
OA21x2_ASAP7_75t_L g621 ( .A1(n_228), .A2(n_506), .B(n_516), .Y(n_621) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_238), .B1(n_239), .B2(n_240), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_237), .A2(n_630), .B(n_631), .Y(n_629) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_238), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_566) );
INVx2_ASAP7_75t_L g256 ( .A(n_242), .Y(n_256) );
INVx1_ASAP7_75t_L g276 ( .A(n_242), .Y(n_276) );
INVx1_ASAP7_75t_L g304 ( .A(n_242), .Y(n_304) );
AND2x2_ASAP7_75t_L g394 ( .A(n_242), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g435 ( .A(n_242), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g451 ( .A(n_242), .B(n_436), .Y(n_451) );
AND2x2_ASAP7_75t_L g477 ( .A(n_242), .B(n_281), .Y(n_477) );
OAI32xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_255), .A3(n_270), .B1(n_271), .B2(n_274), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_253), .B(n_418), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_253), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g287 ( .A(n_254), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g389 ( .A(n_254), .Y(n_389) );
INVx1_ASAP7_75t_L g449 ( .A(n_254), .Y(n_449) );
INVx1_ASAP7_75t_L g387 ( .A(n_255), .Y(n_387) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_SL g291 ( .A(n_256), .Y(n_291) );
AND2x2_ASAP7_75t_L g380 ( .A(n_256), .B(n_295), .Y(n_380) );
AND2x2_ASAP7_75t_L g448 ( .A(n_257), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g273 ( .A(n_258), .Y(n_273) );
AND2x2_ASAP7_75t_L g283 ( .A(n_258), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g319 ( .A(n_258), .Y(n_319) );
AND2x2_ASAP7_75t_L g330 ( .A(n_258), .B(n_288), .Y(n_330) );
AND2x2_ASAP7_75t_L g354 ( .A(n_258), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g364 ( .A(n_258), .B(n_355), .Y(n_364) );
INVxp67_ASAP7_75t_L g418 ( .A(n_258), .Y(n_418) );
BUFx2_ASAP7_75t_L g430 ( .A(n_258), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_258), .Y(n_434) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_269), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_270), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g426 ( .A(n_270), .Y(n_426) );
AND2x2_ASAP7_75t_L g334 ( .A(n_273), .B(n_311), .Y(n_334) );
AND2x2_ASAP7_75t_L g463 ( .A(n_273), .B(n_287), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g351 ( .A1(n_274), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_351) );
O2A1O1Ixp5_ASAP7_75t_R g425 ( .A1(n_274), .A2(n_426), .B(n_427), .C(n_429), .Y(n_425) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g293 ( .A(n_277), .Y(n_293) );
INVx1_ASAP7_75t_L g336 ( .A(n_277), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_277), .B(n_306), .Y(n_412) );
AND2x2_ASAP7_75t_L g424 ( .A(n_277), .B(n_295), .Y(n_424) );
AOI222xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B1(n_285), .B2(n_289), .C1(n_299), .C2(n_307), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_279), .A2(n_321), .B1(n_399), .B2(n_460), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_279), .A2(n_343), .B1(n_479), .B2(n_481), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_280), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_280), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g454 ( .A(n_280), .Y(n_454) );
INVx1_ASAP7_75t_L g484 ( .A(n_280), .Y(n_484) );
INVx1_ASAP7_75t_L g298 ( .A(n_281), .Y(n_298) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
AOI321xp33_ASAP7_75t_L g431 ( .A1(n_285), .A2(n_329), .A3(n_432), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_431) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
OR2x2_ASAP7_75t_L g363 ( .A(n_286), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g383 ( .A(n_287), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g355 ( .A(n_288), .Y(n_355) );
NAND2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
OR2x2_ASAP7_75t_L g356 ( .A(n_291), .B(n_325), .Y(n_356) );
AND2x2_ASAP7_75t_L g376 ( .A(n_291), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g466 ( .A(n_292), .Y(n_466) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g397 ( .A(n_294), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g306 ( .A(n_296), .Y(n_306) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g325 ( .A(n_297), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_300), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_302), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g437 ( .A(n_306), .Y(n_437) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_308), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g370 ( .A(n_309), .Y(n_370) );
INVx1_ASAP7_75t_L g320 ( .A(n_310), .Y(n_320) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
INVx2_ASAP7_75t_L g402 ( .A(n_311), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_337), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_321), .B(n_327), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_320), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_317), .A2(n_404), .B1(n_454), .B2(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g419 ( .A(n_318), .Y(n_419) );
AND2x2_ASAP7_75t_L g343 ( .A(n_319), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g408 ( .A(n_319), .Y(n_408) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g388 ( .A(n_323), .B(n_324), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_323), .B(n_372), .Y(n_404) );
AND2x2_ASAP7_75t_L g450 ( .A(n_323), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_324), .B(n_428), .Y(n_465) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g377 ( .A(n_325), .Y(n_377) );
INVx1_ASAP7_75t_L g436 ( .A(n_326), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B(n_335), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g398 ( .A(n_330), .B(n_353), .Y(n_398) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_333), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g407 ( .A(n_333), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_336), .B(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_351), .Y(n_337) );
OAI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B(n_346), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_339), .A2(n_406), .B1(n_409), .B2(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI311xp33_ASAP7_75t_L g439 ( .A1(n_341), .A2(n_440), .A3(n_441), .B(n_444), .C(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g367 ( .A(n_344), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_344), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g438 ( .A(n_348), .Y(n_438) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx2_ASAP7_75t_L g444 ( .A(n_354), .Y(n_444) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_358), .Y(n_461) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_385), .Y(n_359) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_365), .C(n_373), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AO21x1_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AO221x1_ASAP7_75t_L g446 ( .A1(n_367), .A2(n_447), .B1(n_450), .B2(n_452), .C(n_453), .Y(n_446) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g445 ( .A(n_372), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B(n_381), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B(n_390), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
AOI221x1_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_398), .B1(n_399), .B2(n_403), .C(n_405), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g423 ( .A(n_394), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AO22x1_ASAP7_75t_L g470 ( .A1(n_398), .A2(n_471), .B1(n_473), .B2(n_476), .Y(n_470) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g447 ( .A(n_401), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_402), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp33_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_446), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_431), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_423), .B(n_425), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .C(n_421), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g456 ( .A(n_418), .Y(n_456) );
AND2x2_ASAP7_75t_L g442 ( .A(n_422), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g452 ( .A(n_428), .B(n_437), .Y(n_452) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_434), .B(n_442), .Y(n_480) );
INVx2_ASAP7_75t_L g472 ( .A(n_437), .Y(n_472) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g475 ( .A(n_443), .Y(n_475) );
AND2x2_ASAP7_75t_L g471 ( .A(n_451), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g483 ( .A(n_451), .Y(n_483) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_462), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_464), .B1(n_466), .B2(n_467), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2x1p5_ASAP7_75t_SL g487 ( .A(n_488), .B(n_741), .Y(n_487) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_489), .B(n_677), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_490), .B(n_598), .C(n_638), .D(n_667), .Y(n_489) );
O2A1O1Ixp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_527), .B(n_534), .C(n_582), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_504), .Y(n_491) );
INVx2_ASAP7_75t_L g530 ( .A(n_492), .Y(n_530) );
AND2x2_ASAP7_75t_L g665 ( .A(n_492), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_492), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_492), .B(n_584), .Y(n_760) );
OR2x2_ASAP7_75t_L g796 ( .A(n_492), .B(n_712), .Y(n_796) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g693 ( .A(n_493), .B(n_505), .Y(n_693) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_493), .B(n_532), .Y(n_719) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g654 ( .A(n_494), .Y(n_654) );
AND2x2_ASAP7_75t_L g592 ( .A(n_504), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_504), .B(n_622), .Y(n_637) );
AND2x2_ASAP7_75t_L g645 ( .A(n_504), .B(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_504), .Y(n_668) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_518), .Y(n_504) );
INVx1_ASAP7_75t_L g532 ( .A(n_505), .Y(n_532) );
INVx1_ASAP7_75t_L g584 ( .A(n_505), .Y(n_584) );
AND2x2_ASAP7_75t_L g655 ( .A(n_505), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g716 ( .A(n_505), .B(n_623), .Y(n_716) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g533 ( .A(n_518), .Y(n_533) );
AND2x2_ASAP7_75t_L g585 ( .A(n_518), .B(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_518), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_518), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g699 ( .A(n_518), .B(n_654), .Y(n_699) );
OR2x2_ASAP7_75t_L g712 ( .A(n_518), .B(n_621), .Y(n_712) );
OR2x2_ASAP7_75t_L g722 ( .A(n_518), .B(n_586), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_523), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g548 ( .A(n_524), .Y(n_548) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_530), .B(n_738), .Y(n_784) );
INVx1_ASAP7_75t_L g640 ( .A(n_531), .Y(n_640) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g724 ( .A(n_533), .B(n_586), .Y(n_724) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_558), .Y(n_534) );
AND2x2_ASAP7_75t_L g596 ( .A(n_535), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g659 ( .A(n_535), .Y(n_659) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_545), .Y(n_535) );
BUFx2_ASAP7_75t_L g766 ( .A(n_536), .Y(n_766) );
AND2x2_ASAP7_75t_L g604 ( .A(n_545), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g590 ( .A(n_546), .B(n_572), .Y(n_590) );
INVx2_ASAP7_75t_L g616 ( .A(n_546), .Y(n_616) );
AOI21x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_549), .B(n_557), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
AND2x2_ASAP7_75t_L g763 ( .A(n_558), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_571), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx4_ASAP7_75t_L g589 ( .A(n_560), .Y(n_589) );
BUFx2_ASAP7_75t_L g597 ( .A(n_560), .Y(n_597) );
OR2x2_ASAP7_75t_L g601 ( .A(n_560), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g662 ( .A(n_560), .B(n_605), .Y(n_662) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B(n_570), .Y(n_562) );
INVx1_ASAP7_75t_L g649 ( .A(n_571), .Y(n_649) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_571), .Y(n_663) );
INVx2_ASAP7_75t_L g688 ( .A(n_571), .Y(n_688) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g602 ( .A(n_572), .Y(n_602) );
OAI21x1_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B(n_581), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B1(n_591), .B2(n_595), .Y(n_582) );
INVx1_ASAP7_75t_L g673 ( .A(n_583), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g684 ( .A(n_584), .Y(n_684) );
AND2x2_ASAP7_75t_L g701 ( .A(n_585), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_585), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g594 ( .A(n_586), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_587), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_588), .B(n_604), .Y(n_696) );
AND2x2_ASAP7_75t_L g704 ( .A(n_588), .B(n_670), .Y(n_704) );
AND2x2_ASAP7_75t_L g780 ( .A(n_588), .B(n_727), .Y(n_780) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g614 ( .A(n_589), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g636 ( .A(n_589), .B(n_605), .Y(n_636) );
OR2x2_ASAP7_75t_L g648 ( .A(n_589), .B(n_649), .Y(n_648) );
NAND2x1_ASAP7_75t_L g682 ( .A(n_589), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g687 ( .A(n_589), .Y(n_687) );
INVx2_ASAP7_75t_L g681 ( .A(n_590), .Y(n_681) );
AND2x2_ASAP7_75t_L g707 ( .A(n_590), .B(n_671), .Y(n_707) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_593), .Y(n_643) );
INVx1_ASAP7_75t_L g710 ( .A(n_593), .Y(n_710) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g694 ( .A(n_594), .B(n_623), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_595), .A2(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g767 ( .A(n_597), .B(n_707), .Y(n_767) );
INVx1_ASAP7_75t_L g803 ( .A(n_597), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_607), .B(n_611), .Y(n_598) );
AOI322xp5_ASAP7_75t_L g751 ( .A1(n_599), .A2(n_647), .A3(n_752), .B1(n_753), .B2(n_754), .C1(n_755), .C2(n_758), .Y(n_751) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_601), .B(n_603), .C(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g617 ( .A(n_602), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g747 ( .A(n_602), .B(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_602), .Y(n_799) );
OR2x2_ASAP7_75t_L g695 ( .A(n_603), .B(n_648), .Y(n_695) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g683 ( .A(n_605), .Y(n_683) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g618 ( .A(n_606), .Y(n_618) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_608), .Y(n_744) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g715 ( .A(n_609), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g778 ( .A(n_610), .B(n_738), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_619), .B(n_634), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_613), .B(n_792), .Y(n_791) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
AND2x2_ASAP7_75t_L g670 ( .A(n_615), .B(n_671), .Y(n_670) );
AND3x2_ASAP7_75t_L g714 ( .A(n_615), .B(n_617), .C(n_687), .Y(n_714) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g676 ( .A(n_616), .Y(n_676) );
AND2x2_ASAP7_75t_L g727 ( .A(n_616), .B(n_688), .Y(n_727) );
INVx2_ASAP7_75t_L g750 ( .A(n_616), .Y(n_750) );
AND2x2_ASAP7_75t_L g754 ( .A(n_617), .B(n_750), .Y(n_754) );
INVx2_ASAP7_75t_L g671 ( .A(n_618), .Y(n_671) );
OR2x2_ASAP7_75t_L g805 ( .A(n_618), .B(n_688), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_619), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g757 ( .A(n_620), .Y(n_757) );
AND2x2_ASAP7_75t_L g666 ( .A(n_621), .B(n_656), .Y(n_666) );
AND2x2_ASAP7_75t_L g702 ( .A(n_621), .B(n_623), .Y(n_702) );
AND2x2_ASAP7_75t_L g698 ( .A(n_622), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_622), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g770 ( .A(n_622), .Y(n_770) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g641 ( .A(n_623), .Y(n_641) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_623), .Y(n_646) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_623), .Y(n_692) );
INVx1_ASAP7_75t_L g738 ( .A(n_623), .Y(n_738) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_647), .B(n_650), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .A3(n_642), .B(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g721 ( .A(n_641), .Y(n_721) );
OAI32xp33_ASAP7_75t_L g679 ( .A1(n_642), .A2(n_651), .A3(n_680), .B1(n_684), .B2(n_685), .Y(n_679) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g672 ( .A(n_648), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_657), .B1(n_660), .B2(n_664), .Y(n_650) );
OAI22xp33_ASAP7_75t_SL g735 ( .A1(n_651), .A2(n_696), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx2_ASAP7_75t_L g793 ( .A(n_653), .Y(n_793) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g748 ( .A(n_656), .Y(n_748) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g674 ( .A(n_662), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g749 ( .A(n_662), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g800 ( .A(n_662), .Y(n_800) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g740 ( .A(n_666), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_673), .B2(n_674), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_669), .B(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
AND2x2_ASAP7_75t_L g726 ( .A(n_671), .B(n_687), .Y(n_726) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_674), .A2(n_732), .B(n_735), .C(n_739), .Y(n_731) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_676), .Y(n_789) );
INVx1_ASAP7_75t_L g806 ( .A(n_676), .Y(n_806) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_700), .C(n_713), .D(n_731), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_689), .Y(n_678) );
OR2x6_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_683), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g788 ( .A(n_686), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_689) );
NOR2xp33_ASAP7_75t_SL g690 ( .A(n_691), .B(n_694), .Y(n_690) );
BUFx2_ASAP7_75t_L g703 ( .A(n_691), .Y(n_703) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_697), .B(n_783), .Y(n_782) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g752 ( .A(n_699), .B(n_738), .Y(n_752) );
O2A1O1Ixp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_704), .C(n_705), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_702), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g762 ( .A(n_709), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_717), .B2(n_725), .C(n_728), .Y(n_713) );
AND2x2_ASAP7_75t_L g792 ( .A(n_716), .B(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .C(n_723), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_721), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_721), .B(n_757), .Y(n_787) );
INVx1_ASAP7_75t_L g730 ( .A(n_722), .Y(n_730) );
INVx1_ASAP7_75t_L g734 ( .A(n_722), .Y(n_734) );
AND2x2_ASAP7_75t_L g775 ( .A(n_724), .B(n_764), .Y(n_775) );
NAND2xp33_ASAP7_75t_SL g776 ( .A(n_724), .B(n_746), .Y(n_776) );
AND2x4_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g736 ( .A(n_727), .Y(n_736) );
NOR3x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_771), .C(n_790), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_751), .C(n_761), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g764 ( .A(n_748), .Y(n_764) );
INVx2_ASAP7_75t_L g753 ( .A(n_750), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_752), .A2(n_795), .B1(n_802), .B2(n_842), .Y(n_801) );
O2A1O1Ixp5_ASAP7_75t_L g773 ( .A1(n_753), .A2(n_765), .B(n_774), .C(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AO21x1_ASAP7_75t_L g777 ( .A1(n_756), .A2(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g769 ( .A(n_760), .B(n_770), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_765), .B1(n_767), .B2(n_768), .Y(n_761) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND4xp75_ASAP7_75t_L g771 ( .A(n_772), .B(n_777), .C(n_781), .D(n_785), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .C(n_801), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OR2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
AND2x4_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
NOR2x1p5_ASAP7_75t_SL g804 ( .A(n_805), .B(n_806), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx6_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx10_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_819), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_825), .B(n_829), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx4_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NOR2x1p5_ASAP7_75t_L g835 ( .A(n_823), .B(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_824), .B(n_837), .Y(n_836) );
INVxp33_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
BUFx6f_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
CKINVDCx11_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
INVx6_ASAP7_75t_L g840 ( .A(n_832), .Y(n_840) );
NAND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_834), .Y(n_833) );
INVx5_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
endmodule