module fake_jpeg_22391_n_59 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.C(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_0),
.B(n_2),
.Y(n_36)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_4),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_31),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_30),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_32),
.B1(n_5),
.B2(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_7),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_40),
.B1(n_44),
.B2(n_10),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_51)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_13),
.C(n_15),
.D(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_17),
.B(n_18),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_19),
.C(n_20),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_21),
.Y(n_59)
);


endmodule