module fake_jpeg_23379_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_20),
.Y(n_52)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_20),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_29),
.B1(n_20),
.B2(n_40),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_21),
.B1(n_25),
.B2(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_43),
.B1(n_40),
.B2(n_44),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_28),
.B1(n_23),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_63),
.B(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_65),
.Y(n_105)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_68),
.B1(n_79),
.B2(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_81),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_93),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_87),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_30),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_27),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_35),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_52),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_44),
.B1(n_38),
.B2(n_43),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_58),
.C(n_61),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_43),
.CI(n_38),
.CON(n_92),
.SN(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_42),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_25),
.B1(n_27),
.B2(n_44),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_99),
.B1(n_44),
.B2(n_25),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_35),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_42),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_98),
.Y(n_121)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_35),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_109),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_126),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_128),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_50),
.B1(n_43),
.B2(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_123),
.C(n_90),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_43),
.C(n_38),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_96),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_62),
.C(n_71),
.Y(n_136)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_93),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_135),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_142),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_72),
.B1(n_65),
.B2(n_101),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_140),
.B1(n_148),
.B2(n_127),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_99),
.B1(n_67),
.B2(n_79),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_149),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_62),
.C(n_71),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_150),
.B(n_151),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_81),
.B1(n_70),
.B2(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_73),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_108),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_80),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_121),
.B1(n_128),
.B2(n_104),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_110),
.B(n_76),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_77),
.C(n_43),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_42),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_92),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_78),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_113),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_31),
.B(n_115),
.C(n_130),
.Y(n_180)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_180),
.B1(n_146),
.B2(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_116),
.B(n_126),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_192),
.B(n_133),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_125),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_133),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_121),
.B1(n_120),
.B2(n_104),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_182),
.B1(n_183),
.B2(n_141),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_189),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_113),
.B1(n_115),
.B2(n_118),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_103),
.B1(n_112),
.B2(n_109),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_135),
.C(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_42),
.B(n_31),
.Y(n_192)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_209),
.C(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_203),
.B(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_217),
.B1(n_221),
.B2(n_219),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_152),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_133),
.B1(n_134),
.B2(n_128),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_183),
.B1(n_192),
.B2(n_180),
.Y(n_224)
);

OA21x2_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_41),
.B(n_24),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_216),
.B(n_219),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_122),
.C(n_41),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_26),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_26),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_122),
.C(n_41),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_41),
.C(n_102),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.C(n_218),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_174),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_0),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_31),
.B1(n_35),
.B2(n_24),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_41),
.C(n_26),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_26),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_179),
.B1(n_175),
.B2(n_180),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_224),
.B1(n_226),
.B2(n_228),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_178),
.B1(n_190),
.B2(n_187),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_227),
.B1(n_243),
.B2(n_24),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_220),
.A2(n_180),
.B1(n_164),
.B2(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_189),
.B1(n_163),
.B2(n_162),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_173),
.B1(n_182),
.B2(n_31),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_199),
.B1(n_213),
.B2(n_193),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_236),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_9),
.B1(n_10),
.B2(n_16),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_212),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_198),
.B1(n_195),
.B2(n_196),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_207),
.B(n_211),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_230),
.B(n_10),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_260),
.B1(n_261),
.B2(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_214),
.C(n_215),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_252),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_253),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_209),
.C(n_218),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_216),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_216),
.C(n_217),
.Y(n_257)
);

BUFx12f_ASAP7_75t_SL g258 ( 
.A(n_233),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_7),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_6),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_267),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_239),
.B(n_224),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_6),
.B(n_15),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_254),
.B(n_234),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_277),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_237),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_275),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_241),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_226),
.B1(n_239),
.B2(n_222),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_242),
.B1(n_230),
.B2(n_2),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_279),
.B(n_250),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_255),
.C(n_251),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_270),
.C(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_248),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_41),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_284),
.Y(n_304)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_291),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_5),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_279),
.B(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_304),
.A3(n_300),
.B1(n_292),
.B2(n_301),
.C1(n_11),
.C2(n_14),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_285),
.C(n_266),
.Y(n_305)
);

AOI332xp33_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_306),
.A3(n_307),
.B1(n_296),
.B2(n_11),
.B3(n_14),
.C1(n_10),
.C2(n_5),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_266),
.C(n_6),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_41),
.B(n_5),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_1),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_312),
.B1(n_314),
.B2(n_1),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_3),
.B(n_4),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_301),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_4),
.C(n_24),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_SL g318 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_314),
.Y(n_320)
);


endmodule