module fake_jpeg_21620_n_62 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_12),
.C(n_9),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_11),
.B1(n_29),
.B2(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_8),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_1),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_12),
.B1(n_10),
.B2(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_37),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_12),
.B(n_2),
.C(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.C(n_34),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_1),
.C(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_12),
.B1(n_2),
.B2(n_4),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_34),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_48),
.C(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_40),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_44),
.B1(n_38),
.B2(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_51),
.C(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_57),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_6),
.C(n_7),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_6),
.Y(n_62)
);


endmodule