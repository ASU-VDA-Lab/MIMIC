module fake_jpeg_15579_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_23),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_0),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_3),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_4),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_56),
.B(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_58),
.C(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

AOI22x1_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_44),
.B1(n_25),
.B2(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_65),
.B1(n_45),
.B2(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_39),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_65),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_70),
.B1(n_69),
.B2(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_70),
.B(n_62),
.Y(n_80)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_76),
.B1(n_47),
.B2(n_69),
.Y(n_79)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_82),
.B(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_82),
.B(n_76),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.C(n_44),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_26),
.C(n_19),
.Y(n_91)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_40),
.B(n_72),
.Y(n_90)
);


endmodule