module real_jpeg_10338_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_335, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_335;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_55),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_47),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_47),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_3),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_33),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_33),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_37),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_3),
.A2(n_30),
.B(n_34),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_113),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_4),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_10),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_93),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_93),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_93),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_11),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_129),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_129),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_100),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_100),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_100),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_13),
.A2(n_24),
.B1(n_63),
.B2(n_64),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_13),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_14),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_57),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_16),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_88),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_88),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_88),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_17),
.A2(n_63),
.B1(n_64),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_17),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_17),
.A2(n_47),
.B1(n_48),
.B2(n_148),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_148),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_148),
.Y(n_280)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_75),
.CON(n_18),
.SN(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_23),
.A2(n_27),
.B1(n_37),
.B2(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_29),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_25),
.A2(n_29),
.B(n_113),
.C(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_27),
.A2(n_37),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_28),
.A2(n_32),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_28),
.A2(n_32),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_28),
.A2(n_32),
.B1(n_211),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_28),
.A2(n_32),
.B1(n_236),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_28),
.A2(n_32),
.B1(n_254),
.B2(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_28),
.A2(n_32),
.B1(n_54),
.B2(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_44),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_67),
.C(n_69),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_39),
.A2(n_40),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_52),
.C(n_58),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_41),
.A2(n_42),
.B1(n_58),
.B2(n_307),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_43),
.A2(n_46),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_43),
.A2(n_46),
.B1(n_139),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_43),
.A2(n_46),
.B1(n_156),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_43),
.A2(n_46),
.B1(n_196),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_43),
.A2(n_46),
.B1(n_207),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_43),
.A2(n_46),
.B1(n_233),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_43),
.A2(n_46),
.B1(n_50),
.B2(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_45),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_46),
.B(n_113),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_47),
.B(n_49),
.Y(n_143)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_48),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_52),
.A2(n_53),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_58),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_58),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_66),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_62),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_59),
.A2(n_62),
.B1(n_99),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_62),
.B1(n_126),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_59),
.A2(n_62),
.B1(n_135),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_59),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_59),
.A2(n_62),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_59),
.A2(n_62),
.B1(n_219),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_59),
.A2(n_62),
.B1(n_228),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_60),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_62),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_62),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_63),
.B(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_66),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_67),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_71),
.A2(n_72),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_325),
.B(n_331),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_298),
.A3(n_318),
.B1(n_323),
.B2(n_324),
.C(n_334),
.Y(n_76)
);

AOI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_244),
.A3(n_286),
.B1(n_292),
.B2(n_297),
.C(n_335),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_201),
.C(n_240),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_171),
.B(n_200),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_150),
.B(n_170),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_131),
.B(n_149),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_120),
.B(n_130),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_106),
.B(n_119),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_85),
.B(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_89),
.A2(n_90),
.B1(n_147),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_110),
.B1(n_111),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_105),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_114),
.B(n_118),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_111),
.B1(n_128),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_110),
.A2(n_111),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_110),
.A2(n_111),
.B1(n_182),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_110),
.A2(n_111),
.B1(n_216),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_110),
.A2(n_111),
.B(n_226),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_125),
.C(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.CI(n_140),
.CON(n_133),
.SN(n_133)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_145),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_163),
.B2(n_164),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_166),
.C(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_162),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_160),
.C(n_162),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_165),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_166),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_167),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_172),
.B(n_173),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_186),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_175),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_185),
.C(n_186),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_180),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_194),
.B2(n_195),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_194),
.C(n_197),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_191),
.A2(n_193),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_199),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_202),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_221),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_203),
.B(n_221),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.C(n_220),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_213),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_212),
.C(n_213),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_217),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_238),
.B2(n_239),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_229),
.C(n_239),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_227),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_234),
.C(n_237),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_242),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_263),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_245),
.B(n_263),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_256),
.C(n_262),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_246),
.A2(n_247),
.B1(n_256),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_252),
.C(n_255),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_251),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_256),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_258),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_257),
.A2(n_279),
.B(n_282),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_259),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_259),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_284),
.B2(n_285),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_276),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_276),
.C(n_285),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_271),
.B(n_274),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_271),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_273),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_274),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_274),
.A2(n_300),
.B1(n_309),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_282),
.B2(n_283),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_279),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_311),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_309),
.C(n_310),
.Y(n_299)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_301),
.A2(n_302),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_307),
.C(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_313),
.C(n_317),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_305),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_330),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_327),
.Y(n_329)
);


endmodule