module real_jpeg_6874_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_1),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_1),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_1),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_2),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_2),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_2),
.B(n_115),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_2),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_3),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_3),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_5),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_5),
.B(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_5),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_5),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_7),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_7),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_7),
.B(n_53),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_11),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_11),
.B(n_166),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_13),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_13),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_14),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_14),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_14),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_15),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_15),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_15),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_195),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_193),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_153),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_19),
.B(n_153),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.C(n_137),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_20),
.B(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_65),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_21),
.B(n_66),
.C(n_80),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_56),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_22),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_32),
.B2(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_25),
.B(n_32),
.C(n_37),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_45),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_26),
.B(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_30),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_30),
.Y(n_247)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_31),
.Y(n_218)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_34),
.Y(n_163)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_35),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_41),
.B(n_104),
.Y(n_294)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_43),
.A2(n_56),
.B1(n_57),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.C(n_50),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_44),
.A2(n_50),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_44),
.Y(n_208)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_46),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_47),
.B(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_58),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_58),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_176),
.Y(n_223)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_80),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_68),
.B(n_74),
.C(n_78),
.Y(n_192)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_71),
.Y(n_222)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_75),
.B(n_123),
.Y(n_242)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_76),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_88),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_81),
.B(n_89),
.C(n_95),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_96),
.B(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_101),
.B(n_137),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_118),
.C(n_120),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_102),
.A2(n_118),
.B1(n_119),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_107),
.C(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_104),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B1(n_112),
.B2(n_117),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_120),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_132),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_121),
.A2(n_122),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_324)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_131),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_131),
.Y(n_298)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_152),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_140),
.C(n_152),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_148),
.C(n_151),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_146),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_179),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_170),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_177),
.B2(n_178),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_173),
.A2(n_174),
.B1(n_234),
.B2(n_235),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_174),
.B(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_192),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_227),
.B(n_332),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_198),
.B(n_200),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.C(n_224),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_201),
.A2(n_202),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_205),
.B(n_224),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_223),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_206),
.B(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_210),
.B(n_223),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.C(n_219),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_212),
.B1(n_219),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_220),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_326),
.B(n_331),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_313),
.B(n_325),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_273),
.B(n_312),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_256),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_231),
.B(n_256),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_232),
.B(n_244),
.C(n_253),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_233),
.B(n_239),
.C(n_242),
.Y(n_321)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_258),
.Y(n_257)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.C(n_272),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_259),
.A2(n_260),
.B1(n_272),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_262),
.B1(n_268),
.B2(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_306),
.B(n_311),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_292),
.B(n_305),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_283),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_280),
.C(n_282),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_285),
.B1(n_289),
.B2(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_299),
.B(n_304),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_303),
.Y(n_304)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_315),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_321),
.C(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule