module fake_jpeg_12511_n_515 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_13),
.B(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_60),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_78),
.Y(n_125)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_67),
.B(n_82),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_68),
.Y(n_187)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_1),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_81),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_90),
.Y(n_144)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_96),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_2),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_106),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_21),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_111),
.Y(n_127)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_109),
.B(n_110),
.Y(n_197)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_34),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_115),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

NAND2x1_ASAP7_75t_SL g114 ( 
.A(n_20),
.B(n_3),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_114),
.A2(n_4),
.B(n_5),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_4),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_119),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_25),
.B(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_123),
.Y(n_138)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_41),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_122),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_46),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_85),
.A2(n_47),
.B1(n_30),
.B2(n_24),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_136),
.A2(n_150),
.B1(n_170),
.B2(n_175),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_98),
.B1(n_107),
.B2(n_109),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_140),
.A2(n_169),
.B(n_133),
.C(n_136),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_30),
.C(n_56),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_147),
.B(n_149),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_66),
.A2(n_22),
.B1(n_40),
.B2(n_32),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_148),
.A2(n_154),
.B1(n_174),
.B2(n_193),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_29),
.C(n_56),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_47),
.B1(n_40),
.B2(n_32),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_76),
.A2(n_22),
.B1(n_40),
.B2(n_32),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_92),
.B(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_8),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_58),
.B1(n_22),
.B2(n_26),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_169),
.A2(n_150),
.B1(n_175),
.B2(n_179),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_97),
.A2(n_41),
.B1(n_43),
.B2(n_20),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_171),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_177),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_28),
.B1(n_43),
.B2(n_38),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_80),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_70),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_72),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_179),
.A2(n_199),
.B1(n_192),
.B2(n_135),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_94),
.B(n_55),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_185),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_140),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_79),
.B(n_55),
.Y(n_185)
);

OA22x2_ASAP7_75t_SL g189 ( 
.A1(n_61),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_10),
.B(n_12),
.C(n_14),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_64),
.B(n_37),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_191),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_65),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_68),
.B(n_6),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_195),
.B(n_198),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_75),
.B(n_8),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_113),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_202),
.B(n_206),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_204),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_127),
.A2(n_86),
.B1(n_93),
.B2(n_89),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_205),
.A2(n_211),
.B1(n_222),
.B2(n_226),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_207),
.A2(n_241),
.A3(n_251),
.B1(n_218),
.B2(n_229),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_209),
.B(n_210),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_128),
.A2(n_83),
.B1(n_87),
.B2(n_95),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_10),
.B(n_12),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_212),
.A2(n_214),
.B(n_225),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_213),
.B(n_223),
.Y(n_280)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_145),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_216),
.B(n_219),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_139),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_217),
.B(n_227),
.C(n_203),
.Y(n_315)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_189),
.B1(n_167),
.B2(n_131),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_138),
.A2(n_189),
.B1(n_199),
.B2(n_134),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_142),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_140),
.A2(n_188),
.B1(n_161),
.B2(n_130),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_161),
.A2(n_124),
.B1(n_126),
.B2(n_143),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_132),
.B1(n_196),
.B2(n_156),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_233),
.A2(n_253),
.B1(n_217),
.B2(n_244),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_126),
.A2(n_135),
.B1(n_196),
.B2(n_129),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_234),
.A2(n_236),
.B1(n_246),
.B2(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_137),
.B(n_181),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_235),
.B(n_237),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_129),
.A2(n_159),
.B1(n_153),
.B2(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_152),
.B(n_125),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_132),
.A2(n_200),
.B1(n_153),
.B2(n_164),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_239),
.A2(n_254),
.B1(n_267),
.B2(n_255),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_172),
.A2(n_194),
.B1(n_187),
.B2(n_162),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_249),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_157),
.A2(n_171),
.B(n_183),
.C(n_166),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_172),
.A2(n_194),
.B1(n_187),
.B2(n_162),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_164),
.A2(n_201),
.B1(n_176),
.B2(n_186),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_129),
.A2(n_159),
.B1(n_144),
.B2(n_166),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_258),
.Y(n_284)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_186),
.A2(n_163),
.B1(n_144),
.B2(n_159),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_157),
.Y(n_252)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_189),
.A2(n_136),
.B1(n_150),
.B2(n_140),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_189),
.A2(n_107),
.B1(n_109),
.B2(n_98),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_257),
.Y(n_318)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

BUFx24_ASAP7_75t_L g295 ( 
.A(n_257),
.Y(n_295)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_163),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_182),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_264),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_127),
.B(n_128),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_227),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_263),
.A2(n_268),
.B1(n_249),
.B2(n_252),
.Y(n_288)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_156),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_146),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_266),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_182),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_189),
.A2(n_107),
.B1(n_109),
.B2(n_98),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_140),
.A2(n_47),
.B1(n_96),
.B2(n_85),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_235),
.B(n_237),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_291),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_273),
.A2(n_290),
.B1(n_294),
.B2(n_307),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_222),
.A2(n_216),
.B1(n_219),
.B2(n_213),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_209),
.B1(n_225),
.B2(n_226),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_315),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_216),
.A2(n_205),
.B1(n_211),
.B2(n_261),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_217),
.A2(n_240),
.B1(n_243),
.B2(n_206),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_288),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_208),
.A2(n_232),
.B1(n_259),
.B2(n_223),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_260),
.B(n_266),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_202),
.B(n_221),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_292),
.B(n_303),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_232),
.A2(n_207),
.B1(n_242),
.B2(n_212),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_298),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_227),
.A2(n_220),
.B1(n_224),
.B2(n_215),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_300),
.A2(n_279),
.B1(n_287),
.B2(n_293),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_299),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_275),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_231),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_245),
.B(n_248),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_304),
.B(n_308),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_203),
.A2(n_238),
.B1(n_262),
.B2(n_264),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_204),
.B(n_247),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_252),
.B(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_311),
.B(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_263),
.B(n_250),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_238),
.B(n_262),
.C(n_269),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_274),
.C(n_314),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_318),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_276),
.A2(n_306),
.B1(n_294),
.B2(n_290),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_319),
.A2(n_348),
.B(n_352),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_281),
.A2(n_258),
.B1(n_314),
.B2(n_307),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_310),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_324),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_325),
.B(n_328),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_331),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_302),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_306),
.A2(n_273),
.B1(n_278),
.B2(n_280),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_329),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_335),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_298),
.Y(n_335)
);

BUFx12f_ASAP7_75t_SL g336 ( 
.A(n_295),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_336),
.B(n_337),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_270),
.Y(n_337)
);

NAND2x1_ASAP7_75t_SL g338 ( 
.A(n_315),
.B(n_306),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_338),
.A2(n_340),
.B(n_297),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_275),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_343),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_296),
.A2(n_278),
.B(n_280),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_292),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_282),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

OR2x4_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_282),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_347),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_285),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_303),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_350),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_271),
.A2(n_286),
.B1(n_296),
.B2(n_279),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_351),
.A2(n_271),
.B1(n_316),
.B2(n_284),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_285),
.B(n_318),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_358),
.B1(n_330),
.B2(n_344),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_351),
.A2(n_313),
.B1(n_283),
.B2(n_284),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_343),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_SL g407 ( 
.A(n_359),
.B(n_361),
.C(n_376),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_335),
.A2(n_311),
.B(n_318),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_360),
.A2(n_381),
.B(n_349),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_322),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_272),
.C(n_309),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_365),
.C(n_353),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_272),
.C(n_309),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_339),
.B(n_328),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_367),
.A2(n_338),
.B(n_319),
.Y(n_403)
);

INVx13_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_370),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_332),
.A2(n_305),
.B(n_312),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_322),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_297),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_379),
.B(n_321),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_295),
.B(n_312),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_347),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_384),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_390),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_348),
.Y(n_384)
);

FAx1_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_346),
.CI(n_340),
.CON(n_385),
.SN(n_385)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_385),
.A2(n_388),
.B(n_400),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_364),
.A2(n_362),
.B1(n_326),
.B2(n_345),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_393),
.B1(n_399),
.B2(n_362),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_368),
.B(n_337),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_394),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_403),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_330),
.B1(n_326),
.B2(n_325),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_368),
.B(n_333),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_328),
.C(n_334),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_404),
.C(n_405),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_356),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_401),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_331),
.B1(n_341),
.B2(n_348),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_375),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_369),
.B(n_333),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_359),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_352),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_342),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_341),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_406),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_323),
.Y(n_432)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_412),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_416),
.A2(n_421),
.B(n_426),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_381),
.Y(n_417)
);

AO21x1_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_432),
.B(n_386),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_420),
.B(n_429),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_400),
.A2(n_377),
.B(n_355),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_374),
.Y(n_423)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_371),
.C(n_363),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_427),
.C(n_431),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_387),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_428),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_403),
.A2(n_366),
.B(n_367),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_371),
.C(n_365),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_354),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_394),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_363),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_354),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_433),
.B(n_380),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_430),
.A2(n_406),
.B1(n_389),
.B2(n_399),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_434),
.A2(n_448),
.B1(n_451),
.B2(n_454),
.Y(n_455)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_436),
.Y(n_459)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_438),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_365),
.C(n_404),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_440),
.C(n_445),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_366),
.C(n_386),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_395),
.C(n_402),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_392),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_393),
.C(n_360),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_410),
.A2(n_419),
.B1(n_428),
.B2(n_418),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_413),
.A2(n_401),
.B1(n_388),
.B2(n_380),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_452),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_416),
.A2(n_369),
.B(n_385),
.C(n_373),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_433),
.B(n_378),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_415),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_410),
.A2(n_357),
.B1(n_385),
.B2(n_381),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_447),
.A2(n_418),
.B1(n_419),
.B2(n_413),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_456),
.A2(n_461),
.B1(n_434),
.B2(n_454),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_437),
.A2(n_425),
.B(n_421),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_457),
.A2(n_437),
.B(n_438),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_439),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_462),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_447),
.A2(n_420),
.B1(n_415),
.B2(n_426),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_431),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_422),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_469),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_467),
.C(n_453),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_432),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_423),
.C(n_414),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_468),
.B(n_449),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_412),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_448),
.Y(n_470)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_472),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_468),
.B(n_445),
.C(n_449),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_475),
.Y(n_487)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_466),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_476),
.A2(n_455),
.B1(n_457),
.B2(n_452),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_478),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_458),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_446),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_479),
.B(n_481),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_463),
.B(n_441),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_455),
.C(n_465),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_475),
.A2(n_357),
.B1(n_441),
.B2(n_451),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_483),
.A2(n_473),
.B1(n_470),
.B2(n_471),
.Y(n_494)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_488),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_465),
.C(n_460),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_474),
.C(n_480),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_490),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_476),
.A2(n_443),
.B1(n_378),
.B2(n_411),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_492),
.A2(n_358),
.B1(n_417),
.B2(n_396),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_495),
.Y(n_501)
);

NAND4xp25_ASAP7_75t_SL g496 ( 
.A(n_487),
.B(n_479),
.C(n_295),
.D(n_370),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_496),
.A2(n_417),
.B(n_370),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_480),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_499),
.C(n_488),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_474),
.C(n_462),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_500),
.A2(n_483),
.B1(n_385),
.B2(n_485),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_493),
.A2(n_491),
.B1(n_490),
.B2(n_486),
.Y(n_502)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_414),
.B(n_352),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_493),
.A2(n_498),
.B(n_414),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_504),
.A2(n_469),
.B(n_496),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_506),
.C(n_499),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_509),
.C(n_505),
.Y(n_511)
);

AO21x1_ASAP7_75t_L g512 ( 
.A1(n_510),
.A2(n_501),
.B(n_504),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_512),
.C(n_508),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_502),
.Y(n_515)
);


endmodule