module real_jpeg_6649_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_0),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_0),
.Y(n_237)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_3),
.A2(n_167),
.B1(n_170),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_121),
.B1(n_172),
.B2(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_5),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_5),
.A2(n_97),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_5),
.A2(n_97),
.B1(n_139),
.B2(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_6),
.Y(n_161)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_6),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_6),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_7),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_8),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_11),
.A2(n_92),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_11),
.A2(n_92),
.B1(n_125),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_11),
.A2(n_92),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_12),
.A2(n_47),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_106),
.C(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_12),
.B(n_77),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_12),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_104),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_12),
.B(n_330),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_13),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_13),
.A2(n_122),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_14),
.Y(n_116)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_14),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_15),
.A2(n_53),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_15),
.A2(n_53),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_15),
.A2(n_53),
.B1(n_162),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_245),
.B1(n_246),
.B2(n_365),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_18),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_244),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_205),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_20),
.B(n_205),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_141),
.C(n_184),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_21),
.B(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_140),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_22),
.B(n_59),
.C(n_102),
.Y(n_225)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B(n_50),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_24),
.B(n_52),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_34),
.B(n_47),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_34)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_35),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_37),
.Y(n_190)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_38),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_39),
.A2(n_48),
.A3(n_145),
.B1(n_149),
.B2(n_151),
.Y(n_144)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_43),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_48),
.Y(n_44)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_47),
.A2(n_159),
.B(n_271),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_47),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_57),
.Y(n_238)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_102),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_86),
.B1(n_93),
.B2(n_94),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_60),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_77),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_64),
.Y(n_340)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_66),
.Y(n_346)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_76),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_76),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_76),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_77),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_81),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_81),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_83),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_83),
.Y(n_261)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_86),
.A2(n_93),
.B(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_93),
.B(n_188),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_94),
.Y(n_242)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_117),
.B(n_123),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_103),
.A2(n_117),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_103),
.A2(n_209),
.B1(n_278),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_104),
.B(n_124),
.Y(n_258)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_105),
.A2(n_123),
.B(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_113),
.B2(n_115),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_121),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g338 ( 
.A(n_125),
.Y(n_338)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_128),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_133),
.B1(n_136),
.B2(n_139),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_132),
.Y(n_323)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_141),
.A2(n_142),
.B1(n_184),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_157),
.B2(n_158),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_144),
.B(n_157),
.Y(n_229)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_165),
.B1(n_173),
.B2(n_177),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_159),
.A2(n_266),
.B(n_271),
.Y(n_265)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_166),
.B1(n_196),
.B2(n_202),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_160),
.A2(n_178),
.B1(n_216),
.B2(n_223),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_160),
.B(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_160),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_161),
.Y(n_309)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_169),
.Y(n_274)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_169),
.Y(n_296)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_176),
.Y(n_287)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_176),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.C(n_204),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_185),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_194),
.A2(n_243),
.B(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_195),
.B(n_204),
.Y(n_356)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_196),
.Y(n_334)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_201),
.Y(n_293)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_228),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_209),
.A2(n_253),
.B(n_258),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_209),
.A2(n_258),
.B(n_320),
.Y(n_353)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_240),
.B2(n_241),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_239),
.Y(n_232)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_359),
.B(n_364),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_348),
.B(n_358),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_314),
.B(n_347),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_282),
.B(n_313),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_264),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_264),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_252),
.A2(n_259),
.B1(n_260),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_276),
.C(n_281),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_303),
.B(n_312),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_289),
.B(n_302),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_301),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_301),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_310),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_316),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_332),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_324),
.B2(n_325),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_324),
.C(n_332),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI32xp33_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_337),
.A3(n_338),
.B1(n_339),
.B2(n_341),
.Y(n_336)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_336),
.Y(n_354)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_349),
.B(n_350),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_355),
.B2(n_357),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_354),
.C(n_357),
.Y(n_360)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_360),
.B(n_361),
.Y(n_364)
);


endmodule