module fake_jpeg_30311_n_156 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_15),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_10),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_76),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_89),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_64),
.B1(n_54),
.B2(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_64),
.B1(n_54),
.B2(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_88),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_59),
.B1(n_52),
.B2(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_56),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_60),
.B(n_49),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_98),
.B(n_99),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_76),
.B1(n_63),
.B2(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_56),
.B1(n_48),
.B2(n_2),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_0),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_21),
.C(n_44),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_9),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_105),
.B(n_110),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_3),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_22),
.B(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_3),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_115),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_109),
.A2(n_26),
.B(n_39),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_122),
.B1(n_129),
.B2(n_36),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_4),
.B(n_5),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_7),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_121),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_7),
.B(n_8),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_125),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_92),
.C(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_13),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_32),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_16),
.B1(n_18),
.B2(n_27),
.Y(n_129)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.Y(n_144)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_138),
.C(n_140),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_124),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_128),
.B1(n_113),
.B2(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_131),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_130),
.B(n_133),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_141),
.B(n_115),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_149),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_145),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_150),
.B(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_135),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_123),
.Y(n_156)
);


endmodule