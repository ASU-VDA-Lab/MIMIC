module fake_netlist_1_12592_n_719 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_719, n_722);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_719;
output n_722;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_93), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_32), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_64), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_79), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_83), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_62), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_52), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_86), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_6), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_94), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_10), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_27), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_19), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_67), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_7), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_17), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_69), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_71), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_91), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_99), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_48), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_72), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_6), .Y(n_129) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_59), .B(n_42), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_66), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_47), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_24), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_57), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_44), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_96), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_65), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_102), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_108), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_107), .B(n_0), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_114), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_131), .B(n_0), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_128), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g149 ( .A1(n_110), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_105), .B(n_1), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_119), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_128), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_105), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g156 ( .A1(n_112), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
XOR2x2_ASAP7_75t_L g161 ( .A(n_149), .B(n_4), .Y(n_161) );
AND3x2_ASAP7_75t_L g162 ( .A(n_146), .B(n_129), .C(n_125), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_151), .B(n_127), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_151), .B(n_100), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_150), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_142), .A2(n_158), .B1(n_117), .B2(n_118), .Y(n_174) );
AND3x2_ASAP7_75t_L g175 ( .A(n_146), .B(n_123), .C(n_126), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_151), .B(n_100), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
AOI21x1_ASAP7_75t_L g179 ( .A1(n_140), .A2(n_137), .B(n_132), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_140), .B(n_103), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_141), .B(n_103), .Y(n_181) );
NAND3xp33_ASAP7_75t_L g182 ( .A(n_141), .B(n_133), .C(n_135), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_143), .B(n_104), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_181), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_149), .B1(n_156), .B2(n_147), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_173), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_183), .B(n_143), .Y(n_190) );
NOR2xp33_ASAP7_75t_SL g191 ( .A(n_173), .B(n_104), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_167), .B(n_147), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_165), .B(n_155), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_165), .B(n_155), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_176), .B(n_106), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_180), .B(n_106), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_174), .B(n_109), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_185), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_182), .B(n_109), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_182), .B(n_111), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_172), .A2(n_156), .B1(n_144), .B2(n_153), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_175), .B(n_111), .Y(n_209) );
NAND3xp33_ASAP7_75t_L g210 ( .A(n_172), .B(n_152), .C(n_153), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_152), .B1(n_101), .B2(n_127), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_177), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_179), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_162), .B(n_121), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_179), .B(n_121), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_130), .B(n_124), .C(n_139), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_159), .B(n_124), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_160), .B(n_134), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_161), .B(n_134), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_161), .B(n_136), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_160), .B(n_136), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_213), .A2(n_186), .B(n_184), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_190), .A2(n_184), .B(n_178), .Y(n_225) );
NOR2x1_ASAP7_75t_L g226 ( .A(n_214), .B(n_115), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_204), .A2(n_138), .B1(n_139), .B2(n_120), .Y(n_227) );
AOI21x1_ASAP7_75t_L g228 ( .A1(n_213), .A2(n_178), .B(n_171), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_189), .A2(n_171), .B(n_168), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_187), .B(n_138), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_189), .A2(n_168), .B(n_166), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_192), .A2(n_166), .B(n_164), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_220), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_205), .B(n_5), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_193), .A2(n_128), .B1(n_157), .B2(n_154), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_193), .A2(n_157), .B1(n_154), .B2(n_164), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_195), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_197), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_197), .Y(n_240) );
AOI22x1_ASAP7_75t_L g241 ( .A1(n_215), .A2(n_157), .B1(n_154), .B2(n_163), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_194), .A2(n_157), .B(n_154), .C(n_8), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_203), .B(n_5), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_196), .A2(n_157), .B1(n_154), .B2(n_9), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_192), .A2(n_41), .B(n_95), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_188), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_188), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_191), .B(n_11), .Y(n_248) );
AO32x1_ASAP7_75t_L g249 ( .A1(n_215), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_200), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_200), .A2(n_46), .B(n_92), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_191), .B(n_14), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_199), .B(n_15), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_208), .A2(n_16), .B(n_17), .C(n_18), .Y(n_254) );
CKINVDCx8_ASAP7_75t_R g255 ( .A(n_230), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_253), .A2(n_243), .B(n_250), .C(n_254), .Y(n_256) );
AOI21xp5_ASAP7_75t_SL g257 ( .A1(n_242), .A2(n_217), .B(n_212), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_234), .B(n_220), .Y(n_258) );
AOI21x1_ASAP7_75t_SL g259 ( .A1(n_248), .A2(n_222), .B(n_207), .Y(n_259) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_242), .A2(n_201), .A3(n_212), .B(n_198), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_224), .A2(n_201), .B(n_210), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_233), .Y(n_263) );
BUFx4_ASAP7_75t_SL g264 ( .A(n_239), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_230), .B(n_221), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_238), .A2(n_198), .B1(n_211), .B2(n_206), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_228), .A2(n_216), .B(n_223), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_253), .B(n_208), .Y(n_268) );
OAI21xp33_ASAP7_75t_SL g269 ( .A1(n_235), .A2(n_202), .B(n_219), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_229), .A2(n_216), .B(n_223), .Y(n_270) );
NOR4xp25_ASAP7_75t_L g271 ( .A(n_246), .B(n_210), .C(n_209), .D(n_218), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_244), .A2(n_16), .A3(n_18), .B(n_20), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_225), .A2(n_21), .B(n_22), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_240), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_240), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_226), .B(n_23), .Y(n_276) );
AO32x2_ASAP7_75t_L g277 ( .A1(n_247), .A2(n_25), .A3(n_26), .B1(n_28), .B2(n_29), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_259), .A2(n_241), .B(n_251), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_268), .B(n_252), .Y(n_279) );
NOR2x1_ASAP7_75t_L g280 ( .A(n_257), .B(n_245), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_256), .A2(n_231), .B(n_232), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_269), .A2(n_271), .B(n_266), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
BUFx2_ASAP7_75t_R g286 ( .A(n_255), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_261), .Y(n_287) );
AOI21x1_ASAP7_75t_L g288 ( .A1(n_262), .A2(n_249), .B(n_227), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_260), .B(n_236), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_274), .B(n_237), .Y(n_291) );
INVxp33_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
OR2x6_ASAP7_75t_L g293 ( .A(n_275), .B(n_249), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_270), .A2(n_237), .B(n_236), .Y(n_294) );
OAI21x1_ASAP7_75t_SL g295 ( .A1(n_273), .A2(n_249), .B(n_31), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_259), .A2(n_249), .B(n_33), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_260), .A2(n_30), .B(n_34), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_285), .B(n_260), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_287), .B(n_272), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_285), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_297), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_287), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_282), .A2(n_276), .B(n_277), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_297), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_282), .A2(n_276), .B(n_277), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_279), .B(n_272), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_297), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_278), .A2(n_277), .B(n_272), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_277), .B(n_272), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_295), .A2(n_265), .B(n_36), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_289), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_280), .B(n_265), .Y(n_324) );
AO21x1_ASAP7_75t_SL g325 ( .A1(n_283), .A2(n_35), .B(n_37), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_289), .Y(n_326) );
OR2x6_ASAP7_75t_L g327 ( .A(n_293), .B(n_39), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_279), .A2(n_40), .B(n_43), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_320), .B(n_298), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_311), .B(n_293), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_311), .B(n_320), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_320), .B(n_298), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_322), .B(n_298), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_327), .Y(n_336) );
NOR2x1_ASAP7_75t_SL g337 ( .A(n_327), .B(n_293), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_301), .Y(n_338) );
INVx4_ASAP7_75t_R g339 ( .A(n_304), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_301), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_322), .B(n_298), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_322), .B(n_293), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_327), .B(n_293), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_305), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_326), .B(n_293), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_327), .Y(n_353) );
BUFx4f_ASAP7_75t_L g354 ( .A(n_327), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_303), .Y(n_356) );
OAI222xp33_ASAP7_75t_L g357 ( .A1(n_327), .A2(n_293), .B1(n_290), .B2(n_280), .C1(n_288), .C2(n_291), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_306), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_326), .B(n_292), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_326), .B(n_281), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_308), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_313), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_319), .B(n_281), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_300), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_308), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_319), .A2(n_292), .B1(n_290), .B2(n_291), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_304), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_317), .B(n_281), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_302), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_300), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_302), .B(n_291), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_324), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_323), .B(n_281), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_323), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_375), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_375), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_359), .B(n_324), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_332), .B(n_321), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_359), .B(n_309), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_343), .B(n_321), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_356), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_343), .B(n_314), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_350), .B(n_314), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_329), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_356), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
BUFx4f_ASAP7_75t_L g395 ( .A(n_336), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_332), .B(n_315), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_361), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_350), .B(n_314), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_350), .B(n_340), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_329), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_359), .B(n_307), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
BUFx2_ASAP7_75t_SL g405 ( .A(n_336), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_329), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_338), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_362), .B(n_286), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_354), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_340), .B(n_315), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_354), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_376), .B(n_315), .Y(n_413) );
AND2x4_ASAP7_75t_SL g414 ( .A(n_336), .B(n_291), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_346), .B(n_307), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_376), .B(n_309), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_338), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_337), .A2(n_307), .B1(n_309), .B2(n_318), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_346), .B(n_309), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_336), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_331), .B(n_307), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_367), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_338), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_331), .B(n_307), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_367), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_353), .B(n_328), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_341), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_371), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_337), .B(n_345), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_353), .B(n_328), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
NOR2xp67_ASAP7_75t_L g434 ( .A(n_345), .B(n_288), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_364), .B(n_309), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_333), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_373), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_364), .B(n_360), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_377), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_377), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_365), .B(n_318), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_365), .B(n_318), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_364), .B(n_281), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g444 ( .A(n_345), .B(n_325), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_360), .B(n_325), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_341), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_345), .A2(n_295), .B1(n_294), .B2(n_278), .Y(n_447) );
NOR2x1_ASAP7_75t_SL g448 ( .A(n_378), .B(n_286), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_363), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_360), .B(n_294), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_369), .B(n_45), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_333), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_339), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_345), .B(n_49), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_341), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_438), .B(n_401), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_401), .B(n_344), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_431), .B(n_378), .Y(n_458) );
NOR2xp33_ASAP7_75t_SL g459 ( .A(n_398), .B(n_357), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_438), .B(n_344), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_394), .B(n_373), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_396), .B(n_378), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_380), .B(n_358), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_410), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_381), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_436), .B(n_357), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_439), .B(n_379), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_431), .B(n_379), .Y(n_469) );
NAND2x1_ASAP7_75t_L g470 ( .A(n_398), .B(n_339), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_382), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_384), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_440), .B(n_379), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_388), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_380), .B(n_358), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_389), .B(n_330), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_431), .B(n_374), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_393), .B(n_330), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_399), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_422), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_392), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_423), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_424), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_449), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_427), .Y(n_487) );
AOI211xp5_ASAP7_75t_L g488 ( .A1(n_408), .A2(n_330), .B(n_334), .C(n_335), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_430), .B(n_334), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_421), .B(n_334), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_445), .B(n_335), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_452), .B(n_368), .C(n_374), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_385), .B(n_352), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_392), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_428), .B(n_335), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_445), .B(n_342), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_387), .B(n_342), .Y(n_498) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_402), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_385), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_449), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_402), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_406), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_387), .B(n_355), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_454), .B(n_342), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_383), .B(n_355), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_406), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_407), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_454), .B(n_374), .Y(n_509) );
NAND5xp2_ASAP7_75t_L g510 ( .A(n_444), .B(n_368), .C(n_374), .D(n_53), .E(n_54), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_390), .B(n_374), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_390), .B(n_355), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_421), .B(n_372), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_416), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_391), .B(n_352), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_407), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_417), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_453), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_398), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_426), .B(n_372), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_397), .B(n_352), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_444), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_391), .B(n_351), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_453), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_417), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_397), .B(n_351), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_404), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_444), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_400), .B(n_351), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_400), .B(n_349), .Y(n_530) );
OAI221xp5_ASAP7_75t_SL g531 ( .A1(n_416), .A2(n_368), .B1(n_370), .B2(n_372), .C(n_363), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_425), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_425), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_429), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_420), .B(n_370), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_414), .B(n_349), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_429), .Y(n_537) );
INVx3_ASAP7_75t_SL g538 ( .A(n_414), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_426), .B(n_370), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_446), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_404), .B(n_368), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_446), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_409), .B(n_349), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_455), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_456), .B(n_435), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_524), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_500), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_522), .A2(n_395), .B(n_409), .C(n_412), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_456), .B(n_435), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_469), .B(n_411), .Y(n_550) );
NAND2x2_ASAP7_75t_L g551 ( .A(n_518), .B(n_448), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_466), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_470), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_511), .B(n_411), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_518), .B(n_448), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_462), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
OAI32xp33_ASAP7_75t_L g558 ( .A1(n_522), .A2(n_441), .A3(n_442), .B1(n_432), .B2(n_413), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_514), .B(n_415), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_514), .B(n_415), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_471), .Y(n_561) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_476), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_483), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_538), .Y(n_564) );
NAND5xp2_ASAP7_75t_SL g565 ( .A(n_463), .B(n_447), .C(n_443), .D(n_395), .E(n_405), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_476), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_461), .B(n_413), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_511), .B(n_443), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_472), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_492), .B(n_420), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_539), .B(n_419), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_539), .B(n_386), .Y(n_572) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_510), .B(n_405), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_513), .B(n_403), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_538), .Y(n_575) );
AOI32xp33_ASAP7_75t_L g576 ( .A1(n_459), .A2(n_418), .A3(n_442), .B1(n_441), .B2(n_451), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_491), .B(n_450), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_496), .B(n_434), .Y(n_578) );
NOR2xp33_ASAP7_75t_SL g579 ( .A(n_522), .B(n_395), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_534), .Y(n_580) );
AOI21xp33_ASAP7_75t_SL g581 ( .A1(n_528), .A2(n_455), .B(n_348), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_497), .B(n_363), .Y(n_582) );
OR2x6_ASAP7_75t_L g583 ( .A(n_528), .B(n_348), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_498), .B(n_512), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_474), .Y(n_585) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_481), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_520), .B(n_348), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_481), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_478), .B(n_50), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_458), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_467), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_496), .B(n_51), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_515), .B(n_55), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_528), .A2(n_97), .B(n_58), .C(n_60), .Y(n_595) );
AOI32xp33_ASAP7_75t_L g596 ( .A1(n_527), .A2(n_56), .A3(n_61), .B1(n_73), .B2(n_75), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_468), .B(n_76), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_458), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_464), .B(n_77), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_523), .B(n_78), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_480), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_473), .B(n_80), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_482), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_475), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_458), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_531), .A2(n_81), .B(n_82), .C(n_87), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_484), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_501), .B(n_88), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_485), .Y(n_609) );
NOR2xp33_ASAP7_75t_SL g610 ( .A(n_519), .B(n_89), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_521), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_529), .B(n_90), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_487), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_490), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_457), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_467), .B(n_460), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_465), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_504), .B(n_494), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_576), .A2(n_591), .B(n_616), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_604), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_564), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_552), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_616), .B(n_530), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_615), .B(n_545), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_546), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_557), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_588), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_573), .A2(n_478), .B1(n_488), .B2(n_519), .Y(n_628) );
AOI211xp5_ASAP7_75t_L g629 ( .A1(n_555), .A2(n_493), .B(n_541), .C(n_519), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_549), .B(n_506), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_561), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_546), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_575), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_598), .B(n_478), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_553), .A2(n_541), .B(n_536), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_592), .B(n_533), .C(n_495), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_569), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_585), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_553), .B(n_535), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_563), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_559), .B(n_526), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_568), .B(n_535), .Y(n_642) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_551), .A2(n_477), .A3(n_479), .B1(n_489), .B2(n_509), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_556), .A2(n_505), .B1(n_535), .B2(n_543), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_577), .B(n_486), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_601), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_611), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_594), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_554), .B(n_495), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_603), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_550), .B(n_499), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_607), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_611), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_606), .B(n_544), .C(n_540), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_583), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_609), .Y(n_657) );
NAND2x1_ASAP7_75t_L g658 ( .A(n_583), .B(n_486), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_560), .B(n_499), .Y(n_659) );
OAI22xp33_ASAP7_75t_SL g660 ( .A1(n_579), .A2(n_503), .B1(n_533), .B2(n_507), .Y(n_660) );
NOR2xp33_ASAP7_75t_SL g661 ( .A(n_579), .B(n_503), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_590), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_583), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_628), .A2(n_605), .B1(n_548), .B2(n_562), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_619), .A2(n_558), .B1(n_547), .B2(n_577), .C(n_566), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g666 ( .A1(n_621), .A2(n_606), .B(n_578), .Y(n_666) );
O2A1O1Ixp5_ASAP7_75t_L g667 ( .A1(n_643), .A2(n_586), .B(n_614), .C(n_613), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_650), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_621), .A2(n_610), .B1(n_589), .B2(n_570), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_633), .B(n_618), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_620), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_622), .Y(n_672) );
OAI32xp33_ASAP7_75t_L g673 ( .A1(n_648), .A2(n_567), .A3(n_599), .B1(n_572), .B2(n_571), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_631), .Y(n_674) );
AOI211xp5_ASAP7_75t_SL g675 ( .A1(n_660), .A2(n_661), .B(n_610), .C(n_632), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g676 ( .A1(n_635), .A2(n_581), .B(n_589), .C(n_612), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_625), .A2(n_565), .B(n_595), .C(n_602), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_645), .A2(n_571), .B1(n_572), .B2(n_617), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_645), .A2(n_587), .B1(n_582), .B2(n_574), .C(n_584), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_637), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_624), .B(n_587), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_662), .A2(n_600), .B1(n_593), .B2(n_596), .Y(n_682) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_655), .A2(n_532), .B1(n_508), .B2(n_537), .C1(n_597), .C2(n_608), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_638), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_646), .A2(n_608), .B1(n_516), .B2(n_517), .C(n_525), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_627), .B(n_502), .Y(n_686) );
OA33x2_ASAP7_75t_L g687 ( .A1(n_623), .A2(n_502), .A3(n_516), .B1(n_517), .B2(n_525), .B3(n_542), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_667), .A2(n_639), .B(n_658), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_668), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_675), .B(n_629), .C(n_636), .Y(n_690) );
NOR2xp33_ASAP7_75t_SL g691 ( .A(n_682), .B(n_627), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_677), .B(n_636), .C(n_639), .D(n_644), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_679), .B(n_651), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_665), .A2(n_663), .B(n_656), .C(n_654), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_681), .B(n_657), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_673), .A2(n_653), .B1(n_654), .B2(n_656), .C(n_663), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_669), .A2(n_634), .B(n_650), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_664), .A2(n_659), .B(n_626), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_676), .A2(n_626), .B(n_640), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_688), .A2(n_683), .B(n_666), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_691), .B(n_683), .C(n_685), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_690), .B(n_671), .C(n_670), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_692), .B(n_684), .C(n_680), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_694), .A2(n_674), .B(n_672), .C(n_686), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_695), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_700), .B(n_698), .C(n_696), .D(n_697), .Y(n_706) );
NAND4xp75_ASAP7_75t_L g707 ( .A(n_705), .B(n_693), .C(n_699), .D(n_678), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_701), .B(n_689), .Y(n_708) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_702), .B(n_640), .C(n_647), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_708), .B(n_703), .Y(n_710) );
OA21x2_ASAP7_75t_L g711 ( .A1(n_707), .A2(n_704), .B(n_630), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_706), .B(n_647), .C(n_649), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_710), .B(n_709), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_711), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_714), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_713), .B(n_712), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_715), .Y(n_717) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_717), .A2(n_711), .B1(n_716), .B2(n_649), .Y(n_718) );
UNKNOWN g719 ( );
OAI21xp33_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_652), .B(n_641), .Y(n_720) );
OR2x6_ASAP7_75t_L g721 ( .A(n_720), .B(n_642), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_642), .B1(n_687), .B2(n_542), .Y(n_722) );
endmodule