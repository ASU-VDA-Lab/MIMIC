module fake_jpeg_28024_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_12),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_29),
.B(n_13),
.C(n_20),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_1),
.Y(n_29)
);

OA22x2_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_18),
.B1(n_12),
.B2(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_17),
.B1(n_26),
.B2(n_13),
.Y(n_40)
);

AO22x2_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_18),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_45),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_46),
.B(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_52),
.B1(n_21),
.B2(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_28),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_30),
.C(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_34),
.B1(n_21),
.B2(n_20),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_65),
.B(n_48),
.C(n_43),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_25),
.C(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_8),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_50),
.B(n_40),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_16),
.C(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_44),
.Y(n_74)
);

OAI22x1_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_14),
.B1(n_2),
.B2(n_4),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_65),
.B1(n_54),
.B2(n_63),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_39),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_16),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_61),
.C(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_79),
.B(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_68),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_76),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_67),
.A3(n_62),
.B1(n_69),
.B2(n_59),
.C1(n_73),
.C2(n_66),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_69),
.B(n_2),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_83),
.B1(n_80),
.B2(n_52),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_81),
.C(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_70),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_80),
.A3(n_69),
.B1(n_76),
.B2(n_70),
.C1(n_8),
.C2(n_7),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_97),
.B(n_10),
.Y(n_99)
);

XNOR2x1_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_10),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_92),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_99),
.A3(n_100),
.B1(n_1),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_1),
.B(n_2),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.C(n_6),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_42),
.Y(n_104)
);


endmodule