module real_aes_937_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_602;
wire n_552;
wire n_402;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_246;
wire n_412;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_393;
wire n_294;
wire n_258;
wire n_307;
wire n_601;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
NAND2xp5_ASAP7_75t_L g605 ( .A(n_0), .B(n_383), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_1), .A2(n_73), .B1(n_276), .B2(n_296), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_2), .A2(n_601), .B1(n_602), .B2(n_617), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_2), .Y(n_617) );
AO22x2_ASAP7_75t_L g240 ( .A1(n_3), .A2(n_158), .B1(n_230), .B2(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g597 ( .A(n_3), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_4), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_5), .A2(n_131), .B1(n_307), .B2(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_6), .A2(n_12), .B1(n_428), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_7), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_8), .A2(n_46), .B1(n_339), .B2(n_341), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_9), .A2(n_98), .B1(n_278), .B2(n_279), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_10), .A2(n_187), .B1(n_251), .B2(n_254), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_11), .A2(n_115), .B1(n_313), .B2(n_316), .Y(n_312) );
AO22x2_ASAP7_75t_L g237 ( .A1(n_13), .A2(n_44), .B1(n_230), .B2(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_13), .B(n_596), .Y(n_595) );
AO222x2_ASAP7_75t_L g547 ( .A1(n_14), .A2(n_43), .B1(n_170), .B2(n_226), .C1(n_254), .C2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_15), .A2(n_171), .B1(n_266), .B2(n_267), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_16), .A2(n_191), .B1(n_270), .B2(n_272), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_17), .A2(n_153), .B1(n_325), .B2(n_580), .Y(n_579) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_18), .A2(n_38), .B1(n_124), .B2(n_226), .C1(n_242), .C2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_19), .A2(n_175), .B1(n_339), .B2(n_377), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_20), .A2(n_21), .B1(n_278), .B2(n_279), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_22), .A2(n_176), .B1(n_245), .B2(n_552), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_23), .A2(n_130), .B1(n_179), .B2(n_345), .C1(n_348), .C2(n_351), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_24), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_25), .A2(n_182), .B1(n_331), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_26), .A2(n_82), .B1(n_276), .B2(n_296), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_27), .A2(n_167), .B1(n_334), .B2(n_517), .Y(n_571) );
OA22x2_ASAP7_75t_L g435 ( .A1(n_28), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_28), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g417 ( .A1(n_29), .A2(n_108), .B1(n_206), .B2(n_345), .C1(n_418), .C2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_30), .A2(n_148), .B1(n_251), .B2(n_254), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_31), .A2(n_93), .B1(n_407), .B2(n_517), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_32), .A2(n_95), .B1(n_321), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_33), .A2(n_84), .B1(n_251), .B2(n_257), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_34), .A2(n_65), .B1(n_369), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_35), .A2(n_200), .B1(n_334), .B2(n_336), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_36), .A2(n_201), .B1(n_452), .B2(n_454), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_37), .A2(n_194), .B1(n_351), .B2(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_39), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_40), .A2(n_142), .B1(n_360), .B2(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_41), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_42), .A2(n_135), .B1(n_321), .B2(n_325), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_45), .A2(n_102), .B1(n_307), .B2(n_310), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_47), .A2(n_91), .B1(n_364), .B2(n_365), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_48), .A2(n_105), .B1(n_370), .B2(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_49), .A2(n_196), .B1(n_379), .B2(n_380), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g265 ( .A1(n_50), .A2(n_178), .B1(n_266), .B2(n_267), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_51), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_52), .A2(n_155), .B1(n_369), .B2(n_370), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_53), .A2(n_109), .B1(n_370), .B2(n_401), .Y(n_429) );
OAI22x1_ASAP7_75t_L g513 ( .A1(n_54), .A2(n_514), .B1(n_534), .B2(n_535), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_54), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_55), .A2(n_92), .B1(n_257), .B2(n_260), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_56), .A2(n_136), .B1(n_270), .B2(n_278), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_57), .A2(n_184), .B1(n_272), .B2(n_276), .Y(n_558) );
INVx3_ASAP7_75t_L g230 ( .A(n_58), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_59), .A2(n_126), .B1(n_275), .B2(n_279), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_60), .A2(n_129), .B1(n_405), .B2(n_419), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_61), .A2(n_159), .B1(n_310), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_62), .A2(n_154), .B1(n_336), .B2(n_374), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_63), .A2(n_143), .B1(n_334), .B2(n_517), .Y(n_516) );
OA22x2_ASAP7_75t_L g355 ( .A1(n_64), .A2(n_356), .B1(n_357), .B2(n_384), .Y(n_355) );
INVxp67_ASAP7_75t_L g384 ( .A(n_64), .Y(n_384) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_66), .B(n_603), .Y(n_622) );
INVxp67_ASAP7_75t_L g627 ( .A(n_66), .Y(n_627) );
AO222x2_ASAP7_75t_L g225 ( .A1(n_67), .A2(n_113), .B1(n_134), .B2(n_226), .C1(n_242), .C2(n_245), .Y(n_225) );
INVx1_ASAP7_75t_L g353 ( .A(n_68), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_69), .A2(n_145), .B1(n_267), .B2(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_70), .A2(n_118), .B1(n_257), .B2(n_260), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_71), .A2(n_192), .B1(n_379), .B2(n_380), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_72), .Y(n_462) );
INVx1_ASAP7_75t_SL g231 ( .A(n_74), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_74), .B(n_100), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_75), .Y(n_444) );
INVx2_ASAP7_75t_L g214 ( .A(n_76), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_77), .A2(n_147), .B1(n_316), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_78), .A2(n_138), .B1(n_365), .B2(n_524), .Y(n_616) );
OA22x2_ASAP7_75t_L g390 ( .A1(n_79), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_79), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_80), .A2(n_117), .B1(n_310), .B2(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_81), .A2(n_188), .B1(n_275), .B2(n_276), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_83), .A2(n_177), .B1(n_424), .B2(n_426), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_85), .A2(n_202), .B1(n_401), .B2(n_472), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_86), .A2(n_156), .B1(n_327), .B2(n_330), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_87), .A2(n_114), .B1(n_446), .B2(n_448), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_88), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_89), .A2(n_111), .B1(n_407), .B2(n_408), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_90), .B(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_94), .A2(n_112), .B1(n_307), .B2(n_424), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_96), .A2(n_204), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_97), .A2(n_104), .B1(n_313), .B2(n_362), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_99), .A2(n_186), .B1(n_339), .B2(n_405), .Y(n_404) );
AO22x2_ASAP7_75t_L g233 ( .A1(n_100), .A2(n_164), .B1(n_230), .B2(n_234), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_101), .A2(n_183), .B1(n_407), .B2(n_408), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_103), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_106), .A2(n_123), .B1(n_334), .B2(n_408), .Y(n_500) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_107), .A2(n_208), .B(n_215), .C(n_599), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_110), .A2(n_189), .B1(n_313), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_116), .A2(n_125), .B1(n_321), .B2(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g232 ( .A(n_119), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_120), .A2(n_174), .B1(n_242), .B2(n_245), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_121), .A2(n_151), .B1(n_313), .B2(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_122), .B(n_345), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_127), .A2(n_139), .B1(n_270), .B2(n_272), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_128), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_132), .A2(n_161), .B1(n_321), .B2(n_323), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_133), .A2(n_166), .B1(n_377), .B2(n_419), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_137), .A2(n_150), .B1(n_379), .B2(n_380), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_140), .A2(n_160), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_141), .A2(n_152), .B1(n_396), .B2(n_397), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_144), .A2(n_193), .B1(n_313), .B2(n_360), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_146), .A2(n_195), .B1(n_419), .B2(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_149), .B(n_569), .Y(n_568) );
CKINVDCx16_ASAP7_75t_R g298 ( .A(n_157), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_162), .A2(n_544), .B1(n_545), .B2(n_560), .Y(n_543) );
INVx1_ASAP7_75t_L g560 ( .A(n_162), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_163), .A2(n_203), .B1(n_360), .B2(n_531), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_165), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_168), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g593 ( .A(n_168), .Y(n_593) );
OA22x2_ASAP7_75t_L g412 ( .A1(n_169), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_169), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_172), .A2(n_198), .B1(n_341), .B2(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g211 ( .A(n_173), .Y(n_211) );
AND2x2_ASAP7_75t_R g619 ( .A(n_173), .B(n_593), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_180), .A2(n_197), .B1(n_351), .B2(n_379), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_181), .A2(n_205), .B1(n_351), .B2(n_379), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_185), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_190), .B(n_226), .Y(n_284) );
AOI22x1_ASAP7_75t_L g491 ( .A1(n_199), .A2(n_492), .B1(n_493), .B2(n_512), .Y(n_491) );
INVx1_ASAP7_75t_L g512 ( .A(n_199), .Y(n_512) );
XNOR2x1_ASAP7_75t_L g538 ( .A(n_199), .B(n_493), .Y(n_538) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_209), .B(n_212), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g626 ( .A(n_210), .B(n_212), .Y(n_626) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_211), .B(n_593), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_430), .B1(n_588), .B2(n_589), .C(n_590), .Y(n_215) );
INVx1_ASAP7_75t_L g588 ( .A(n_216), .Y(n_588) );
AOI22xp5_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_218), .B1(n_387), .B2(n_388), .Y(n_216) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_301), .B1(n_385), .B2(n_386), .Y(n_218) );
INVx1_ASAP7_75t_L g385 ( .A(n_219), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_280), .B1(n_299), .B2(n_300), .Y(n_219) );
INVx1_ASAP7_75t_L g299 ( .A(n_220), .Y(n_299) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
XNOR2x1_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_263), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_249), .Y(n_224) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_235), .Y(n_226) );
AND2x2_ASAP7_75t_L g254 ( .A(n_227), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g260 ( .A(n_227), .B(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g337 ( .A(n_227), .B(n_261), .Y(n_337) );
AND2x4_ASAP7_75t_L g343 ( .A(n_227), .B(n_255), .Y(n_343) );
AND2x2_ASAP7_75t_L g347 ( .A(n_227), .B(n_235), .Y(n_347) );
AND2x2_ASAP7_75t_L g521 ( .A(n_227), .B(n_255), .Y(n_521) );
AND2x2_ASAP7_75t_L g548 ( .A(n_227), .B(n_261), .Y(n_548) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_233), .Y(n_227) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
AND2x2_ASAP7_75t_L g247 ( .A(n_228), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
OAI22x1_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B1(n_231), .B2(n_232), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g234 ( .A(n_230), .Y(n_234) );
INVx2_ASAP7_75t_L g238 ( .A(n_230), .Y(n_238) );
INVx1_ASAP7_75t_L g241 ( .A(n_230), .Y(n_241) );
INVx2_ASAP7_75t_L g248 ( .A(n_233), .Y(n_248) );
AND2x2_ASAP7_75t_L g252 ( .A(n_233), .B(n_253), .Y(n_252) );
BUFx2_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
AND2x2_ASAP7_75t_L g270 ( .A(n_235), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_235), .B(n_247), .Y(n_275) );
AND2x6_ASAP7_75t_L g278 ( .A(n_235), .B(n_252), .Y(n_278) );
AND2x2_ASAP7_75t_L g296 ( .A(n_235), .B(n_247), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_235), .B(n_252), .Y(n_309) );
AND2x4_ASAP7_75t_L g315 ( .A(n_235), .B(n_271), .Y(n_315) );
AND2x4_ASAP7_75t_L g329 ( .A(n_235), .B(n_247), .Y(n_329) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_239), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g244 ( .A(n_237), .B(n_240), .Y(n_244) );
AND2x4_ASAP7_75t_L g246 ( .A(n_237), .B(n_239), .Y(n_246) );
INVx1_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
INVxp67_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g258 ( .A(n_240), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_SL g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g352 ( .A(n_243), .B(n_244), .Y(n_352) );
AND2x2_ASAP7_75t_SL g552 ( .A(n_243), .B(n_244), .Y(n_552) );
AND2x4_ASAP7_75t_L g267 ( .A(n_244), .B(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g276 ( .A(n_244), .B(n_271), .Y(n_276) );
AND2x4_ASAP7_75t_L g325 ( .A(n_244), .B(n_268), .Y(n_325) );
AND2x4_ASAP7_75t_L g331 ( .A(n_244), .B(n_271), .Y(n_331) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_245), .Y(n_533) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g251 ( .A(n_246), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g272 ( .A(n_246), .B(n_271), .Y(n_272) );
AND2x4_ASAP7_75t_L g311 ( .A(n_246), .B(n_271), .Y(n_311) );
AND2x4_ASAP7_75t_L g340 ( .A(n_246), .B(n_252), .Y(n_340) );
AND2x2_ASAP7_75t_L g350 ( .A(n_246), .B(n_247), .Y(n_350) );
AND2x2_ASAP7_75t_L g520 ( .A(n_246), .B(n_252), .Y(n_520) );
AND2x4_ASAP7_75t_L g257 ( .A(n_247), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g335 ( .A(n_247), .B(n_258), .Y(n_335) );
AND2x4_ASAP7_75t_L g271 ( .A(n_248), .B(n_253), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_256), .Y(n_249) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_252), .B(n_258), .Y(n_266) );
AND2x2_ASAP7_75t_L g292 ( .A(n_252), .B(n_258), .Y(n_292) );
AND2x2_ASAP7_75t_L g322 ( .A(n_252), .B(n_258), .Y(n_322) );
AND2x6_ASAP7_75t_L g279 ( .A(n_258), .B(n_271), .Y(n_279) );
AND2x4_ASAP7_75t_L g318 ( .A(n_258), .B(n_271), .Y(n_318) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_259), .Y(n_262) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_273), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
XOR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_298), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_282), .B(n_289), .Y(n_281) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NOR2x1_ASAP7_75t_L g289 ( .A(n_290), .B(n_294), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx2_ASAP7_75t_SL g386 ( .A(n_301), .Y(n_386) );
OA22x2_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_354), .B2(n_355), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
XOR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_353), .Y(n_303) );
NAND4xp75_ASAP7_75t_L g304 ( .A(n_305), .B(n_319), .C(n_332), .D(n_344), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_312), .Y(n_305) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g396 ( .A(n_308), .Y(n_396) );
INVx2_ASAP7_75t_SL g426 ( .A(n_308), .Y(n_426) );
INVx2_ASAP7_75t_L g477 ( .A(n_308), .Y(n_477) );
INVx3_ASAP7_75t_L g577 ( .A(n_308), .Y(n_577) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g526 ( .A(n_309), .Y(n_526) );
BUFx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_311), .Y(n_360) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_311), .Y(n_464) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_SL g469 ( .A(n_314), .Y(n_469) );
INVx4_ASAP7_75t_L g511 ( .A(n_314), .Y(n_511) );
INVx2_ASAP7_75t_L g531 ( .A(n_314), .Y(n_531) );
INVx8_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g362 ( .A(n_317), .Y(n_362) );
INVx1_ASAP7_75t_SL g397 ( .A(n_317), .Y(n_397) );
INVx2_ASAP7_75t_SL g424 ( .A(n_317), .Y(n_424) );
INVx2_ASAP7_75t_L g480 ( .A(n_317), .Y(n_480) );
INVx2_ASAP7_75t_SL g578 ( .A(n_317), .Y(n_578) );
INVx8_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_326), .Y(n_319) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g367 ( .A(n_322), .Y(n_367) );
BUFx3_ASAP7_75t_L g580 ( .A(n_322), .Y(n_580) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx3_ASAP7_75t_L g428 ( .A(n_324), .Y(n_428) );
OAI22xp33_ASAP7_75t_SL g482 ( .A1(n_324), .A2(n_483), .B1(n_486), .B2(n_487), .Y(n_482) );
INVx5_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
BUFx2_ASAP7_75t_L g524 ( .A(n_325), .Y(n_524) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g369 ( .A(n_328), .Y(n_369) );
INVx2_ASAP7_75t_L g401 ( .A(n_328), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_328), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_460) );
INVx6_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx3_ASAP7_75t_L g529 ( .A(n_329), .Y(n_529) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g371 ( .A(n_331), .Y(n_371) );
BUFx2_ASAP7_75t_SL g472 ( .A(n_331), .Y(n_472) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_338), .Y(n_332) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_335), .Y(n_407) );
BUFx6f_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx4f_ASAP7_75t_L g408 ( .A(n_337), .Y(n_408) );
BUFx3_ASAP7_75t_L g455 ( .A(n_337), .Y(n_455) );
INVx2_ASAP7_75t_L g518 ( .A(n_337), .Y(n_518) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g419 ( .A(n_340), .Y(n_419) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_340), .Y(n_458) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
INVx2_ASAP7_75t_SL g405 ( .A(n_342), .Y(n_405) );
INVx2_ASAP7_75t_SL g418 ( .A(n_342), .Y(n_418) );
INVx2_ASAP7_75t_L g573 ( .A(n_342), .Y(n_573) );
INVx6_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g496 ( .A(n_345), .Y(n_496) );
INVx4_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
INVx3_ASAP7_75t_SL g443 ( .A(n_346), .Y(n_443) );
INVx3_ASAP7_75t_L g569 ( .A(n_346), .Y(n_569) );
INVx6_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g567 ( .A(n_349), .Y(n_567) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx5_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
BUFx3_ASAP7_75t_L g449 ( .A(n_350), .Y(n_449) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
NOR2x1_ASAP7_75t_L g357 ( .A(n_358), .B(n_372), .Y(n_357) );
NAND4xp25_ASAP7_75t_SL g358 ( .A(n_359), .B(n_361), .C(n_363), .D(n_368), .Y(n_358) );
INVx1_ASAP7_75t_L g613 ( .A(n_360), .Y(n_613) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g485 ( .A(n_366), .Y(n_485) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g615 ( .A(n_371), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .C(n_378), .D(n_382), .Y(n_372) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g453 ( .A(n_375), .Y(n_453) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g447 ( .A(n_381), .Y(n_447) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_390), .B1(n_410), .B2(n_411), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_402), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .C(n_399), .D(n_400), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .C(n_406), .D(n_409), .Y(n_402) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_422), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .C(n_421), .Y(n_416) );
NAND4xp25_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .C(n_427), .D(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g589 ( .A(n_430), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_541), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_488), .B1(n_489), .B2(n_539), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_435), .Y(n_540) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND3x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_459), .C(n_473), .Y(n_438) );
NOR2xp67_ASAP7_75t_SL g439 ( .A(n_440), .B(n_450), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_444), .B(n_445), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_451), .B(n_456), .Y(n_450) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_465), .Y(n_459) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B1(n_470), .B2(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
OAI22xp33_ASAP7_75t_SL g474 ( .A1(n_475), .A2(n_478), .B1(n_479), .B2(n_481), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g505 ( .A(n_485), .Y(n_505) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AO22x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_513), .B1(n_536), .B2(n_537), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_502), .Y(n_493) );
NOR2xp67_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .Y(n_494) );
OAI21xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_497), .B(n_498), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g536 ( .A(n_513), .Y(n_536) );
NAND4xp25_ASAP7_75t_SL g514 ( .A(n_515), .B(n_522), .C(n_527), .D(n_532), .Y(n_514) );
AND4x1_ASAP7_75t_L g534 ( .A(n_515), .B(n_522), .C(n_527), .D(n_532), .Y(n_534) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_561), .B1(n_585), .B2(n_586), .Y(n_541) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_542), .Y(n_587) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_553), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g585 ( .A(n_561), .Y(n_585) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
XOR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_584), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_564), .B(n_574), .Y(n_563) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_570), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_581), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_592), .B(n_595), .Y(n_625) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
OAI222xp33_ASAP7_75t_R g599 ( .A1(n_600), .A2(n_618), .B1(n_620), .B2(n_623), .C1(n_626), .C2(n_627), .Y(n_599) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVxp33_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2xp67_ASAP7_75t_L g603 ( .A(n_604), .B(n_609), .Y(n_603) );
NAND4xp25_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .C(n_607), .D(n_608), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .C(n_614), .D(n_616), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
CKINVDCx6p67_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
endmodule