module real_aes_752_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_0), .B(n_136), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_1), .A2(n_130), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_2), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_3), .B(n_136), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_4), .B(n_147), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_5), .B(n_147), .Y(n_222) );
INVx1_ASAP7_75t_L g135 ( .A(n_6), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_7), .B(n_147), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g752 ( .A(n_8), .Y(n_752) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_9), .B(n_145), .Y(n_198) );
AND2x2_ASAP7_75t_L g449 ( .A(n_10), .B(n_192), .Y(n_449) );
AND2x2_ASAP7_75t_L g457 ( .A(n_11), .B(n_159), .Y(n_457) );
INVx2_ASAP7_75t_L g127 ( .A(n_12), .Y(n_127) );
AOI221x1_ASAP7_75t_L g129 ( .A1(n_13), .A2(n_25), .B1(n_130), .B2(n_136), .C(n_143), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_14), .B(n_147), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_15), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_16), .Y(n_104) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_17), .A2(n_192), .B(n_193), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_18), .B(n_136), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_19), .B(n_125), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_20), .B(n_147), .Y(n_206) );
AO21x1_ASAP7_75t_L g217 ( .A1(n_21), .A2(n_136), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_22), .B(n_136), .Y(n_488) );
INVx1_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_24), .A2(n_88), .B1(n_136), .B2(n_518), .Y(n_517) );
NAND2x1_ASAP7_75t_L g155 ( .A(n_26), .B(n_147), .Y(n_155) );
NAND2x1_ASAP7_75t_L g185 ( .A(n_27), .B(n_145), .Y(n_185) );
OR2x2_ASAP7_75t_L g128 ( .A(n_28), .B(n_85), .Y(n_128) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_28), .A2(n_85), .B(n_127), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_29), .B(n_145), .Y(n_180) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_30), .A2(n_114), .B1(n_727), .B2(n_730), .C(n_731), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g730 ( .A(n_30), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_31), .B(n_147), .Y(n_197) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_32), .A2(n_159), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_33), .B(n_145), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_34), .A2(n_130), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_35), .B(n_147), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_36), .A2(n_130), .B(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g131 ( .A(n_37), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g142 ( .A(n_37), .B(n_135), .Y(n_142) );
INVx1_ASAP7_75t_L g526 ( .A(n_37), .Y(n_526) );
OR2x6_ASAP7_75t_L g109 ( .A(n_38), .B(n_110), .Y(n_109) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_38), .B(n_751), .C(n_753), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_39), .B(n_136), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_40), .B(n_136), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_41), .B(n_147), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_42), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_43), .B(n_145), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_44), .B(n_136), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_45), .A2(n_130), .B(n_453), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_46), .A2(n_130), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_47), .B(n_145), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_48), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_49), .B(n_145), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_50), .B(n_136), .Y(n_462) );
INVx1_ASAP7_75t_L g134 ( .A(n_51), .Y(n_134) );
INVx1_ASAP7_75t_L g139 ( .A(n_51), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_52), .B(n_147), .Y(n_455) );
OAI22xp33_ASAP7_75t_SL g742 ( .A1(n_53), .A2(n_425), .B1(n_426), .B2(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_53), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_54), .Y(n_732) );
AND2x2_ASAP7_75t_L g479 ( .A(n_55), .B(n_125), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_56), .B(n_145), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_57), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_58), .B(n_145), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_59), .A2(n_130), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_60), .B(n_136), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_61), .B(n_136), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_62), .A2(n_130), .B(n_470), .Y(n_469) );
AO21x1_ASAP7_75t_L g219 ( .A1(n_63), .A2(n_130), .B(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g494 ( .A(n_64), .B(n_126), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_65), .B(n_136), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_66), .B(n_145), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_67), .B(n_136), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_68), .B(n_145), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_69), .A2(n_93), .B1(n_130), .B2(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g170 ( .A(n_70), .B(n_126), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_71), .B(n_147), .Y(n_491) );
INVx1_ASAP7_75t_L g132 ( .A(n_72), .Y(n_132) );
INVx1_ASAP7_75t_L g141 ( .A(n_72), .Y(n_141) );
AND2x2_ASAP7_75t_L g189 ( .A(n_73), .B(n_159), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_74), .B(n_145), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_75), .A2(n_130), .B(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_76), .A2(n_130), .B(n_436), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_77), .A2(n_130), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g474 ( .A(n_78), .B(n_126), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_79), .B(n_125), .Y(n_515) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_80), .B(n_111), .Y(n_754) );
AND2x2_ASAP7_75t_L g174 ( .A(n_81), .B(n_159), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_82), .B(n_136), .Y(n_208) );
AND2x2_ASAP7_75t_L g439 ( .A(n_83), .B(n_192), .Y(n_439) );
AND2x2_ASAP7_75t_L g218 ( .A(n_84), .B(n_199), .Y(n_218) );
AND2x2_ASAP7_75t_L g162 ( .A(n_86), .B(n_159), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_87), .B(n_145), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_89), .B(n_147), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_90), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_91), .A2(n_130), .B(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_92), .A2(n_130), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_94), .B(n_147), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_95), .B(n_147), .Y(n_179) );
BUFx2_ASAP7_75t_L g493 ( .A(n_96), .Y(n_493) );
BUFx2_ASAP7_75t_L g738 ( .A(n_97), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_98), .A2(n_130), .B(n_196), .Y(n_195) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_745), .B(n_755), .Y(n_99) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_734), .B(n_739), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_113), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
AOI21xp5_ASAP7_75t_SL g741 ( .A1(n_103), .A2(n_742), .B(n_744), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g744 ( .A(n_106), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x6_ASAP7_75t_SL g424 ( .A(n_107), .B(n_108), .Y(n_424) );
AND2x6_ASAP7_75t_SL g726 ( .A(n_107), .B(n_109), .Y(n_726) );
OR2x2_ASAP7_75t_L g733 ( .A(n_107), .B(n_109), .Y(n_733) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_107), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OAI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_422), .B1(n_425), .B2(n_725), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_116), .A2(n_424), .B1(n_426), .B2(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_334), .Y(n_116) );
AND4x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_246), .C(n_273), .D(n_308), .Y(n_117) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_171), .B1(n_211), .B2(n_226), .C(n_230), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_150), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_121), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g287 ( .A(n_122), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g342 ( .A(n_122), .B(n_297), .Y(n_342) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g245 ( .A(n_123), .B(n_163), .Y(n_245) );
AND2x4_ASAP7_75t_L g281 ( .A(n_123), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g295 ( .A(n_123), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g212 ( .A(n_124), .Y(n_212) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_124), .Y(n_384) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_149), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_125), .A2(n_176), .B(n_177), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_125), .Y(n_188) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_125), .A2(n_129), .B(n_149), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_125), .A2(n_434), .B(n_435), .Y(n_433) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_125), .A2(n_517), .B(n_523), .Y(n_516) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g199 ( .A(n_127), .B(n_128), .Y(n_199) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
BUFx3_ASAP7_75t_L g522 ( .A(n_131), .Y(n_522) );
AND2x6_ASAP7_75t_L g145 ( .A(n_132), .B(n_138), .Y(n_145) );
INVx2_ASAP7_75t_L g528 ( .A(n_132), .Y(n_528) );
AND2x4_ASAP7_75t_L g524 ( .A(n_133), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g147 ( .A(n_134), .B(n_140), .Y(n_147) );
INVx2_ASAP7_75t_L g520 ( .A(n_134), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_135), .Y(n_521) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_142), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_146), .B(n_148), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_145), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_148), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_148), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_148), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_148), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_148), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_148), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_148), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_148), .A2(n_437), .B(n_438), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_148), .A2(n_446), .B(n_447), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_148), .A2(n_454), .B(n_455), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_148), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_148), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_148), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_148), .A2(n_491), .B(n_492), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_SL g239 ( .A1(n_150), .A2(n_212), .B(n_240), .C(n_244), .Y(n_239) );
AND2x2_ASAP7_75t_L g260 ( .A(n_150), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_150), .B(n_212), .Y(n_400) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_163), .Y(n_150) );
INVx2_ASAP7_75t_L g280 ( .A(n_151), .Y(n_280) );
BUFx3_ASAP7_75t_L g296 ( .A(n_151), .Y(n_296) );
INVxp67_ASAP7_75t_L g300 ( .A(n_151), .Y(n_300) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_158), .B(n_162), .Y(n_151) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_152), .A2(n_158), .B(n_162), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_158), .A2(n_164), .B(n_170), .Y(n_163) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_158), .A2(n_164), .B(n_170), .Y(n_225) );
AO21x1_ASAP7_75t_SL g467 ( .A1(n_158), .A2(n_468), .B(n_474), .Y(n_467) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_158), .A2(n_468), .B(n_474), .Y(n_501) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_160), .A2(n_451), .B(n_457), .Y(n_450) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx4f_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
INVx2_ASAP7_75t_L g279 ( .A(n_163), .Y(n_279) );
AND2x2_ASAP7_75t_L g285 ( .A(n_163), .B(n_258), .Y(n_285) );
AND2x2_ASAP7_75t_L g311 ( .A(n_163), .B(n_280), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_165), .B(n_169), .Y(n_164) );
AOI211xp5_ASAP7_75t_L g308 ( .A1(n_171), .A2(n_309), .B(n_312), .C(n_322), .Y(n_308) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_172), .B(n_190), .Y(n_171) );
OAI321xp33_ASAP7_75t_L g283 ( .A1(n_172), .A2(n_231), .A3(n_284), .B1(n_286), .B2(n_287), .C(n_289), .Y(n_283) );
AND2x2_ASAP7_75t_L g404 ( .A(n_172), .B(n_379), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_172), .Y(n_407) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_181), .Y(n_172) );
INVx5_ASAP7_75t_L g229 ( .A(n_173), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_173), .B(n_243), .Y(n_242) );
NOR2x1_ASAP7_75t_SL g274 ( .A(n_173), .B(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
AND2x2_ASAP7_75t_L g421 ( .A(n_173), .B(n_191), .Y(n_421) );
OR2x6_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
AND2x2_ASAP7_75t_L g228 ( .A(n_181), .B(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_181), .Y(n_238) );
INVx4_ASAP7_75t_L g243 ( .A(n_181), .Y(n_243) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_188), .B(n_189), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
AOI21x1_ASAP7_75t_L g442 ( .A1(n_188), .A2(n_443), .B(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g286 ( .A(n_190), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_R g389 ( .A1(n_190), .A2(n_228), .B(n_260), .C(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g409 ( .A(n_190), .B(n_234), .Y(n_409) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
INVx1_ASAP7_75t_L g227 ( .A(n_191), .Y(n_227) );
INVx2_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
OR2x2_ASAP7_75t_L g252 ( .A(n_191), .B(n_243), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_191), .B(n_275), .Y(n_321) );
BUFx3_ASAP7_75t_L g328 ( .A(n_191), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_192), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_199), .Y(n_193) );
INVx1_ASAP7_75t_SL g202 ( .A(n_199), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_199), .B(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_199), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_199), .A2(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g291 ( .A(n_200), .Y(n_291) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_200), .Y(n_304) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g237 ( .A(n_201), .Y(n_237) );
INVx1_ASAP7_75t_L g346 ( .A(n_201), .Y(n_346) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_209), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_202), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_202), .A2(n_203), .B(n_209), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_208), .Y(n_203) );
AND2x2_ASAP7_75t_L g247 ( .A(n_211), .B(n_248), .Y(n_247) );
OAI31xp33_ASAP7_75t_L g398 ( .A1(n_211), .A2(n_399), .A3(n_401), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_SL g416 ( .A(n_211), .Y(n_416) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AOI21xp33_ASAP7_75t_L g230 ( .A1(n_212), .A2(n_231), .B(n_239), .Y(n_230) );
NAND2x1_ASAP7_75t_L g310 ( .A(n_212), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g339 ( .A(n_212), .Y(n_339) );
INVx2_ASAP7_75t_L g288 ( .A(n_213), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_213), .B(n_271), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_213), .B(n_270), .Y(n_380) );
NOR2xp33_ASAP7_75t_SL g388 ( .A(n_213), .B(n_339), .Y(n_388) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
AND2x2_ASAP7_75t_SL g257 ( .A(n_214), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g268 ( .A(n_214), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g297 ( .A(n_214), .B(n_279), .Y(n_297) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g261 ( .A(n_215), .Y(n_261) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g282 ( .A(n_216), .Y(n_282) );
OAI21x1_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_219), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g224 ( .A(n_218), .Y(n_224) );
INVx2_ASAP7_75t_L g269 ( .A(n_225), .Y(n_269) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_225), .Y(n_329) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
AND2x2_ASAP7_75t_L g344 ( .A(n_227), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g255 ( .A(n_228), .B(n_249), .Y(n_255) );
INVx2_ASAP7_75t_SL g303 ( .A(n_228), .Y(n_303) );
INVx4_ASAP7_75t_L g234 ( .A(n_229), .Y(n_234) );
AND2x2_ASAP7_75t_L g332 ( .A(n_229), .B(n_275), .Y(n_332) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_229), .B(n_345), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_229), .B(n_243), .Y(n_367) );
INVx1_ASAP7_75t_L g373 ( .A(n_231), .Y(n_373) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
OR2x2_ASAP7_75t_L g305 ( .A(n_232), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
OR2x2_ASAP7_75t_L g357 ( .A(n_233), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g387 ( .A(n_233), .B(n_275), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_234), .B(n_237), .Y(n_263) );
AND2x2_ASAP7_75t_L g355 ( .A(n_234), .B(n_345), .Y(n_355) );
AND2x4_ASAP7_75t_L g417 ( .A(n_234), .B(n_296), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
INVx2_ASAP7_75t_L g241 ( .A(n_236), .Y(n_241) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp67_ASAP7_75t_SL g240 ( .A(n_241), .B(n_242), .Y(n_240) );
OAI322xp33_ASAP7_75t_SL g253 ( .A1(n_241), .A2(n_254), .A3(n_256), .B1(n_259), .B2(n_262), .C1(n_264), .C2(n_266), .Y(n_253) );
INVx1_ASAP7_75t_L g411 ( .A(n_241), .Y(n_411) );
OR2x2_ASAP7_75t_L g264 ( .A(n_242), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g290 ( .A(n_243), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_243), .B(n_291), .Y(n_306) );
INVx2_ASAP7_75t_L g333 ( .A(n_243), .Y(n_333) );
AND2x4_ASAP7_75t_L g345 ( .A(n_243), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_245), .B(n_261), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_251), .B(n_253), .Y(n_246) );
AND2x2_ASAP7_75t_L g314 ( .A(n_248), .B(n_281), .Y(n_314) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_249), .B(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g272 ( .A(n_250), .Y(n_272) );
AND2x4_ASAP7_75t_SL g354 ( .A(n_250), .B(n_269), .Y(n_354) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g262 ( .A(n_252), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_255), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g390 ( .A(n_257), .B(n_354), .Y(n_390) );
NOR4xp25_ASAP7_75t_L g394 ( .A(n_257), .B(n_271), .C(n_311), .D(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g271 ( .A(n_258), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g307 ( .A(n_258), .B(n_282), .Y(n_307) );
AND2x4_ASAP7_75t_L g371 ( .A(n_258), .B(n_282), .Y(n_371) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_261), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
OR2x2_ASAP7_75t_L g360 ( .A(n_268), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g414 ( .A(n_268), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_269), .B(n_281), .Y(n_315) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AOI211xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_276), .B(n_283), .C(n_298), .Y(n_273) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_279), .B(n_282), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_280), .B(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g362 ( .A(n_280), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_281), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g377 ( .A(n_281), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .B(n_293), .Y(n_289) );
AND2x4_ASAP7_75t_L g326 ( .A(n_290), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g420 ( .A(n_290), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_SL g324 ( .A(n_296), .Y(n_324) );
AND2x2_ASAP7_75t_L g383 ( .A(n_297), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g397 ( .A(n_297), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_301), .B(n_305), .C(n_307), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_299), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g375 ( .A(n_300), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g396 ( .A(n_300), .B(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
OR2x2_ASAP7_75t_L g385 ( .A(n_303), .B(n_327), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_306), .A2(n_313), .B1(n_315), .B2(n_316), .Y(n_312) );
INVx1_ASAP7_75t_SL g403 ( .A(n_307), .Y(n_403) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_318), .B(n_327), .Y(n_369) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_321), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B1(n_329), .B2(n_330), .Y(n_322) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI21xp5_ASAP7_75t_SL g336 ( .A1(n_327), .A2(n_337), .B(n_340), .Y(n_336) );
AND2x2_ASAP7_75t_L g365 ( .A(n_327), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND3x2_ASAP7_75t_L g331 ( .A(n_328), .B(n_332), .C(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g393 ( .A(n_328), .B(n_350), .Y(n_393) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g378 ( .A(n_333), .B(n_379), .Y(n_378) );
NOR2xp67_ASAP7_75t_L g334 ( .A(n_335), .B(n_391), .Y(n_334) );
NAND4xp25_ASAP7_75t_L g335 ( .A(n_336), .B(n_351), .C(n_372), .D(n_389), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_347), .B2(n_349), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_343), .A2(n_357), .B1(n_377), .B2(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g358 ( .A(n_345), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_347), .A2(n_370), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_356), .B2(n_359), .C(n_363), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_368), .B1(n_369), .B2(n_370), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_366), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_366), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_378), .B2(n_380), .C(n_381), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_375), .B(n_377), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B1(n_386), .B2(n_388), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g406 ( .A1(n_387), .A2(n_407), .B(n_408), .C(n_410), .Y(n_406) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_398), .C(n_405), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_418), .Y(n_405) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
CKINVDCx11_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_427), .B(n_633), .Y(n_426) );
NOR3xp33_ASAP7_75t_SL g427 ( .A(n_428), .B(n_556), .C(n_591), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_458), .B(n_508), .C(n_546), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_440), .Y(n_430) );
AND2x2_ASAP7_75t_L g539 ( .A(n_431), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_431), .B(n_545), .Y(n_579) );
AND2x2_ASAP7_75t_L g604 ( .A(n_431), .B(n_559), .Y(n_604) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g511 ( .A(n_432), .Y(n_511) );
OR2x2_ASAP7_75t_L g542 ( .A(n_432), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g550 ( .A(n_432), .B(n_450), .Y(n_550) );
AND2x2_ASAP7_75t_L g558 ( .A(n_432), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g585 ( .A(n_432), .B(n_586), .Y(n_585) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_432), .B(n_588), .Y(n_596) );
AND2x4_ASAP7_75t_L g613 ( .A(n_432), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g651 ( .A(n_432), .Y(n_651) );
AND2x4_ASAP7_75t_SL g656 ( .A(n_432), .B(n_441), .Y(n_656) );
OR2x6_ASAP7_75t_L g432 ( .A(n_433), .B(n_439), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_440), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_440), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_450), .Y(n_440) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_441), .Y(n_551) );
INVx2_ASAP7_75t_L g587 ( .A(n_441), .Y(n_587) );
INVx1_ASAP7_75t_L g614 ( .A(n_441), .Y(n_614) );
AND2x2_ASAP7_75t_L g713 ( .A(n_441), .B(n_623), .Y(n_713) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_442), .Y(n_545) );
AND2x2_ASAP7_75t_L g559 ( .A(n_442), .B(n_450), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_448), .Y(n_443) );
INVx2_ASAP7_75t_L g588 ( .A(n_450), .Y(n_588) );
INVx2_ASAP7_75t_L g623 ( .A(n_450), .Y(n_623) );
OR2x2_ASAP7_75t_L g708 ( .A(n_450), .B(n_540), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_456), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_475), .B(n_495), .C(n_502), .Y(n_458) );
INVx2_ASAP7_75t_SL g597 ( .A(n_459), .Y(n_597) );
AND2x2_ASAP7_75t_L g603 ( .A(n_459), .B(n_476), .Y(n_603) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
INVx1_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
INVx2_ASAP7_75t_L g530 ( .A(n_460), .Y(n_530) );
AND2x2_ASAP7_75t_L g554 ( .A(n_460), .B(n_478), .Y(n_554) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_460), .Y(n_583) );
OR2x2_ASAP7_75t_L g663 ( .A(n_460), .B(n_486), .Y(n_663) );
AND2x2_ASAP7_75t_L g529 ( .A(n_467), .B(n_530), .Y(n_529) );
NOR2x1_ASAP7_75t_SL g561 ( .A(n_467), .B(n_486), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g575 ( .A(n_476), .B(n_498), .Y(n_575) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
OR2x2_ASAP7_75t_L g507 ( .A(n_477), .B(n_486), .Y(n_507) );
BUFx2_ASAP7_75t_L g531 ( .A(n_477), .Y(n_531) );
NOR2xp67_ASAP7_75t_L g582 ( .A(n_477), .B(n_583), .Y(n_582) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
AND2x2_ASAP7_75t_L g560 ( .A(n_478), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g570 ( .A(n_478), .Y(n_570) );
NAND2x1_ASAP7_75t_L g608 ( .A(n_478), .B(n_486), .Y(n_608) );
OR2x2_ASAP7_75t_L g683 ( .A(n_478), .B(n_500), .Y(n_683) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx2_ASAP7_75t_SL g496 ( .A(n_486), .Y(n_496) );
AND2x2_ASAP7_75t_L g555 ( .A(n_486), .B(n_500), .Y(n_555) );
AND2x2_ASAP7_75t_L g626 ( .A(n_486), .B(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g647 ( .A(n_486), .Y(n_647) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_494), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g569 ( .A(n_498), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
BUFx2_ASAP7_75t_L g564 ( .A(n_499), .Y(n_564) );
AND2x2_ASAP7_75t_L g536 ( .A(n_500), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g627 ( .A(n_500), .Y(n_627) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
OR2x2_ASAP7_75t_L g573 ( .A(n_504), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_SL g615 ( .A(n_504), .B(n_616), .Y(n_615) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_504), .A2(n_531), .A3(n_653), .B1(n_655), .B2(n_658), .C1(n_660), .C2(n_662), .Y(n_652) );
AND2x2_ASAP7_75t_L g717 ( .A(n_504), .B(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_505), .B(n_531), .Y(n_541) );
AOI322xp5_ASAP7_75t_L g592 ( .A1(n_506), .A2(n_593), .A3(n_597), .B1(n_598), .B2(n_601), .C1(n_603), .C2(n_604), .Y(n_592) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g644 ( .A(n_507), .B(n_597), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_507), .A2(n_704), .B1(n_706), .B2(n_709), .Y(n_703) );
OR2x2_ASAP7_75t_L g721 ( .A(n_507), .B(n_670), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_531), .B(n_532), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
AOI221xp5_ASAP7_75t_SL g571 ( .A1(n_510), .A2(n_547), .B1(n_572), .B2(n_575), .C(n_576), .Y(n_571) );
AND2x2_ASAP7_75t_L g598 ( .A(n_510), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_511), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g640 ( .A(n_511), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g669 ( .A(n_512), .Y(n_669) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_529), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_513), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g611 ( .A(n_513), .Y(n_611) );
OR2x2_ASAP7_75t_L g618 ( .A(n_513), .B(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g661 ( .A(n_514), .B(n_623), .Y(n_661) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AND2x4_ASAP7_75t_L g540 ( .A(n_515), .B(n_516), .Y(n_540) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
NOR2x1p5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_529), .B(n_590), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_529), .B(n_570), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_529), .Y(n_670) );
INVx1_ASAP7_75t_L g537 ( .A(n_530), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_538), .B1(n_541), .B2(n_542), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_SL g648 ( .A(n_536), .Y(n_648) );
AND2x2_ASAP7_75t_L g705 ( .A(n_537), .B(n_561), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_539), .B(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_SL g577 ( .A(n_539), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_539), .B(n_698), .Y(n_697) );
BUFx3_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
INVx2_ASAP7_75t_L g595 ( .A(n_540), .Y(n_595) );
AND2x2_ASAP7_75t_L g638 ( .A(n_540), .B(n_622), .Y(n_638) );
INVx1_ASAP7_75t_L g552 ( .A(n_542), .Y(n_552) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI21xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_552), .B(n_553), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g631 ( .A(n_550), .Y(n_631) );
INVx2_ASAP7_75t_L g619 ( .A(n_551), .Y(n_619) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g616 ( .A(n_555), .B(n_570), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_555), .A2(n_653), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_557), .B(n_571), .Y(n_556) );
AOI32xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .A3(n_562), .B1(n_566), .B2(n_569), .Y(n_557) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_558), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_558), .A2(n_647), .B1(n_665), .B2(n_667), .C(n_673), .Y(n_664) );
AND2x2_ASAP7_75t_L g684 ( .A(n_558), .B(n_565), .Y(n_684) );
BUFx2_ASAP7_75t_L g568 ( .A(n_559), .Y(n_568) );
INVx1_ASAP7_75t_L g693 ( .A(n_559), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_559), .Y(n_698) );
INVx1_ASAP7_75t_SL g691 ( .A(n_560), .Y(n_691) );
INVx2_ASAP7_75t_L g574 ( .A(n_561), .Y(n_574) );
AND2x2_ASAP7_75t_L g686 ( .A(n_562), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g658 ( .A(n_564), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g630 ( .A(n_565), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_565), .B(n_656), .Y(n_678) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g590 ( .A(n_570), .Y(n_590) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g580 ( .A(n_574), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g589 ( .A(n_574), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g694 ( .A(n_575), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B1(n_584), .B2(n_589), .Y(n_576) );
INVx2_ASAP7_75t_SL g668 ( .A(n_578), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_578), .B(n_707), .Y(n_709) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_580), .A2(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g625 ( .A(n_582), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g653 ( .A(n_585), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g600 ( .A(n_586), .Y(n_600) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g642 ( .A(n_588), .Y(n_642) );
INVx1_ASAP7_75t_L g687 ( .A(n_589), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_605), .C(n_628), .Y(n_591) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_L g654 ( .A(n_594), .Y(n_654) );
AND2x2_ASAP7_75t_L g672 ( .A(n_594), .B(n_613), .Y(n_672) );
OR2x2_ASAP7_75t_L g711 ( .A(n_594), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_595), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g607 ( .A(n_597), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g674 ( .A(n_600), .B(n_611), .Y(n_674) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_603), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g715 ( .A(n_603), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B1(n_613), .B2(n_615), .C(n_617), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_606), .A2(n_629), .B(n_632), .Y(n_628) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx3_ASAP7_75t_L g659 ( .A(n_608), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_608), .B(n_702), .Y(n_701) );
INVxp33_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g620 ( .A(n_616), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_621), .B2(n_624), .Y(n_617) );
INVx2_ASAP7_75t_L g723 ( .A(n_619), .Y(n_723) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g702 ( .A(n_627), .Y(n_702) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_634), .B(n_679), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_652), .C(n_664), .D(n_676), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .B(n_643), .C(n_645), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g675 ( .A(n_638), .Y(n_675) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_640), .A2(n_646), .B(n_649), .Y(n_645) );
INVx2_ASAP7_75t_L g724 ( .A(n_641), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_642), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g657 ( .A(n_642), .Y(n_657) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
OR2x2_ASAP7_75t_L g719 ( .A(n_647), .B(n_683), .Y(n_719) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_654), .Y(n_690) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g660 ( .A(n_656), .B(n_661), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_656), .A2(n_686), .B(n_688), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_656), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g714 ( .A(n_656), .Y(n_714) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp33_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_685), .C(n_695), .D(n_716), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B1(n_692), .B2(n_694), .Y(n_688) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI211xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_699), .B(n_703), .C(n_710), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .B(n_715), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_720), .B(n_722), .Y(n_716) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx3_ASAP7_75t_SL g729 ( .A(n_725), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
CKINVDCx6p67_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_736), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
BUFx8_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
BUFx4f_ASAP7_75t_SL g758 ( .A(n_749), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_750), .B(n_754), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule