module fake_netlist_6_486_n_1044 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1044);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1044;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_114),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_10),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_190),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_86),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_104),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_162),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_24),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_74),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_107),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_79),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_12),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_166),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_93),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_30),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_56),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_31),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_85),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_60),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_160),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_208),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_106),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_21),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_21),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_28),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_13),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_50),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_48),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_65),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_172),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_141),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_92),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_67),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_26),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_218),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_167),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_24),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_153),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_209),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_73),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_28),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_188),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_134),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_33),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_158),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_53),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_195),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_119),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_142),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_165),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_78),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_58),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_170),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_22),
.Y(n_305)
);

BUFx8_ASAP7_75t_SL g306 ( 
.A(n_29),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_31),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_131),
.Y(n_309)
);

BUFx8_ASAP7_75t_SL g310 ( 
.A(n_200),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_59),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_148),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_82),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_133),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_41),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_41),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_137),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_175),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_243),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_254),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_246),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_284),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_252),
.B(n_0),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_257),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_1),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_1),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_264),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_224),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_267),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_224),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_223),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_2),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_229),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_262),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_265),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_270),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_231),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_236),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_236),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_232),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_233),
.Y(n_355)
);

BUFx2_ASAP7_75t_SL g356 ( 
.A(n_229),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_268),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_271),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_290),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_305),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g361 ( 
.A(n_241),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_241),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_310),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_247),
.B(n_2),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_310),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_247),
.B(n_3),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_293),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_300),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_253),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_235),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_307),
.B(n_3),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_237),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_238),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_328),
.B(n_225),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_249),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_356),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_R g384 ( 
.A(n_364),
.B(n_240),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_361),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_226),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_364),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_371),
.B(n_302),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_320),
.B(n_249),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_323),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_227),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_347),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

INVx4_ASAP7_75t_R g405 ( 
.A(n_353),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_332),
.A2(n_286),
.B1(n_312),
.B2(n_230),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_331),
.B(n_276),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_322),
.B(n_276),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_366),
.B(n_242),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_333),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_366),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_374),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_371),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_354),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_355),
.B(n_228),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_348),
.B(n_244),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_239),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_352),
.B(n_248),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_357),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_368),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_358),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_396),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_358),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_392),
.B(n_359),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_359),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_412),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_392),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_379),
.B(n_234),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_360),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_360),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_377),
.B(n_319),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_325),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_315),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_379),
.B(n_258),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_404),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_427),
.B(n_386),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_387),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_406),
.B(n_394),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_234),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_256),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_390),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_407),
.A2(n_292),
.B1(n_281),
.B2(n_260),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_234),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_400),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_259),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_417),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_398),
.B(n_261),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_430),
.B(n_319),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_274),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_411),
.B(n_275),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_403),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_234),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

NAND2x1p5_ASAP7_75t_L g492 ( 
.A(n_420),
.B(n_272),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_408),
.B(n_277),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_382),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_433),
.B(n_368),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_417),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_411),
.B(n_428),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_421),
.B(n_370),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_430),
.B(n_297),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_429),
.B(n_285),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_411),
.B(n_429),
.Y(n_504)
);

INVx4_ASAP7_75t_SL g505 ( 
.A(n_429),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_431),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_278),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_431),
.B(n_263),
.Y(n_509)
);

AO22x1_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_450),
.B1(n_451),
.B2(n_506),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_490),
.A2(n_402),
.B1(n_397),
.B2(n_424),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_445),
.B(n_424),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_445),
.B(n_391),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_380),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_449),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_230),
.B1(n_308),
.B2(n_303),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_437),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_434),
.B(n_380),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_434),
.B(n_385),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_508),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_437),
.B(n_419),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_465),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_436),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_466),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_291),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_493),
.A2(n_418),
.B1(n_385),
.B2(n_389),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_493),
.A2(n_343),
.B1(n_340),
.B2(n_363),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_461),
.B(n_389),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g531 ( 
.A(n_509),
.B(n_297),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_459),
.Y(n_532)
);

OAI22x1_ASAP7_75t_L g533 ( 
.A1(n_508),
.A2(n_370),
.B1(n_432),
.B2(n_418),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_436),
.B(n_432),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_446),
.B(n_296),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_444),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_441),
.B(n_416),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_438),
.B(n_299),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_438),
.B(n_297),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_438),
.B(n_297),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_466),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_449),
.B(n_313),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_484),
.B(n_314),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_495),
.B(n_405),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_492),
.B(n_263),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_485),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_450),
.A2(n_416),
.B1(n_346),
.B2(n_288),
.Y(n_548)
);

AND2x6_ASAP7_75t_SL g549 ( 
.A(n_501),
.B(n_303),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_279),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_488),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_469),
.B(n_280),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_457),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_492),
.A2(n_317),
.B1(n_283),
.B2(n_287),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_485),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_470),
.B(n_289),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_504),
.A2(n_295),
.B(n_294),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_464),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_488),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_470),
.B(n_298),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_464),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_467),
.B(n_384),
.Y(n_563)
);

NAND2x1_ASAP7_75t_L g564 ( 
.A(n_440),
.B(n_47),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_499),
.A2(n_308),
.B1(n_415),
.B2(n_422),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_471),
.B(n_301),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_482),
.B(n_304),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_440),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_457),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_492),
.B(n_263),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_467),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_475),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_480),
.B(n_309),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_467),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_509),
.A2(n_263),
.B1(n_236),
.B2(n_413),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_480),
.B(n_263),
.Y(n_578)
);

AND2x6_ASAP7_75t_SL g579 ( 
.A(n_454),
.B(n_395),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_435),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_477),
.B(n_5),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_505),
.B(n_458),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_505),
.B(n_263),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_486),
.Y(n_586)
);

BUFx4_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_460),
.B(n_458),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_448),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_494),
.B(n_263),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_489),
.B(n_49),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_478),
.B(n_5),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_489),
.B(n_51),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_494),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_522),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_525),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_551),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_545),
.B(n_496),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_515),
.B(n_498),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_571),
.B(n_496),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_460),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_537),
.B(n_505),
.Y(n_602)
);

BUFx4f_ASAP7_75t_L g603 ( 
.A(n_545),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_452),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_553),
.A2(n_460),
.B1(n_503),
.B2(n_462),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_SL g607 ( 
.A(n_577),
.B(n_472),
.C(n_481),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_594),
.B(n_503),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_579),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_538),
.B(n_500),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_592),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_516),
.B(n_505),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_560),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_519),
.B(n_503),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_517),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_516),
.B(n_476),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_519),
.B(n_476),
.Y(n_620)
);

BUFx8_ASAP7_75t_L g621 ( 
.A(n_563),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_517),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_573),
.B(n_439),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_528),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_580),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_512),
.B(n_476),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_547),
.B(n_479),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_513),
.Y(n_628)
);

NAND2x1p5_ASAP7_75t_L g629 ( 
.A(n_534),
.B(n_593),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_587),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_SL g631 ( 
.A(n_581),
.B(n_439),
.C(n_448),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_576),
.Y(n_634)
);

BUFx4f_ASAP7_75t_L g635 ( 
.A(n_547),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_548),
.Y(n_636)
);

AOI221xp5_ASAP7_75t_SL g637 ( 
.A1(n_524),
.A2(n_566),
.B1(n_526),
.B2(n_542),
.C(n_589),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_582),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_511),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_517),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_547),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_547),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_555),
.B(n_486),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_569),
.B(n_458),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_569),
.B(n_458),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_518),
.B(n_443),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

AOI22x1_ASAP7_75t_L g649 ( 
.A1(n_583),
.A2(n_440),
.B1(n_455),
.B2(n_491),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_514),
.B(n_458),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_593),
.B(n_491),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_531),
.A2(n_502),
.B1(n_447),
.B2(n_487),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_533),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_518),
.B(n_474),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_SL g655 ( 
.A(n_581),
.B(n_521),
.C(n_520),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_SL g656 ( 
.A(n_577),
.B(n_455),
.C(n_443),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_510),
.B(n_474),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_556),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_555),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_628),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_607),
.A2(n_550),
.B(n_552),
.C(n_531),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_596),
.B(n_529),
.Y(n_663)
);

AO31x2_ASAP7_75t_L g664 ( 
.A1(n_657),
.A2(n_539),
.A3(n_578),
.B(n_527),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_649),
.A2(n_588),
.B(n_584),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_600),
.B(n_550),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_645),
.A2(n_534),
.B(n_463),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_601),
.B(n_626),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_607),
.A2(n_552),
.B(n_590),
.C(n_543),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_638),
.B(n_650),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_627),
.A2(n_584),
.B(n_536),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_629),
.B(n_591),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_620),
.B(n_555),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_616),
.B(n_555),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_647),
.A2(n_591),
.B1(n_529),
.B2(n_544),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_651),
.B(n_523),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_643),
.A2(n_564),
.B(n_562),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_656),
.A2(n_572),
.B(n_546),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_618),
.B(n_623),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_646),
.A2(n_463),
.B(n_497),
.Y(n_680)
);

AO31x2_ASAP7_75t_L g681 ( 
.A1(n_657),
.A2(n_599),
.A3(n_554),
.B(n_604),
.Y(n_681)
);

OAI21x1_ASAP7_75t_SL g682 ( 
.A1(n_648),
.A2(n_561),
.B(n_557),
.Y(n_682)
);

AO21x1_ASAP7_75t_L g683 ( 
.A1(n_613),
.A2(n_541),
.B(n_540),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_643),
.A2(n_567),
.B(n_559),
.Y(n_684)
);

AO22x2_ASAP7_75t_L g685 ( 
.A1(n_654),
.A2(n_549),
.B1(n_521),
.B2(n_520),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_595),
.Y(n_686)
);

AO21x2_ASAP7_75t_L g687 ( 
.A1(n_655),
.A2(n_585),
.B(n_541),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_635),
.A2(n_463),
.B(n_497),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_599),
.A2(n_575),
.B(n_568),
.C(n_530),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_635),
.A2(n_619),
.B(n_629),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_SL g691 ( 
.A(n_655),
.B(n_540),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_651),
.B(n_574),
.Y(n_692)
);

AOI221x1_ASAP7_75t_L g693 ( 
.A1(n_656),
.A2(n_558),
.B1(n_483),
.B2(n_474),
.C(n_586),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_637),
.A2(n_585),
.B(n_447),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_644),
.A2(n_453),
.B(n_474),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_622),
.B(n_660),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_651),
.B(n_474),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_602),
.A2(n_456),
.B(n_447),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_652),
.A2(n_606),
.B1(n_631),
.B2(n_624),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_651),
.B(n_632),
.Y(n_700)
);

AOI221x1_ASAP7_75t_L g701 ( 
.A1(n_614),
.A2(n_456),
.B1(n_502),
.B2(n_473),
.C(n_468),
.Y(n_701)
);

AOI21xp33_ASAP7_75t_L g702 ( 
.A1(n_612),
.A2(n_6),
.B(n_7),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_597),
.A2(n_615),
.B(n_617),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_623),
.A2(n_447),
.B1(n_502),
.B2(n_473),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_617),
.A2(n_640),
.B(n_658),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_644),
.A2(n_453),
.B(n_447),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_632),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_631),
.A2(n_502),
.B(n_487),
.C(n_473),
.Y(n_708)
);

NOR2x1_ASAP7_75t_SL g709 ( 
.A(n_622),
.B(n_453),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_640),
.A2(n_447),
.B(n_468),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_608),
.A2(n_502),
.B(n_473),
.Y(n_711)
);

AOI221xp5_ASAP7_75t_L g712 ( 
.A1(n_605),
.A2(n_636),
.B1(n_639),
.B2(n_653),
.C(n_611),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_659),
.A2(n_502),
.A3(n_487),
.B(n_473),
.Y(n_713)
);

AOI21xp33_ASAP7_75t_L g714 ( 
.A1(n_634),
.A2(n_6),
.B(n_7),
.Y(n_714)
);

AOI221x1_ASAP7_75t_L g715 ( 
.A1(n_622),
.A2(n_487),
.B1(n_473),
.B2(n_468),
.C(n_11),
.Y(n_715)
);

AOI21x1_ASAP7_75t_L g716 ( 
.A1(n_642),
.A2(n_453),
.B(n_468),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_618),
.B(n_453),
.Y(n_717)
);

AO21x2_ASAP7_75t_L g718 ( 
.A1(n_662),
.A2(n_610),
.B(n_642),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_665),
.A2(n_652),
.B(n_634),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_684),
.A2(n_651),
.B(n_622),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_696),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_668),
.B(n_641),
.Y(n_723)
);

AO21x2_ASAP7_75t_L g724 ( 
.A1(n_678),
.A2(n_610),
.B(n_487),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_705),
.A2(n_660),
.B(n_633),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_686),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_703),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_677),
.A2(n_671),
.B(n_678),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_707),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_699),
.A2(n_625),
.B1(n_621),
.B2(n_598),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_679),
.B(n_690),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_663),
.A2(n_609),
.B1(n_603),
.B2(n_598),
.Y(n_732)
);

OA21x2_ASAP7_75t_L g733 ( 
.A1(n_693),
.A2(n_487),
.B(n_468),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_698),
.B(n_660),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_666),
.A2(n_699),
.B1(n_675),
.B2(n_670),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_669),
.A2(n_660),
.B(n_633),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_680),
.A2(n_633),
.B(n_598),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_673),
.B(n_621),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_675),
.A2(n_603),
.B1(n_468),
.B2(n_630),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_692),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_SL g741 ( 
.A1(n_689),
.A2(n_717),
.B(n_676),
.C(n_694),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_694),
.A2(n_54),
.B(n_52),
.Y(n_742)
);

OAI21xp5_ASAP7_75t_L g743 ( 
.A1(n_674),
.A2(n_57),
.B(n_55),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_696),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_712),
.B(n_8),
.Y(n_745)
);

AO21x2_ASAP7_75t_L g746 ( 
.A1(n_683),
.A2(n_62),
.B(n_61),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_700),
.Y(n_747)
);

OA21x2_ASAP7_75t_L g748 ( 
.A1(n_701),
.A2(n_8),
.B(n_9),
.Y(n_748)
);

BUFx12f_ASAP7_75t_L g749 ( 
.A(n_702),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_697),
.B(n_63),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_710),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_681),
.B(n_10),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_714),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_17),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_667),
.A2(n_124),
.B(n_220),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_691),
.A2(n_123),
.B(n_217),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_681),
.Y(n_757)
);

OR2x4_ASAP7_75t_L g758 ( 
.A(n_685),
.B(n_14),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_687),
.B(n_15),
.Y(n_759)
);

OA21x2_ASAP7_75t_L g760 ( 
.A1(n_711),
.A2(n_16),
.B(n_18),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_681),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_711),
.A2(n_18),
.B(n_19),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_664),
.B(n_19),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_709),
.B(n_64),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_687),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_716),
.A2(n_127),
.B(n_216),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_695),
.B(n_66),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_685),
.Y(n_768)
);

OAI21x1_ASAP7_75t_L g769 ( 
.A1(n_688),
.A2(n_126),
.B(n_215),
.Y(n_769)
);

AO21x1_ASAP7_75t_L g770 ( 
.A1(n_672),
.A2(n_20),
.B(n_23),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_706),
.A2(n_125),
.B(n_214),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_719),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_723),
.B(n_664),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_SL g774 ( 
.A1(n_745),
.A2(n_715),
.B(n_708),
.Y(n_774)
);

AOI222xp33_ASAP7_75t_L g775 ( 
.A1(n_749),
.A2(n_672),
.B1(n_23),
.B2(n_25),
.C1(n_26),
.C2(n_27),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_719),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_SL g777 ( 
.A(n_730),
.B(n_756),
.C(n_770),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_723),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_729),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_726),
.B(n_664),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_747),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_763),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_749),
.A2(n_704),
.B1(n_713),
.B2(n_27),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_758),
.A2(n_20),
.B1(n_25),
.B2(n_29),
.Y(n_784)
);

NAND3xp33_ASAP7_75t_SL g785 ( 
.A(n_770),
.B(n_30),
.C(n_32),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_763),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_740),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_R g788 ( 
.A(n_738),
.B(n_68),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_735),
.A2(n_713),
.B1(n_33),
.B2(n_34),
.Y(n_789)
);

BUFx12f_ASAP7_75t_L g790 ( 
.A(n_753),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_722),
.Y(n_791)
);

BUFx2_ASAP7_75t_SL g792 ( 
.A(n_722),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_758),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_740),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_747),
.B(n_713),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_722),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_741),
.A2(n_136),
.B(n_212),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_732),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_758),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_753),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_768),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_739),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_722),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_731),
.B(n_718),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_752),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_752),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_722),
.Y(n_807)
);

BUFx4f_ASAP7_75t_SL g808 ( 
.A(n_744),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_731),
.B(n_42),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_754),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_757),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_731),
.B(n_44),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_718),
.B(n_45),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_743),
.A2(n_46),
.B1(n_70),
.B2(n_71),
.Y(n_814)
);

OAI222xp33_ASAP7_75t_L g815 ( 
.A1(n_757),
.A2(n_46),
.B1(n_72),
.B2(n_75),
.C1(n_76),
.C2(n_77),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_761),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_SL g817 ( 
.A1(n_760),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_764),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_750),
.A2(n_84),
.B1(n_87),
.B2(n_90),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_744),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_744),
.Y(n_821)
);

OAI221xp5_ASAP7_75t_L g822 ( 
.A1(n_759),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.C(n_96),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_718),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_750),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_764),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_761),
.B(n_750),
.Y(n_826)
);

OAI221xp5_ASAP7_75t_L g827 ( 
.A1(n_760),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.C(n_105),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_720),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_764),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_736),
.A2(n_108),
.B(n_109),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_796),
.Y(n_831)
);

BUFx4f_ASAP7_75t_SL g832 ( 
.A(n_803),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_782),
.B(n_765),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_793),
.A2(n_760),
.B1(n_762),
.B2(n_767),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_787),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_830),
.A2(n_728),
.B(n_755),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_780),
.B(n_765),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_798),
.A2(n_767),
.B1(n_760),
.B2(n_762),
.C(n_734),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_775),
.A2(n_762),
.B1(n_767),
.B2(n_746),
.Y(n_839)
);

OR2x6_ASAP7_75t_SL g840 ( 
.A(n_813),
.B(n_727),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_794),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_830),
.A2(n_728),
.B(n_755),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_775),
.A2(n_762),
.B1(n_746),
.B2(n_724),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_SL g844 ( 
.A1(n_793),
.A2(n_734),
.B1(n_727),
.B2(n_751),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_814),
.A2(n_769),
.B(n_748),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_800),
.B(n_748),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_777),
.A2(n_737),
.B1(n_746),
.B2(n_724),
.Y(n_847)
);

OAI211xp5_ASAP7_75t_L g848 ( 
.A1(n_801),
.A2(n_748),
.B(n_769),
.C(n_742),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_786),
.B(n_724),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_772),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_776),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_778),
.B(n_748),
.Y(n_852)
);

AO221x1_ASAP7_75t_L g853 ( 
.A1(n_799),
.A2(n_784),
.B1(n_815),
.B2(n_810),
.C(n_802),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_829),
.A2(n_734),
.B1(n_751),
.B2(n_733),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_805),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_788),
.A2(n_733),
.B1(n_742),
.B2(n_737),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_789),
.A2(n_733),
.B1(n_720),
.B2(n_771),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_828),
.A2(n_721),
.B(n_771),
.Y(n_858)
);

OAI21xp33_ASAP7_75t_L g859 ( 
.A1(n_799),
.A2(n_785),
.B(n_802),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_SL g860 ( 
.A1(n_822),
.A2(n_733),
.B1(n_766),
.B2(n_725),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_790),
.A2(n_766),
.B1(n_721),
.B2(n_725),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_822),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_779),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_811),
.Y(n_864)
);

AOI221xp5_ASAP7_75t_L g865 ( 
.A1(n_827),
.A2(n_813),
.B1(n_774),
.B2(n_783),
.C(n_797),
.Y(n_865)
);

AOI222xp33_ASAP7_75t_L g866 ( 
.A1(n_827),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.C1(n_121),
.C2(n_122),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_812),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_867)
);

OAI221xp5_ASAP7_75t_L g868 ( 
.A1(n_824),
.A2(n_132),
.B1(n_135),
.B2(n_140),
.C(n_143),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_819),
.A2(n_144),
.B(n_145),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_773),
.B(n_221),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_808),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_809),
.B(n_151),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_817),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_825),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_874)
);

AOI222xp33_ASAP7_75t_L g875 ( 
.A1(n_781),
.A2(n_163),
.B1(n_164),
.B2(n_168),
.C1(n_169),
.C2(n_174),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_796),
.Y(n_876)
);

OAI221xp5_ASAP7_75t_L g877 ( 
.A1(n_804),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.C(n_180),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_825),
.B(n_182),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_863),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_840),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_849),
.B(n_804),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_833),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_855),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_837),
.B(n_823),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_855),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_837),
.B(n_816),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_864),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_864),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_850),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_850),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_840),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_835),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_865),
.A2(n_795),
.B(n_806),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_846),
.B(n_826),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_833),
.Y(n_895)
);

AOI221xp5_ASAP7_75t_L g896 ( 
.A1(n_859),
.A2(n_825),
.B1(n_795),
.B2(n_820),
.C(n_791),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_835),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_841),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_846),
.B(n_807),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_852),
.B(n_807),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_852),
.B(n_818),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_851),
.B(n_818),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_841),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_858),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_831),
.Y(n_906)
);

AO31x2_ASAP7_75t_L g907 ( 
.A1(n_845),
.A2(n_821),
.A3(n_792),
.B(n_796),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_870),
.B(n_821),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_870),
.B(n_847),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_838),
.A2(n_183),
.B(n_184),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_843),
.B(n_185),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_839),
.A2(n_187),
.B1(n_189),
.B2(n_191),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_858),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_R g914 ( 
.A(n_908),
.B(n_832),
.Y(n_914)
);

OAI211xp5_ASAP7_75t_L g915 ( 
.A1(n_910),
.A2(n_866),
.B(n_834),
.C(n_875),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_883),
.Y(n_916)
);

AND2x2_ASAP7_75t_SL g917 ( 
.A(n_880),
.B(n_862),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_880),
.B(n_854),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_910),
.A2(n_869),
.B(n_877),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_879),
.Y(n_920)
);

AOI33xp33_ASAP7_75t_L g921 ( 
.A1(n_879),
.A2(n_873),
.A3(n_856),
.B1(n_853),
.B2(n_867),
.B3(n_874),
.Y(n_921)
);

NAND4xp25_ASAP7_75t_SL g922 ( 
.A(n_896),
.B(n_868),
.C(n_848),
.D(n_853),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_911),
.B(n_878),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_891),
.B(n_836),
.Y(n_924)
);

NOR2x1_ASAP7_75t_SL g925 ( 
.A(n_909),
.B(n_887),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_883),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_908),
.B(n_876),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_887),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_883),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_895),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_889),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_912),
.A2(n_872),
.B(n_871),
.C(n_836),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_911),
.A2(n_844),
.B1(n_860),
.B2(n_857),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_888),
.Y(n_934)
);

AO21x2_ASAP7_75t_L g935 ( 
.A1(n_905),
.A2(n_842),
.B(n_861),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_925),
.B(n_891),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_930),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_918),
.B(n_920),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_931),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_916),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_916),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_926),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_926),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_918),
.B(n_894),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_929),
.B(n_894),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_929),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_928),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_899),
.Y(n_948)
);

INVx5_ASAP7_75t_SL g949 ( 
.A(n_935),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_934),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_936),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_947),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_939),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_936),
.B(n_924),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_938),
.B(n_922),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_944),
.B(n_927),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_948),
.B(n_899),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_947),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_956),
.B(n_944),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_955),
.B(n_938),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_951),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_951),
.A2(n_919),
.B(n_915),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_956),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_954),
.B(n_945),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_953),
.B(n_937),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_957),
.Y(n_966)
);

NAND2x1p5_ASAP7_75t_L g967 ( 
.A(n_953),
.B(n_939),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_961),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_966),
.Y(n_969)
);

AOI222xp33_ASAP7_75t_L g970 ( 
.A1(n_962),
.A2(n_917),
.B1(n_923),
.B2(n_933),
.C1(n_909),
.C2(n_912),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_961),
.Y(n_971)
);

OAI32xp33_ASAP7_75t_L g972 ( 
.A1(n_962),
.A2(n_953),
.A3(n_957),
.B1(n_948),
.B2(n_954),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_970),
.A2(n_963),
.B1(n_917),
.B2(n_969),
.Y(n_973)
);

OAI22xp33_ASAP7_75t_SL g974 ( 
.A1(n_968),
.A2(n_967),
.B1(n_960),
.B2(n_965),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_971),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_972),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_975),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_L g978 ( 
.A1(n_976),
.A2(n_967),
.B1(n_972),
.B2(n_939),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_973),
.B(n_959),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_974),
.B(n_964),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_975),
.Y(n_981)
);

AOI221xp5_ASAP7_75t_L g982 ( 
.A1(n_978),
.A2(n_932),
.B1(n_958),
.B2(n_952),
.C(n_896),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_979),
.A2(n_932),
.B(n_893),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_980),
.B(n_939),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_977),
.A2(n_893),
.B(n_950),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_981),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_921),
.C(n_906),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_977),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_977),
.B(n_950),
.Y(n_989)
);

OAI211xp5_ASAP7_75t_SL g990 ( 
.A1(n_986),
.A2(n_921),
.B(n_943),
.C(n_941),
.Y(n_990)
);

BUFx4f_ASAP7_75t_SL g991 ( 
.A(n_988),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_989),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_983),
.A2(n_949),
.B1(n_943),
.B2(n_941),
.Y(n_993)
);

AOI322xp5_ASAP7_75t_L g994 ( 
.A1(n_987),
.A2(n_949),
.A3(n_945),
.B1(n_902),
.B2(n_923),
.C1(n_886),
.C2(n_900),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_984),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_982),
.A2(n_949),
.B1(n_923),
.B2(n_903),
.Y(n_996)
);

OAI221xp5_ASAP7_75t_L g997 ( 
.A1(n_985),
.A2(n_906),
.B1(n_946),
.B2(n_942),
.C(n_940),
.Y(n_997)
);

AOI211x1_ASAP7_75t_L g998 ( 
.A1(n_995),
.A2(n_949),
.B(n_903),
.C(n_888),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_991),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_992),
.B(n_946),
.Y(n_1000)
);

AOI31xp33_ASAP7_75t_L g1001 ( 
.A1(n_996),
.A2(n_914),
.A3(n_882),
.B(n_902),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_990),
.A2(n_949),
.B1(n_923),
.B2(n_906),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_997),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_993),
.B(n_906),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_994),
.Y(n_1005)
);

AOI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_995),
.A2(n_935),
.B(n_876),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_942),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1005),
.B(n_1003),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_L g1009 ( 
.A(n_1001),
.B(n_1004),
.C(n_1006),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_1000),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_998),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1002),
.Y(n_1012)
);

NAND3x1_ASAP7_75t_L g1013 ( 
.A(n_1003),
.B(n_900),
.C(n_886),
.Y(n_1013)
);

NOR3x1_ASAP7_75t_L g1014 ( 
.A(n_1005),
.B(n_904),
.C(n_905),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_1000),
.B(n_831),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_1010),
.Y(n_1016)
);

OR3x1_ASAP7_75t_L g1017 ( 
.A(n_1012),
.B(n_913),
.C(n_897),
.Y(n_1017)
);

AO22x2_ASAP7_75t_L g1018 ( 
.A1(n_1008),
.A2(n_940),
.B1(n_831),
.B2(n_913),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_1009),
.B(n_842),
.C(n_892),
.Y(n_1019)
);

OAI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1011),
.A2(n_890),
.B1(n_897),
.B2(n_889),
.C(n_898),
.Y(n_1020)
);

XNOR2xp5_ASAP7_75t_L g1021 ( 
.A(n_1007),
.B(n_192),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1013),
.A2(n_923),
.B1(n_935),
.B2(n_931),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_892),
.C(n_898),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_SL g1024 ( 
.A(n_1014),
.B(n_904),
.C(n_890),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1016),
.Y(n_1025)
);

NAND3xp33_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_895),
.C(n_885),
.Y(n_1026)
);

XNOR2xp5_ASAP7_75t_L g1027 ( 
.A(n_1021),
.B(n_193),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1018),
.B(n_901),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_1020),
.A2(n_923),
.B(n_881),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1025),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1027),
.B(n_1018),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1026),
.A2(n_1022),
.B1(n_1017),
.B2(n_1023),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1028),
.Y(n_1033)
);

XNOR2xp5_ASAP7_75t_L g1034 ( 
.A(n_1030),
.B(n_1024),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1033),
.A2(n_1029),
.B1(n_931),
.B2(n_885),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_1034),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1035),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_L g1038 ( 
.A(n_1036),
.B(n_1031),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_1037),
.A2(n_1032),
.B(n_196),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_SL g1040 ( 
.A1(n_1038),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_1039),
.Y(n_1041)
);

AOI322xp5_ASAP7_75t_L g1042 ( 
.A1(n_1041),
.A2(n_1040),
.A3(n_901),
.B1(n_885),
.B2(n_884),
.C1(n_907),
.C2(n_206),
.Y(n_1042)
);

OAI221xp5_ASAP7_75t_R g1043 ( 
.A1(n_1042),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1043),
.A2(n_205),
.B(n_210),
.C(n_211),
.Y(n_1044)
);


endmodule