module real_aes_16778_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_82;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_0), .A2(n_2), .B1(n_120), .B2(n_121), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g88 ( .A1(n_1), .A2(n_16), .B1(n_89), .B2(n_91), .Y(n_88) );
AND2x2_ASAP7_75t_L g505 ( .A(n_3), .B(n_69), .Y(n_505) );
AND2x2_ASAP7_75t_L g568 ( .A(n_3), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g592 ( .A(n_3), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_4), .A2(n_43), .B1(n_179), .B2(n_188), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_5), .A2(n_9), .B1(n_96), .B2(n_171), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_6), .Y(n_142) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_7), .Y(n_90) );
INVx1_ASAP7_75t_L g458 ( .A(n_8), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_10), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_10), .Y(n_457) );
INVx1_ASAP7_75t_L g480 ( .A(n_11), .Y(n_480) );
INVx1_ASAP7_75t_L g497 ( .A(n_11), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_12), .A2(n_67), .B1(n_541), .B2(n_546), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_12), .A2(n_47), .B1(n_603), .B2(n_607), .C(n_608), .Y(n_602) );
INVx2_ASAP7_75t_L g483 ( .A(n_13), .Y(n_483) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_14), .A2(n_40), .B(n_105), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
INVx4_ASAP7_75t_R g207 ( .A(n_17), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_18), .B(n_94), .Y(n_149) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_19), .A2(n_31), .B1(n_538), .B2(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_19), .A2(n_41), .B1(n_594), .B2(n_596), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_20), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_21), .Y(n_570) );
INVx1_ASAP7_75t_L g128 ( .A(n_22), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_23), .B(n_91), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_SL g140 ( .A1(n_24), .A2(n_93), .B(n_96), .C(n_141), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g95 ( .A1(n_25), .A2(n_37), .B1(n_96), .B2(n_97), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_26), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_27), .Y(n_137) );
INVx1_ASAP7_75t_L g464 ( .A(n_28), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_29), .A2(n_41), .B1(n_535), .B2(n_538), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_29), .A2(n_31), .B1(n_582), .B2(n_587), .C(n_589), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_30), .Y(n_511) );
INVx2_ASAP7_75t_L g485 ( .A(n_32), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_32), .B(n_483), .Y(n_500) );
INVx1_ASAP7_75t_L g555 ( .A(n_32), .Y(n_555) );
INVx1_ASAP7_75t_L g154 ( .A(n_33), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_34), .B(n_96), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_35), .Y(n_172) );
INVx2_ASAP7_75t_L g641 ( .A(n_36), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_38), .A2(n_70), .B1(n_96), .B2(n_97), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_39), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_42), .Y(n_565) );
BUFx3_ASAP7_75t_L g477 ( .A(n_44), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_45), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_46), .A2(n_47), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_46), .A2(n_67), .B1(n_594), .B2(n_596), .Y(n_593) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_48), .A2(n_622), .B(n_631), .Y(n_621) );
INVx1_ASAP7_75t_L g105 ( .A(n_49), .Y(n_105) );
AND2x4_ASAP7_75t_L g107 ( .A(n_50), .B(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_50), .Y(n_651) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_51), .Y(n_510) );
BUFx3_ASAP7_75t_L g463 ( .A(n_52), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_53), .A2(n_72), .B1(n_97), .B2(n_117), .Y(n_116) );
AO22x1_ASAP7_75t_L g192 ( .A1(n_54), .A2(n_61), .B1(n_150), .B2(n_193), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_54), .A2(n_461), .B1(n_462), .B2(n_467), .Y(n_460) );
INVx1_ASAP7_75t_L g467 ( .A(n_54), .Y(n_467) );
INVx1_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
AND2x2_ASAP7_75t_L g144 ( .A(n_56), .B(n_102), .Y(n_144) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_57), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_58), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_59), .B(n_179), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_60), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_62), .B(n_91), .Y(n_173) );
INVx2_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_64), .A2(n_468), .B1(n_469), .B2(n_653), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_64), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_65), .B(n_102), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_66), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_68), .B(n_112), .Y(n_190) );
INVx1_ASAP7_75t_L g569 ( .A(n_69), .Y(n_569) );
BUFx3_ASAP7_75t_L g591 ( .A(n_69), .Y(n_591) );
INVx1_ASAP7_75t_L g489 ( .A(n_71), .Y(n_489) );
INVx1_ASAP7_75t_L g503 ( .A(n_71), .Y(n_503) );
INVx2_ASAP7_75t_L g533 ( .A(n_71), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_73), .B(n_102), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_74), .A2(n_124), .B(n_179), .C(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g212 ( .A(n_75), .B(n_213), .Y(n_212) );
NAND2xp33_ASAP7_75t_L g177 ( .A(n_76), .B(n_118), .Y(n_177) );
AOI21xp33_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_444), .B(n_452), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x4_ASAP7_75t_L g79 ( .A(n_80), .B(n_336), .Y(n_79) );
NOR2xp67_ASAP7_75t_L g80 ( .A(n_81), .B(n_278), .Y(n_80) );
NAND3xp33_ASAP7_75t_SL g81 ( .A(n_82), .B(n_214), .C(n_260), .Y(n_81) );
OAI21xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_159), .B(n_182), .Y(n_82) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_83), .A2(n_215), .B1(n_234), .B2(n_247), .Y(n_214) );
AOI22x1_ASAP7_75t_L g340 ( .A1(n_83), .A2(n_341), .B1(n_345), .B2(n_346), .Y(n_340) );
INVx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
OR2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_129), .Y(n_84) );
OR2x2_ASAP7_75t_L g301 ( .A(n_85), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_86), .B(n_113), .Y(n_85) );
OR2x2_ASAP7_75t_L g164 ( .A(n_86), .B(n_113), .Y(n_164) );
AND2x2_ASAP7_75t_L g218 ( .A(n_86), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_SL g226 ( .A(n_86), .Y(n_226) );
BUFx2_ASAP7_75t_L g277 ( .A(n_86), .Y(n_277) );
AO31x2_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_101), .A3(n_106), .B(n_109), .Y(n_86) );
OAI22xp5_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_92), .B1(n_95), .B2(n_98), .Y(n_87) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_89), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
INVx3_ASAP7_75t_L g96 ( .A(n_90), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_90), .Y(n_97) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
INVx1_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
INVx1_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx1_ASAP7_75t_L g179 ( .A(n_90), .Y(n_179) );
INVx1_ASAP7_75t_L g189 ( .A(n_90), .Y(n_189) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_90), .Y(n_194) );
INVx1_ASAP7_75t_L g208 ( .A(n_90), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_91), .B(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_92), .A2(n_116), .B1(n_119), .B2(n_123), .Y(n_115) );
OAI22x1_ASAP7_75t_L g241 ( .A1(n_92), .A2(n_123), .B1(n_242), .B2(n_243), .Y(n_241) );
INVx6_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_93), .A2(n_177), .B(n_178), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_93), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_93), .A2(n_186), .B(n_192), .C(n_196), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_93), .B(n_449), .Y(n_448) );
BUFx8_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g100 ( .A(n_94), .Y(n_100) );
INVx1_ASAP7_75t_L g124 ( .A(n_94), .Y(n_124) );
INVx1_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
INVx4_ASAP7_75t_L g171 ( .A(n_96), .Y(n_171) );
INVx2_ASAP7_75t_L g120 ( .A(n_97), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_97), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_98), .A2(n_156), .B(n_157), .Y(n_155) );
OAI21x1_ASAP7_75t_L g186 ( .A1(n_98), .A2(n_187), .B(n_190), .Y(n_186) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g175 ( .A(n_100), .Y(n_175) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NOR2x1_ASAP7_75t_L g180 ( .A(n_102), .B(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g158 ( .A(n_103), .B(n_106), .Y(n_158) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g112 ( .A(n_104), .Y(n_112) );
INVx1_ASAP7_75t_L g181 ( .A(n_106), .Y(n_181) );
BUFx10_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g126 ( .A(n_107), .Y(n_126) );
INVx1_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
BUFx10_ASAP7_75t_L g211 ( .A(n_107), .Y(n_211) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_108), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
BUFx2_ASAP7_75t_L g114 ( .A(n_111), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_111), .B(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g213 ( .A(n_111), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_111), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI21xp33_ASAP7_75t_L g196 ( .A1(n_112), .A2(n_143), .B(n_190), .Y(n_196) );
INVx2_ASAP7_75t_L g200 ( .A(n_112), .Y(n_200) );
INVx2_ASAP7_75t_L g244 ( .A(n_112), .Y(n_244) );
AND2x2_ASAP7_75t_L g221 ( .A(n_113), .B(n_145), .Y(n_221) );
INVx1_ASAP7_75t_L g228 ( .A(n_113), .Y(n_228) );
INVx1_ASAP7_75t_L g233 ( .A(n_113), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_113), .B(n_226), .Y(n_296) );
INVx1_ASAP7_75t_L g317 ( .A(n_113), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_113), .B(n_219), .Y(n_387) );
AO31x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_115), .A3(n_125), .B(n_127), .Y(n_113) );
AOI21x1_ASAP7_75t_L g131 ( .A1(n_114), .A2(n_132), .B(n_144), .Y(n_131) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp33_ASAP7_75t_L g206 ( .A1(n_118), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_206) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_122), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_123), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g280 ( .A(n_129), .Y(n_280) );
OR2x2_ASAP7_75t_L g332 ( .A(n_129), .B(n_296), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_145), .Y(n_129) );
AND2x2_ASAP7_75t_L g165 ( .A(n_130), .B(n_166), .Y(n_165) );
OR2x2_ASAP7_75t_L g224 ( .A(n_130), .B(n_225), .Y(n_224) );
INVxp67_ASAP7_75t_L g230 ( .A(n_130), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_130), .B(n_162), .Y(n_308) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_143), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_136), .B(n_138), .Y(n_133) );
BUFx4f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_139), .B(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g162 ( .A(n_145), .Y(n_162) );
INVx1_ASAP7_75t_L g274 ( .A(n_145), .Y(n_274) );
AND2x2_ASAP7_75t_L g276 ( .A(n_145), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g294 ( .A(n_145), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g316 ( .A(n_145), .B(n_317), .Y(n_316) );
NAND2x1p5_ASAP7_75t_SL g327 ( .A(n_145), .B(n_303), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_145), .B(n_233), .Y(n_417) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_155), .B(n_158), .Y(n_147) );
OAI21xp33_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_150), .B(n_152), .Y(n_148) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_165), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_160), .A2(n_356), .B1(n_357), .B2(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_161), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_161), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g434 ( .A(n_161), .B(n_292), .Y(n_434) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g232 ( .A(n_162), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_162), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g322 ( .A(n_162), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g273 ( .A(n_163), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g363 ( .A(n_164), .Y(n_363) );
OR2x2_ASAP7_75t_L g437 ( .A(n_164), .B(n_364), .Y(n_437) );
INVx1_ASAP7_75t_L g268 ( .A(n_165), .Y(n_268) );
INVx3_ASAP7_75t_L g272 ( .A(n_166), .Y(n_272) );
BUFx2_ASAP7_75t_L g283 ( .A(n_166), .Y(n_283) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g253 ( .A(n_167), .B(n_197), .Y(n_253) );
INVx2_ASAP7_75t_L g299 ( .A(n_167), .Y(n_299) );
INVx1_ASAP7_75t_L g331 ( .A(n_167), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_167), .B(n_240), .Y(n_344) );
AND2x2_ASAP7_75t_L g366 ( .A(n_167), .B(n_265), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_176), .B(n_180), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_174), .Y(n_170) );
INVx2_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g357 ( .A(n_183), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_183), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g382 ( .A(n_183), .B(n_250), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_183), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_197), .Y(n_183) );
INVx2_ASAP7_75t_L g238 ( .A(n_184), .Y(n_238) );
AND2x2_ASAP7_75t_L g266 ( .A(n_184), .B(n_267), .Y(n_266) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_191), .B(n_195), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g451 ( .A(n_188), .Y(n_451) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_189), .B(n_204), .Y(n_203) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g239 ( .A(n_197), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g259 ( .A(n_197), .Y(n_259) );
INVx2_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
OR2x2_ASAP7_75t_L g287 ( .A(n_197), .B(n_240), .Y(n_287) );
AND2x2_ASAP7_75t_L g298 ( .A(n_197), .B(n_299), .Y(n_298) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_201), .B(n_212), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_205), .B(n_210), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_207), .A2(n_468), .B1(n_469), .B2(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_207), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_209), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_210), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_211), .A2(n_241), .A3(n_244), .B(n_245), .Y(n_240) );
OAI221xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B1(n_222), .B2(n_227), .C(n_229), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OAI32xp33_ASAP7_75t_L g328 ( .A1(n_217), .A2(n_231), .A3(n_329), .B1(n_332), .B2(n_333), .Y(n_328) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g318 ( .A(n_218), .Y(n_318) );
AND2x2_ASAP7_75t_L g354 ( .A(n_218), .B(n_232), .Y(n_354) );
INVx1_ASAP7_75t_L g418 ( .A(n_218), .Y(n_418) );
OR2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_226), .Y(n_292) );
INVx2_ASAP7_75t_L g303 ( .A(n_219), .Y(n_303) );
BUFx2_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g442 ( .A(n_221), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVxp67_ASAP7_75t_L g429 ( .A(n_224), .Y(n_429) );
INVx1_ASAP7_75t_L g443 ( .A(n_224), .Y(n_443) );
OR2x2_ASAP7_75t_L g323 ( .A(n_225), .B(n_303), .Y(n_323) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_227), .B(n_323), .Y(n_345) );
INVx1_ASAP7_75t_L g376 ( .A(n_227), .Y(n_376) );
BUFx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g410 ( .A(n_228), .Y(n_410) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2x1_ASAP7_75t_L g379 ( .A(n_230), .B(n_380), .Y(n_379) );
OAI21xp5_ASAP7_75t_SL g401 ( .A1(n_231), .A2(n_402), .B(n_407), .Y(n_401) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_239), .Y(n_235) );
AND2x2_ASAP7_75t_L g311 ( .A(n_236), .B(n_253), .Y(n_311) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_236), .Y(n_441) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g343 ( .A(n_237), .Y(n_343) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g325 ( .A(n_238), .B(n_299), .Y(n_325) );
AND2x2_ASAP7_75t_L g396 ( .A(n_238), .B(n_267), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_239), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g324 ( .A(n_239), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g403 ( .A(n_239), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g252 ( .A(n_240), .Y(n_252) );
INVx2_ASAP7_75t_L g265 ( .A(n_240), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_240), .B(n_256), .Y(n_313) );
AND2x2_ASAP7_75t_L g373 ( .A(n_240), .B(n_267), .Y(n_373) );
NAND2xp33_ASAP7_75t_SL g247 ( .A(n_248), .B(n_254), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g348 ( .A(n_251), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_251), .B(n_331), .Y(n_423) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g255 ( .A(n_252), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g384 ( .A(n_252), .B(n_299), .Y(n_384) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
OR2x2_ASAP7_75t_L g329 ( .A(n_255), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g312 ( .A(n_259), .B(n_313), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_273), .B1(n_275), .B2(n_276), .Y(n_260) );
OAI21xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_268), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g275 ( .A(n_263), .B(n_272), .Y(n_275) );
BUFx2_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g304 ( .A(n_264), .Y(n_304) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g319 ( .A(n_266), .B(n_283), .Y(n_319) );
INVx2_ASAP7_75t_L g335 ( .A(n_266), .Y(n_335) );
AND2x2_ASAP7_75t_L g377 ( .A(n_266), .B(n_299), .Y(n_377) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g352 ( .A(n_272), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g399 ( .A(n_273), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g430 ( .A(n_274), .Y(n_430) );
INVx2_ASAP7_75t_L g369 ( .A(n_277), .Y(n_369) );
NAND4xp25_ASAP7_75t_L g278 ( .A(n_279), .B(n_288), .C(n_305), .D(n_320), .Y(n_278) );
NAND2xp33_ASAP7_75t_SL g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_281), .A2(n_359), .B1(n_375), .B2(n_377), .C(n_378), .Y(n_374) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g356 ( .A(n_285), .Y(n_356) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
INVx2_ASAP7_75t_L g421 ( .A(n_287), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_293), .B1(n_294), .B2(n_297), .C1(n_300), .C2(n_304), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g375 ( .A(n_291), .B(n_376), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_291), .A2(n_403), .B(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g414 ( .A(n_292), .B(n_358), .Y(n_414) );
OAI21xp33_ASAP7_75t_SL g388 ( .A1(n_293), .A2(n_314), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g307 ( .A(n_296), .B(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_296), .Y(n_359) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g364 ( .A(n_303), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_309), .B1(n_314), .B2(n_319), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_311), .A2(n_321), .B1(n_324), .B2(n_326), .C(n_328), .Y(n_320) );
INVx3_ASAP7_75t_R g435 ( .A(n_312), .Y(n_435) );
INVx1_ASAP7_75t_L g353 ( .A(n_313), .Y(n_353) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_316), .Y(n_370) );
INVx1_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_325), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g398 ( .A(n_325), .Y(n_398) );
AND2x2_ASAP7_75t_L g426 ( .A(n_325), .B(n_373), .Y(n_426) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g420 ( .A(n_330), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_392), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_374), .C(n_388), .Y(n_337) );
NOR3xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_350), .C(n_360), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_341), .A2(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g391 ( .A(n_343), .Y(n_391) );
AND2x2_ASAP7_75t_L g432 ( .A(n_343), .B(n_421), .Y(n_432) );
NAND2x1_ASAP7_75t_L g390 ( .A(n_344), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g404 ( .A(n_358), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_365), .B1(n_367), .B2(n_371), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_366), .B(n_396), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g439 ( .A(n_372), .Y(n_439) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI22xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_381), .B1(n_383), .B2(n_385), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_419), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_399), .C(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_395), .A2(n_409), .B(n_411), .Y(n_408) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_SL g419 ( .A1(n_399), .A2(n_420), .B(n_422), .C(n_424), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_403), .A2(n_408), .B1(n_413), .B2(n_415), .Y(n_407) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B(n_431), .C(n_438), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_431) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI21xp5_ASAP7_75t_SL g668 ( .A1(n_448), .A2(n_657), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_635), .B1(n_652), .B2(n_654), .C(n_658), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B1(n_468), .B2(n_469), .Y(n_453) );
CKINVDCx14_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
XNOR2xp5_ASAP7_75t_SL g455 ( .A(n_456), .B(n_460), .Y(n_455) );
INVx1_ASAP7_75t_SL g459 ( .A(n_458), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g466 ( .A(n_463), .Y(n_466) );
INVx1_ASAP7_75t_L g465 ( .A(n_464), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_562), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_490), .B1(n_491), .B2(n_511), .C(n_512), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_475), .B(n_481), .Y(n_474) );
BUFx3_ASAP7_75t_L g537 ( .A(n_475), .Y(n_537) );
INVx8_ASAP7_75t_L g558 ( .A(n_475), .Y(n_558) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
AND2x4_ASAP7_75t_L g544 ( .A(n_476), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_477), .B(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
AND2x4_ASAP7_75t_L g539 ( .A(n_477), .B(n_527), .Y(n_539) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g545 ( .A(n_480), .Y(n_545) );
AND2x4_ASAP7_75t_L g520 ( .A(n_481), .B(n_502), .Y(n_520) );
AND2x6_ASAP7_75t_L g640 ( .A(n_481), .B(n_517), .Y(n_640) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
NAND3x1_ASAP7_75t_L g553 ( .A(n_482), .B(n_554), .C(n_555), .Y(n_553) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g531 ( .A(n_483), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g647 ( .A(n_483), .B(n_485), .Y(n_647) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND3x4_ASAP7_75t_L g530 ( .A(n_485), .B(n_531), .C(n_532), .Y(n_530) );
INVxp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g623 ( .A(n_487), .B(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g499 ( .A(n_488), .Y(n_499) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_490), .A2(n_577), .B1(n_581), .B2(n_593), .C(n_597), .Y(n_576) );
INVx8_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g527 ( .A(n_497), .Y(n_527) );
INVx1_ASAP7_75t_L g630 ( .A(n_497), .Y(n_630) );
OR2x2_ASAP7_75t_L g627 ( .A(n_498), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g633 ( .A(n_498), .Y(n_633) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g554 ( .A(n_503), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x6_ASAP7_75t_L g597 ( .A(n_505), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_505), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_505), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g567 ( .A(n_506), .B(n_568), .Y(n_567) );
INVx3_ASAP7_75t_L g595 ( .A(n_506), .Y(n_595) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
AND2x2_ASAP7_75t_L g586 ( .A(n_508), .B(n_510), .Y(n_586) );
INVx1_ASAP7_75t_L g626 ( .A(n_508), .Y(n_626) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g575 ( .A(n_510), .Y(n_575) );
AND2x2_ASAP7_75t_L g579 ( .A(n_510), .B(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g616 ( .A(n_510), .Y(n_616) );
NAND3xp33_ASAP7_75t_SL g512 ( .A(n_513), .B(n_528), .C(n_559), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_521), .B2(n_522), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g599 ( .A1(n_514), .A2(n_521), .B1(n_600), .B2(n_602), .C1(n_611), .C2(n_612), .Y(n_599) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2x1_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_517), .B(n_643), .C(n_646), .Y(n_642) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g547 ( .A(n_519), .B(n_526), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_519), .B(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g522 ( .A(n_520), .B(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g560 ( .A(n_520), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI33xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_534), .A3(n_540), .B1(n_548), .B2(n_551), .B3(n_556), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g620 ( .A(n_533), .Y(n_620) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g561 ( .A(n_539), .Y(n_561) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx8_ASAP7_75t_L g549 ( .A(n_544), .Y(n_549) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g550 ( .A(n_547), .Y(n_550) );
AND2x4_ASAP7_75t_L g634 ( .A(n_549), .B(n_633), .Y(n_634) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g632 ( .A(n_557), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_617), .B(n_621), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g563 ( .A(n_564), .B(n_576), .C(n_599), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_570), .B2(n_571), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_565), .A2(n_570), .B1(n_632), .B2(n_634), .Y(n_631) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g572 ( .A(n_568), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g577 ( .A(n_568), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_568), .B(n_598), .Y(n_601) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx3_ASAP7_75t_L g588 ( .A(n_574), .Y(n_588) );
INVx2_ASAP7_75t_L g606 ( .A(n_574), .Y(n_606) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g596 ( .A(n_579), .Y(n_596) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_586), .Y(n_598) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx4_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g610 ( .A(n_591), .Y(n_610) );
AND2x4_ASAP7_75t_L g609 ( .A(n_592), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
BUFx3_ASAP7_75t_L g607 ( .A(n_598), .Y(n_607) );
BUFx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .Y(n_622) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx8_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B(n_642), .C(n_648), .Y(n_638) );
AND2x2_ASAP7_75t_L g663 ( .A(n_639), .B(n_642), .Y(n_663) );
INVx4_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g645 ( .A(n_641), .Y(n_645) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g662 ( .A(n_648), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
BUFx2_ASAP7_75t_L g657 ( .A(n_649), .Y(n_657) );
AND2x2_ASAP7_75t_L g669 ( .A(n_649), .B(n_650), .Y(n_669) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g656 ( .A(n_651), .B(n_657), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_664), .B1(n_666), .B2(n_667), .Y(n_658) );
CKINVDCx14_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
BUFx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x6_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
endmodule