module fake_jpeg_5013_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_22),
.B1(n_11),
.B2(n_13),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_35),
.B(n_38),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_22),
.B1(n_19),
.B2(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_17),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_22),
.B1(n_13),
.B2(n_19),
.Y(n_42)
);

OAI22x1_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_43),
.B1(n_35),
.B2(n_29),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_14),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_23),
.B(n_24),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_36),
.C(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_33),
.B1(n_43),
.B2(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_72),
.B1(n_62),
.B2(n_60),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_16),
.B(n_20),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_55),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_57),
.B1(n_30),
.B2(n_21),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_83),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_82),
.B(n_84),
.C(n_29),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_49),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_23),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_66),
.B(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_89),
.C(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_20),
.C(n_12),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_74),
.B(n_23),
.C(n_26),
.D(n_18),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_94),
.C(n_12),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_60),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_79),
.B(n_18),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_14),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_95),
.B1(n_16),
.B2(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_6),
.B(n_9),
.C(n_3),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_3),
.B(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_8),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_103),
.C(n_10),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_0),
.B(n_1),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_0),
.Y(n_108)
);


endmodule