module fake_jpeg_19420_n_287 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_273;
wire n_182;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_24),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_43),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_89),
.B1(n_91),
.B2(n_16),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_70),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_42),
.B(n_37),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_97),
.B(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_27),
.B1(n_18),
.B2(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_63),
.A2(n_73),
.B1(n_78),
.B2(n_99),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_77),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_27),
.B1(n_18),
.B2(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_18),
.B1(n_39),
.B2(n_34),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_75),
.B1(n_0),
.B2(n_1),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_14),
.B1(n_31),
.B2(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_14),
.B1(n_31),
.B2(n_29),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_22),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_0),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_111)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_0),
.B(n_1),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_16),
.B1(n_20),
.B2(n_32),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_97),
.B1(n_80),
.B2(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_16),
.B1(n_20),
.B2(n_32),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_110),
.B1(n_111),
.B2(n_129),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_91),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_125),
.B(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_115),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_0),
.B(n_1),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_2),
.B(n_3),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_91),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_7),
.C(n_10),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_9),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_9),
.B1(n_11),
.B2(n_4),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_81),
.A2(n_82),
.B1(n_67),
.B2(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_65),
.B1(n_66),
.B2(n_84),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_137),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_158),
.B1(n_132),
.B2(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_65),
.C(n_90),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_141),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_79),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_144),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_76),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_98),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_87),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_87),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_151),
.Y(n_175)
);

AO21x2_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_69),
.B(n_64),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_96),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_88),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_155),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_9),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_122),
.B1(n_115),
.B2(n_130),
.Y(n_166)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_127),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_11),
.Y(n_185)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_167),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_129),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_154),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_138),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_164),
.A2(n_174),
.B(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_154),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_130),
.C(n_118),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_173),
.C(n_134),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_114),
.C(n_133),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_112),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_147),
.B(n_105),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_107),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_135),
.B(n_105),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_124),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_191),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_195),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_192),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_145),
.B(n_135),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_175),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_145),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_134),
.C(n_151),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_202),
.C(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_152),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_140),
.C(n_141),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_158),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_147),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_150),
.C(n_133),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_163),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_164),
.B(n_181),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_224),
.B(n_187),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_171),
.B1(n_177),
.B2(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_223),
.B1(n_189),
.B2(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_192),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_166),
.B1(n_184),
.B2(n_170),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_195),
.B(n_206),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_175),
.C(n_173),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.C(n_202),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_181),
.C(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_241),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_192),
.C(n_194),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_235),
.C(n_238),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_225),
.A2(n_210),
.B1(n_224),
.B2(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_203),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_243),
.B(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_246),
.C(n_221),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_226),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_225),
.B1(n_223),
.B2(n_217),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_256),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_227),
.B1(n_211),
.B2(n_189),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_255),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_230),
.A2(n_215),
.B(n_212),
.Y(n_257)
);

AOI31xp33_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_201),
.A3(n_183),
.B(n_207),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_258),
.B1(n_245),
.B2(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_235),
.CI(n_234),
.CON(n_260),
.SN(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_193),
.B1(n_212),
.B2(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_250),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_211),
.B(n_244),
.C(n_213),
.D(n_246),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_265),
.B(n_266),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_208),
.B(n_199),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_256),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_264),
.B(n_259),
.Y(n_276)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_273),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_250),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_277),
.B(n_268),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_267),
.B(n_260),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_267),
.B(n_272),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_281),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_275),
.B(n_270),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_274),
.Y(n_284)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_282),
.A3(n_182),
.B1(n_251),
.B2(n_198),
.C1(n_147),
.C2(n_126),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_182),
.B(n_119),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_155),
.Y(n_287)
);


endmodule