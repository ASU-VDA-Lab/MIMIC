module fake_aes_9745_n_636 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_636);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_636;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g74 ( .A(n_34), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_9), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_43), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_28), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_21), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_52), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_35), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_72), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_7), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_32), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_17), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_25), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_13), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_45), .Y(n_90) );
OR2x2_ASAP7_75t_L g91 ( .A(n_55), .B(n_42), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_66), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_71), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_56), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_24), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_51), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_58), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_49), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_40), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_20), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_39), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_73), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_17), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_48), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_70), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_26), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_60), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_95), .B(n_99), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_75), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_116), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_95), .B(n_0), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_116), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_116), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_116), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_86), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_74), .Y(n_140) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_88), .A2(n_30), .B(n_67), .Y(n_141) );
NAND2xp33_ASAP7_75t_SL g142 ( .A(n_114), .B(n_1), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_96), .B(n_2), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_102), .B(n_3), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_76), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_79), .Y(n_147) );
INVxp67_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_79), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_106), .B(n_3), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_90), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_77), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_118), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_78), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_132), .B(n_103), .Y(n_158) );
INVx5_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_127), .B(n_91), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_127), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_132), .B(n_103), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
INVx1_ASAP7_75t_SL g167 ( .A(n_152), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
INVx5_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_135), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_123), .B(n_111), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_152), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_127), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_143), .B(n_94), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_125), .B(n_111), .Y(n_182) );
NAND3x1_ASAP7_75t_L g183 ( .A(n_144), .B(n_117), .C(n_112), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_148), .B(n_82), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_124), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_124), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_152), .B(n_80), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_121), .B(n_100), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_129), .Y(n_191) );
OR2x2_ASAP7_75t_SL g192 ( .A(n_139), .B(n_113), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_146), .B(n_82), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_133), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_119), .B(n_100), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_156), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_119), .B(n_84), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_137), .B(n_91), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_142), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_143), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_146), .B(n_84), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_155), .A2(n_115), .B1(n_87), .B2(n_97), .Y(n_203) );
AND3x4_ASAP7_75t_L g204 ( .A(n_149), .B(n_110), .C(n_147), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_124), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_130), .B(n_97), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_130), .B(n_104), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_134), .B(n_107), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_162), .B(n_134), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_195), .B(n_136), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_191), .B(n_157), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_191), .A2(n_136), .B(n_145), .C(n_150), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_195), .B(n_157), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_176), .B(n_155), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
AO22x1_ASAP7_75t_L g221 ( .A1(n_194), .A2(n_87), .B1(n_109), .B2(n_101), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_162), .B(n_120), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_197), .B(n_210), .Y(n_223) );
OR2x6_ASAP7_75t_L g224 ( .A(n_198), .B(n_122), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_206), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_198), .A2(n_120), .B1(n_122), .B2(n_149), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_197), .B(n_120), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g228 ( .A1(n_198), .A2(n_141), .B1(n_98), .B2(n_93), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_162), .B(n_153), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_210), .B(n_120), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_206), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_176), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_193), .B(n_122), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g236 ( .A(n_194), .B(n_153), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_180), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_169), .B(n_153), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_190), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_202), .B(n_122), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g241 ( .A1(n_198), .A2(n_147), .B1(n_138), .B2(n_151), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_182), .B(n_151), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_180), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_188), .B(n_151), .Y(n_244) );
AOI22xp5_ASAP7_75t_SL g245 ( .A1(n_196), .A2(n_141), .B1(n_5), .B2(n_6), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_182), .B(n_147), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_169), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_179), .A2(n_141), .B(n_131), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_158), .B(n_131), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_164), .B(n_131), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_179), .B(n_128), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_200), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_179), .Y(n_257) );
NOR3xp33_ASAP7_75t_SL g258 ( .A(n_203), .B(n_4), .C(n_5), .Y(n_258) );
BUFx12f_ASAP7_75t_L g259 ( .A(n_192), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_201), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_161), .B(n_128), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_189), .A2(n_126), .B(n_128), .C(n_8), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_161), .B(n_135), .Y(n_263) );
NOR2x2_ASAP7_75t_L g264 ( .A(n_192), .B(n_4), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_161), .B(n_135), .Y(n_265) );
INVx5_ASAP7_75t_L g266 ( .A(n_180), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_247), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_225), .A2(n_199), .B1(n_184), .B2(n_187), .C(n_177), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_259), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_215), .B(n_167), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_232), .B(n_187), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_250), .A2(n_183), .B(n_178), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_266), .B(n_208), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_233), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_233), .A2(n_209), .B(n_183), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_223), .B(n_204), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_224), .B(n_207), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_218), .B(n_204), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_216), .A2(n_208), .B(n_126), .C(n_173), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_239), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_242), .B(n_207), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_214), .B(n_207), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_239), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_255), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_220), .Y(n_291) );
AND2x2_ASAP7_75t_SL g292 ( .A(n_220), .B(n_209), .Y(n_292) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_229), .Y(n_293) );
BUFx12f_ASAP7_75t_L g294 ( .A(n_224), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_211), .A2(n_209), .B(n_163), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_256), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_241), .A2(n_163), .B(n_173), .C(n_166), .Y(n_297) );
CKINVDCx6p67_ASAP7_75t_R g298 ( .A(n_224), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_229), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
O2A1O1Ixp5_ASAP7_75t_SL g301 ( .A1(n_263), .A2(n_171), .B(n_181), .C(n_166), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_229), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_221), .Y(n_303) );
BUFx2_ASAP7_75t_SL g304 ( .A(n_266), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_211), .A2(n_175), .B(n_171), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_260), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_241), .A2(n_207), .B1(n_159), .B2(n_170), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_226), .A2(n_207), .B1(n_205), .B2(n_186), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_227), .B(n_207), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_295), .A2(n_228), .B(n_252), .Y(n_311) );
OAI21x1_ASAP7_75t_SL g312 ( .A1(n_279), .A2(n_262), .B(n_261), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_301), .A2(n_265), .B(n_263), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_296), .B(n_226), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_281), .B(n_237), .Y(n_316) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_294), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_301), .A2(n_265), .B(n_251), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_296), .B(n_244), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_276), .A2(n_238), .B(n_230), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_280), .A2(n_248), .B1(n_257), .B2(n_249), .Y(n_322) );
AOI21x1_ASAP7_75t_L g323 ( .A1(n_276), .A2(n_175), .B(n_181), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_278), .Y(n_324) );
NOR2x1_ASAP7_75t_R g325 ( .A(n_294), .B(n_266), .Y(n_325) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_271), .Y(n_326) );
BUFx2_ASAP7_75t_SL g327 ( .A(n_281), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_274), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_297), .A2(n_235), .B(n_240), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_267), .A2(n_222), .B(n_254), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_281), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_306), .B(n_244), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_278), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_267), .A2(n_230), .B(n_238), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_281), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_303), .A2(n_236), .B1(n_231), .B2(n_243), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_308), .A2(n_290), .B(n_305), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_290), .A2(n_288), .B(n_289), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_307), .B(n_266), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_315), .Y(n_340) );
OAI211xp5_ASAP7_75t_L g341 ( .A1(n_326), .A2(n_258), .B(n_268), .C(n_303), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_327), .A2(n_271), .B1(n_282), .B2(n_245), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_328), .B(n_272), .Y(n_343) );
OR2x6_ASAP7_75t_L g344 ( .A(n_327), .B(n_304), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_324), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_314), .A2(n_309), .B1(n_298), .B2(n_288), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_333), .B(n_275), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_333), .B(n_275), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_314), .A2(n_269), .B1(n_258), .B2(n_283), .C(n_287), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_328), .B(n_298), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_320), .B(n_306), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_320), .A2(n_286), .B1(n_264), .B2(n_289), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_310), .B1(n_212), .B2(n_213), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_335), .A2(n_292), .B1(n_217), .B2(n_270), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_319), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_332), .B(n_217), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_332), .A2(n_257), .B1(n_248), .B2(n_249), .C(n_277), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_311), .B(n_159), .C(n_170), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_331), .A2(n_292), .B1(n_300), .B2(n_302), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_319), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_354), .B(n_338), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_356), .A2(n_331), .B1(n_339), .B2(n_317), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_354), .B(n_338), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_365), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_342), .A2(n_339), .B1(n_317), .B2(n_311), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_358), .B(n_330), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_358), .B(n_330), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_345), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_345), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_348), .A2(n_339), .B1(n_317), .B2(n_312), .Y(n_377) );
INVx8_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_346), .B(n_329), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_351), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_346), .B(n_321), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_347), .B(n_321), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_352), .A2(n_312), .B1(n_322), .B2(n_336), .C(n_339), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_349), .B(n_316), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_344), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_360), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_349), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_350), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_344), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_347), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_341), .A2(n_316), .B1(n_323), .B2(n_126), .C(n_300), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_350), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_379), .A2(n_363), .B(n_323), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_373), .B(n_366), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_373), .B(n_355), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_372), .B(n_343), .C(n_359), .Y(n_402) );
NAND2x1_ASAP7_75t_L g403 ( .A(n_373), .B(n_385), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_397), .B(n_353), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_367), .A2(n_377), .B1(n_384), .B2(n_353), .C(n_396), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_378), .B(n_325), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_397), .B(n_325), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_380), .B(n_361), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_366), .B(n_329), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_392), .A2(n_357), .B1(n_362), .B2(n_364), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_374), .B(n_313), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_384), .B(n_396), .C(n_375), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_392), .B(n_7), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_383), .B(n_337), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_391), .B(n_334), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_378), .A2(n_334), .B(n_292), .C(n_337), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_374), .B(n_313), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_378), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_385), .B(n_300), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_370), .B(n_318), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx4_ASAP7_75t_L g427 ( .A(n_378), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g428 ( .A1(n_386), .A2(n_8), .A3(n_10), .B1(n_11), .B2(n_12), .B3(n_13), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_391), .B(n_318), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_368), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_391), .A2(n_300), .B1(n_304), .B2(n_302), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_379), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_382), .B(n_12), .Y(n_433) );
AOI33xp33_ASAP7_75t_L g434 ( .A1(n_382), .A2(n_383), .A3(n_393), .B1(n_390), .B2(n_389), .B3(n_387), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_371), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_371), .B(n_14), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_389), .B(n_14), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_368), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_390), .B(n_15), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_378), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_386), .B(n_368), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_378), .Y(n_442) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_388), .B(n_291), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_440), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_430), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_401), .B(n_381), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_401), .B(n_381), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_434), .B(n_388), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_418), .A2(n_393), .B(n_369), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_412), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_404), .B(n_381), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_400), .B(n_409), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_400), .B(n_383), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_398), .B(n_383), .Y(n_456) );
OR2x6_ASAP7_75t_L g457 ( .A(n_403), .B(n_393), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_398), .B(n_394), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_428), .A2(n_395), .B1(n_394), .B2(n_369), .C1(n_135), .C2(n_16), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_438), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_419), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_426), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_423), .B(n_369), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_423), .B(n_395), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_424), .B(n_394), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_416), .B(n_394), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_427), .B(n_18), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_435), .B(n_135), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_424), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_436), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_438), .Y(n_472) );
NAND3xp33_ASAP7_75t_SL g473 ( .A(n_406), .B(n_178), .C(n_174), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_410), .B(n_135), .Y(n_474) );
OAI31xp33_ASAP7_75t_L g475 ( .A1(n_405), .A2(n_302), .A3(n_284), .B(n_160), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_410), .B(n_174), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_435), .B(n_168), .Y(n_478) );
AOI32xp33_ASAP7_75t_L g479 ( .A1(n_415), .A2(n_160), .A3(n_168), .B1(n_284), .B2(n_205), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_441), .B(n_186), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_413), .B(n_170), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_432), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_408), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_413), .B(n_170), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_440), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_437), .B(n_170), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_420), .B(n_159), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_437), .B(n_159), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_408), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_439), .B(n_159), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_439), .B(n_185), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_417), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_420), .B(n_19), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_422), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_425), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_425), .B(n_185), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_452), .B(n_403), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_448), .A2(n_433), .B(n_414), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_429), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_444), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_453), .B(n_443), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_448), .A2(n_427), .B1(n_442), .B2(n_421), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_461), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_461), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_462), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_457), .Y(n_509) );
AOI21xp33_ASAP7_75t_SL g510 ( .A1(n_459), .A2(n_421), .B(n_442), .Y(n_510) );
NOR2xp33_ASAP7_75t_R g511 ( .A(n_486), .B(n_442), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_453), .B(n_483), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_462), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_450), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_496), .B(n_402), .C(n_422), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_490), .B(n_416), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_454), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_470), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_482), .B(n_416), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_465), .B(n_443), .Y(n_521) );
OAI21xp5_ASAP7_75t_SL g522 ( .A1(n_475), .A2(n_421), .B(n_411), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_446), .Y(n_523) );
NOR2xp67_ASAP7_75t_SL g524 ( .A(n_495), .B(n_427), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_491), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_482), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_485), .B(n_416), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_465), .B(n_443), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_485), .B(n_399), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_456), .B(n_399), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_447), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_469), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_457), .B(n_431), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_471), .B(n_411), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_457), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_477), .B(n_399), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_497), .B(n_431), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_466), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_474), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_464), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_497), .B(n_29), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_494), .B(n_33), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_494), .B(n_37), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_451), .Y(n_544) );
OAI211xp5_ASAP7_75t_SL g545 ( .A1(n_479), .A2(n_299), .B(n_293), .C(n_46), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_464), .B(n_474), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_445), .Y(n_547) );
AOI21xp33_ASAP7_75t_L g548 ( .A1(n_500), .A2(n_498), .B(n_495), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_510), .A2(n_468), .B(n_449), .C(n_473), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_525), .B(n_467), .Y(n_550) );
OAI22x1_ASAP7_75t_L g551 ( .A1(n_535), .A2(n_467), .B1(n_457), .B2(n_458), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_544), .B(n_456), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_504), .Y(n_553) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_505), .A2(n_492), .B1(n_489), .B2(n_487), .C(n_498), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_505), .A2(n_493), .B1(n_480), .B2(n_484), .C(n_481), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_522), .A2(n_467), .B1(n_484), .B2(n_481), .Y(n_556) );
AND2x2_ASAP7_75t_SL g557 ( .A(n_509), .B(n_458), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_515), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_538), .B(n_476), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_518), .Y(n_560) );
OAI221xp5_ASAP7_75t_SL g561 ( .A1(n_533), .A2(n_488), .B1(n_480), .B2(n_476), .C(n_478), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_539), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_519), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_516), .B(n_488), .C(n_478), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_511), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_545), .A2(n_458), .B(n_460), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_534), .A2(n_472), .B1(n_460), .B2(n_455), .C(n_445), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_502), .A2(n_472), .B(n_455), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_523), .B(n_38), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_531), .B(n_44), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_506), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_536), .A2(n_172), .B1(n_284), .B2(n_273), .C(n_291), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_507), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_540), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_547), .Y(n_575) );
O2A1O1Ixp33_ASAP7_75t_SL g576 ( .A1(n_499), .A2(n_50), .B(n_53), .C(n_54), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_508), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_512), .B(n_57), .Y(n_578) );
AOI322xp5_ASAP7_75t_L g579 ( .A1(n_530), .A2(n_59), .A3(n_61), .B1(n_62), .B2(n_63), .C1(n_64), .C2(n_65), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g580 ( .A1(n_542), .A2(n_69), .B(n_172), .C(n_237), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_526), .Y(n_581) );
OAI222xp33_ASAP7_75t_L g582 ( .A1(n_561), .A2(n_524), .B1(n_533), .B2(n_509), .C1(n_503), .C2(n_546), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_565), .B(n_546), .Y(n_583) );
NAND4xp75_ASAP7_75t_L g584 ( .A(n_556), .B(n_517), .C(n_532), .D(n_528), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_558), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_574), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_564), .B(n_513), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_564), .A2(n_517), .B1(n_514), .B2(n_527), .C(n_520), .Y(n_588) );
NAND4xp25_ASAP7_75t_SL g589 ( .A(n_549), .B(n_521), .C(n_501), .D(n_527), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_567), .B(n_520), .Y(n_590) );
XOR2x2_ASAP7_75t_L g591 ( .A(n_550), .B(n_537), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_553), .B(n_529), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_568), .B(n_529), .C(n_533), .Y(n_593) );
NOR2xp33_ASAP7_75t_SL g594 ( .A(n_557), .B(n_541), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_551), .A2(n_543), .B1(n_542), .B2(n_172), .C(n_291), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_574), .Y(n_596) );
OAI21xp33_ASAP7_75t_L g597 ( .A1(n_550), .A2(n_543), .B(n_172), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_557), .B(n_273), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_560), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_563), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_562), .B(n_172), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_571), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_589), .A2(n_555), .B1(n_554), .B2(n_559), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_598), .A2(n_576), .B(n_580), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_602), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_583), .Y(n_606) );
NOR2x1p5_ASAP7_75t_L g607 ( .A(n_584), .B(n_552), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_586), .A2(n_548), .B(n_579), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_590), .A2(n_577), .B(n_573), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_588), .A2(n_570), .B1(n_566), .B2(n_581), .C(n_575), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_593), .A2(n_570), .B1(n_578), .B2(n_569), .C(n_576), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_582), .A2(n_572), .B1(n_273), .B2(n_291), .C(n_243), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_585), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_596), .B(n_273), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_586), .A2(n_237), .B(n_243), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_607), .B(n_591), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_605), .Y(n_617) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_608), .A2(n_595), .B(n_597), .C(n_587), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_606), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_609), .A2(n_582), .B1(n_600), .B2(n_599), .C(n_592), .Y(n_620) );
OAI22x1_ASAP7_75t_L g621 ( .A1(n_603), .A2(n_598), .B1(n_594), .B2(n_601), .Y(n_621) );
XNOR2xp5_ASAP7_75t_SL g622 ( .A(n_613), .B(n_237), .Y(n_622) );
NOR4xp75_ASAP7_75t_SL g623 ( .A(n_621), .B(n_612), .C(n_610), .D(n_611), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_616), .B(n_604), .Y(n_624) );
OR5x1_ASAP7_75t_L g625 ( .A(n_618), .B(n_604), .C(n_615), .D(n_614), .E(n_291), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_617), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_624), .B(n_619), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_624), .B(n_619), .Y(n_628) );
INVxp33_ASAP7_75t_SL g629 ( .A(n_623), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_629), .A2(n_620), .B(n_626), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_628), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_631), .A2(n_627), .B1(n_625), .B2(n_622), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_632), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_633), .A2(n_630), .B(n_253), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_634), .A2(n_243), .B1(n_253), .B2(n_273), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_253), .B(n_628), .Y(n_636) );
endmodule