module fake_netlist_5_509_n_21 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_21);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_21;

wire n_16;
wire n_12;
wire n_18;
wire n_10;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_20;
wire n_14;
wire n_13;

NAND2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_9),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_2),
.B(n_7),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_1),
.A2(n_3),
.B1(n_8),
.B2(n_0),
.Y(n_12)
);

NAND2xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_4),
.Y(n_14)
);

AND2x4_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_15),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_11),
.B(n_16),
.C(n_10),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_SL g20 ( 
.A(n_19),
.B(n_12),
.C(n_15),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_15),
.B(n_4),
.Y(n_21)
);


endmodule