module fake_jpeg_19898_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_68),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_58),
.Y(n_77)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_58),
.B1(n_49),
.B2(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_56),
.Y(n_81)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_42),
.B1(n_60),
.B2(n_50),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_47),
.B1(n_73),
.B2(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_90),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_54),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_2),
.C(n_3),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_48),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_71),
.B1(n_76),
.B2(n_45),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_104),
.B1(n_86),
.B2(n_7),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_85),
.B1(n_73),
.B2(n_46),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_2),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_19),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_105),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_112),
.B1(n_98),
.B2(n_100),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_114),
.B(n_96),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_102),
.C(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.C(n_111),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_109),
.B1(n_95),
.B2(n_108),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_13),
.B(n_14),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_15),
.A3(n_17),
.B1(n_18),
.B2(n_20),
.C1(n_23),
.C2(n_24),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_25),
.B(n_27),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_29),
.B(n_31),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.C(n_38),
.Y(n_124)
);


endmodule