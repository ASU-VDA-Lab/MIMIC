module fake_jpeg_10014_n_143 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_1),
.C(n_2),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_21),
.C(n_19),
.Y(n_48)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_33),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_26),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_30),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_67),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_32),
.B1(n_37),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_59),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_57),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_22),
.B(n_24),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_33),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_1),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_33),
.B(n_16),
.C(n_31),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_64),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_32),
.B1(n_37),
.B2(n_29),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_22),
.C(n_20),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_26),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_58),
.C(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_86),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_27),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_51),
.B1(n_63),
.B2(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_44),
.C(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_91),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_57),
.B1(n_67),
.B2(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_94),
.B1(n_83),
.B2(n_74),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_55),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_28),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_20),
.B1(n_27),
.B2(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_14),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_24),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_103),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_77),
.C(n_81),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_107),
.C(n_105),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_106),
.B1(n_96),
.B2(n_88),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_81),
.B(n_86),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_112),
.B(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_82),
.B1(n_71),
.B2(n_84),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_97),
.C(n_100),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.C(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_115),
.C(n_120),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_117),
.B(n_121),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_91),
.B(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

AOI211xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_94),
.B(n_95),
.C(n_98),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_82),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_106),
.B1(n_109),
.B2(n_117),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_50),
.B1(n_15),
.B2(n_17),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_107),
.C(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_84),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_39),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_60),
.C(n_17),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_111),
.B(n_99),
.C(n_25),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_127),
.C(n_123),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_17),
.B1(n_60),
.B2(n_39),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_50),
.B1(n_15),
.B2(n_34),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_134),
.A3(n_39),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_3),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_2),
.B(n_3),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_136),
.C(n_5),
.Y(n_141)
);

OAI21x1_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_3),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_8),
.A3(n_12),
.B1(n_11),
.B2(n_10),
.C1(n_7),
.C2(n_13),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_141),
.B(n_4),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_6),
.Y(n_143)
);


endmodule