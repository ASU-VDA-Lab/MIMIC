module fake_netlist_5_403_n_81 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_81);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_81;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_0),
.B(n_20),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

OAI21x1_ASAP7_75t_L g30 ( 
.A1(n_9),
.A2(n_4),
.B(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_4),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_14),
.B1(n_1),
.B2(n_7),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_0),
.C(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_19),
.B1(n_12),
.B2(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

OAI221xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.C(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_27),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_24),
.B(n_30),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_40),
.B(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_30),
.B(n_24),
.C(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_42),
.B(n_44),
.Y(n_54)
);

AO21x2_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_47),
.B(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp67_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_50),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_43),
.B(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_25),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_59),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_55),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_60),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_62),
.Y(n_70)
);

NAND4xp25_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_65),
.C(n_67),
.D(n_63),
.Y(n_71)
);

NAND5xp2_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_55),
.C(n_27),
.D(n_56),
.E(n_29),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_72),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_25),
.B1(n_29),
.B2(n_63),
.Y(n_77)
);

AOI221x1_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_25),
.B1(n_29),
.B2(n_46),
.C(n_63),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_54),
.B1(n_57),
.B2(n_77),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_54),
.Y(n_80)
);

NAND4xp75_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_54),
.C(n_57),
.D(n_80),
.Y(n_81)
);


endmodule