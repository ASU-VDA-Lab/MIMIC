module fake_netlist_5_2524_n_100 (n_29, n_16, n_43, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_100);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_100;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_78;
wire n_65;
wire n_74;
wire n_57;
wire n_96;
wire n_66;
wire n_98;
wire n_60;
wire n_58;
wire n_69;
wire n_94;
wire n_80;
wire n_73;
wire n_92;
wire n_84;
wire n_79;
wire n_47;
wire n_53;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_55;
wire n_99;
wire n_49;
wire n_54;
wire n_67;
wire n_76;
wire n_87;
wire n_64;
wire n_77;
wire n_81;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_12),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_2),
.B1(n_28),
.B2(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_5),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_47),
.B(n_49),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_0),
.C(n_1),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

OAI21x1_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_53),
.B(n_61),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_54),
.B1(n_64),
.B2(n_70),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

OAI222xp33_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_51),
.B1(n_58),
.B2(n_65),
.C1(n_56),
.C2(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_88),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_91),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_85),
.B1(n_75),
.B2(n_77),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_73),
.B1(n_66),
.B2(n_62),
.C(n_68),
.Y(n_98)
);

AOI222xp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_60),
.B1(n_69),
.B2(n_67),
.C1(n_82),
.C2(n_41),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_39),
.B1(n_36),
.B2(n_37),
.Y(n_100)
);


endmodule