module fake_jpeg_1510_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_0),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_41),
.B1(n_44),
.B2(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_71),
.B1(n_50),
.B2(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_67),
.B1(n_40),
.B2(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_42),
.B1(n_52),
.B2(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_40),
.B1(n_46),
.B2(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_77),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_43),
.B1(n_64),
.B2(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_60),
.B(n_59),
.C(n_52),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_49),
.B(n_53),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_62),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_82),
.B(n_43),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_18),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_62),
.B(n_63),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_19),
.B(n_34),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_89),
.B1(n_96),
.B2(n_99),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_3),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_59),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_53),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_5),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_108),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_5),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_6),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_7),
.B(n_8),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_21),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.C(n_107),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_15),
.B(n_33),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_7),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_22),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_123),
.B(n_128),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_117),
.B1(n_112),
.B2(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_8),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_117),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_137),
.B(n_120),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_133),
.B1(n_131),
.B2(n_122),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_124),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_131),
.B1(n_123),
.B2(n_121),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_119),
.B(n_129),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_137),
.C(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_142),
.B(n_143),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_140),
.B(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_9),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_10),
.C(n_11),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_13),
.Y(n_151)
);


endmodule