module fake_netlist_6_764_n_196 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_196);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_196;

wire n_52;
wire n_119;
wire n_146;
wire n_46;
wire n_91;
wire n_163;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_85;
wire n_99;
wire n_66;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_29;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_151;
wire n_110;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_31;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

INVxp33_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_R g66 ( 
.A(n_46),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_40),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_52),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_34),
.B1(n_38),
.B2(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_30),
.B1(n_47),
.B2(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_68),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_34),
.C(n_38),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_43),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_52),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_55),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_81),
.B(n_79),
.C(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_R g94 ( 
.A(n_89),
.B(n_58),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_74),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_63),
.B(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_50),
.B(n_42),
.C(n_36),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_87),
.B(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_68),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_68),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_48),
.B1(n_39),
.B2(n_51),
.C(n_36),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.C(n_98),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_78),
.B1(n_87),
.B2(n_88),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

AO31x2_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_92),
.A3(n_42),
.B(n_100),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_82),
.B(n_88),
.Y(n_109)
);

AO31x2_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_86),
.A3(n_81),
.B(n_85),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_56),
.C(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_66),
.B1(n_64),
.B2(n_78),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_R g116 ( 
.A(n_104),
.B(n_90),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_115),
.Y(n_118)
);

AOI211xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_76),
.B(n_84),
.C(n_48),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_107),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_117),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_117),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_112),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_115),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_108),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_82),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_108),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_76),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_108),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_125),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_109),
.B(n_128),
.Y(n_145)
);

OAI221xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_131),
.B1(n_126),
.B2(n_133),
.C(n_39),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_129),
.A3(n_78),
.B1(n_88),
.B2(n_51),
.Y(n_149)
);

NAND2x1_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_140),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_130),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_68),
.B1(n_88),
.B2(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_132),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_149),
.B(n_91),
.C(n_85),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_153),
.A3(n_157),
.B1(n_159),
.B2(n_151),
.C1(n_156),
.C2(n_152),
.Y(n_162)
);

NOR4xp25_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_0),
.C(n_2),
.D(n_3),
.Y(n_163)
);

NAND4xp25_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_75),
.C(n_5),
.D(n_6),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_108),
.Y(n_165)
);

AOI211xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_3),
.B(n_5),
.C(n_7),
.Y(n_166)
);

OAI211xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_75),
.B(n_9),
.C(n_10),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_110),
.Y(n_168)
);

NOR4xp75_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_8),
.C(n_11),
.D(n_12),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_70),
.B1(n_111),
.B2(n_104),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_70),
.B1(n_13),
.B2(n_16),
.C(n_17),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_113),
.C(n_104),
.Y(n_174)
);

AOI221x1_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_8),
.B1(n_17),
.B2(n_18),
.C(n_111),
.Y(n_175)
);

NAND2x1p5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_172),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_174),
.B1(n_161),
.B2(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

OR3x1_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_182),
.C(n_183),
.Y(n_186)
);

OAI221xp5_ASAP7_75t_R g187 ( 
.A1(n_180),
.A2(n_162),
.B1(n_70),
.B2(n_20),
.C(n_22),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_179),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_181),
.B1(n_180),
.B2(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_192),
.B1(n_191),
.B2(n_188),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_194),
.A2(n_188),
.B1(n_187),
.B2(n_185),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_193),
.B(n_70),
.Y(n_196)
);


endmodule