module fake_netlist_1_5384_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_2), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_0), .B(n_5), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_11), .B(n_0), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_1), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_14), .B(n_15), .C(n_13), .Y(n_19) );
INVx6_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
AO21x2_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_17), .B(n_14), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OAI22xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_20), .B1(n_22), .B2(n_21), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_23), .B1(n_21), .B2(n_2), .C(n_3), .Y(n_27) );
AND4x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_3), .C(n_4), .D(n_6), .Y(n_28) );
NAND4xp75_ASAP7_75t_L g29 ( .A(n_28), .B(n_25), .C(n_21), .D(n_3), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_21), .B1(n_6), .B2(n_7), .Y(n_30) );
OAI22x1_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_28), .B1(n_7), .B2(n_8), .Y(n_31) );
AOI22xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_4), .B1(n_8), .B2(n_9), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_31), .Y(n_33) );
AOI22xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_10), .B1(n_32), .B2(n_31), .Y(n_34) );
endmodule