module fake_jpeg_18669_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_19),
.B(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_47),
.B1(n_56),
.B2(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_24),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_28),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_30),
.B1(n_29),
.B2(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_61),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_30),
.B1(n_29),
.B2(n_15),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_70),
.B1(n_74),
.B2(n_36),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_35),
.B1(n_32),
.B2(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_81),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_35),
.B1(n_32),
.B2(n_29),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_15),
.B1(n_19),
.B2(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_33),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_50),
.C(n_41),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_64),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_97),
.B1(n_81),
.B2(n_62),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_45),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_100),
.B(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_41),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_82),
.B(n_70),
.C(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_102),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_36),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_62),
.B1(n_72),
.B2(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_1),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_106),
.B1(n_97),
.B2(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_119),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_86),
.Y(n_145)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_73),
.C(n_60),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_128),
.B1(n_104),
.B2(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_125),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_66),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_89),
.B(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_104),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_73),
.B1(n_83),
.B2(n_59),
.Y(n_128)
);

OAI22x1_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_97),
.B1(n_89),
.B2(n_88),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_111),
.B1(n_115),
.B2(n_121),
.Y(n_157)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_103),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_99),
.C(n_86),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_137),
.C(n_158),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_127),
.B1(n_31),
.B2(n_23),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_118),
.C(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_149),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_157),
.B(n_26),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_101),
.B1(n_108),
.B2(n_83),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_26),
.B1(n_31),
.B2(n_23),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_93),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_150),
.B1(n_108),
.B2(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_92),
.B1(n_94),
.B2(n_100),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_105),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_4),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_107),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_4),
.C(n_5),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_104),
.C(n_108),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_23),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_161),
.A2(n_169),
.B1(n_135),
.B2(n_159),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_181),
.B1(n_156),
.B2(n_139),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_20),
.B(n_5),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_168),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_20),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_170),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_31),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_31),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_26),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_180),
.B1(n_159),
.B2(n_151),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_22),
.B1(n_7),
.B2(n_8),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_136),
.C(n_142),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_196),
.B1(n_176),
.B2(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_150),
.C(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_192),
.C(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_157),
.C(n_149),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_158),
.C(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_146),
.C(n_156),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_162),
.C(n_168),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_180),
.B1(n_190),
.B2(n_192),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_138),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_199),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_138),
.B1(n_22),
.B2(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_167),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_210),
.C(n_22),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_173),
.B(n_176),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_161),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_174),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_212),
.A2(n_213),
.B1(n_197),
.B2(n_184),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_196),
.B(n_195),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_217),
.A2(n_216),
.B(n_219),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_174),
.B(n_165),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_188),
.B(n_194),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_223),
.Y(n_233)
);

FAx1_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_193),
.CI(n_181),
.CON(n_222),
.SN(n_222)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_202),
.B(n_210),
.C(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_202),
.C(n_201),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_217),
.Y(n_240)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

AOI31xp67_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_189),
.A3(n_10),
.B(n_13),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_9),
.C(n_10),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_234),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_14),
.C(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_240),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_229),
.Y(n_241)
);

NAND2xp67_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_234),
.C(n_226),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_226),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_247),
.B(n_245),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_252),
.Y(n_254)
);


endmodule