module real_aes_8799_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g238 ( .A1(n_0), .A2(n_239), .B(n_240), .C(n_244), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_1), .B(n_180), .Y(n_245) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g461 ( .A(n_2), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_3), .B(n_152), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_4), .A2(n_138), .B(n_143), .C(n_506), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_5), .A2(n_133), .B(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_6), .A2(n_133), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_7), .B(n_180), .Y(n_550) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_8), .A2(n_168), .B(n_184), .Y(n_183) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_10), .A2(n_138), .B(n_143), .C(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g488 ( .A(n_11), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_12), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_12), .B(n_42), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_13), .B(n_243), .Y(n_508) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_15), .B(n_152), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_153), .B(n_496), .C(n_498), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_17), .B(n_180), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_18), .A2(n_470), .B1(n_747), .B2(n_753), .C1(n_756), .C2(n_757), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_19), .B(n_217), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_20), .A2(n_143), .B(n_194), .C(n_213), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_21), .A2(n_192), .B(n_242), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_22), .B(n_243), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_23), .B(n_243), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_24), .Y(n_535) );
INVx1_ASAP7_75t_L g527 ( .A(n_25), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_26), .A2(n_143), .B(n_187), .C(n_194), .Y(n_186) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_28), .Y(n_504) );
INVx1_ASAP7_75t_L g584 ( .A(n_29), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_30), .A2(n_133), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_32), .A2(n_141), .B(n_156), .C(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_33), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_34), .A2(n_242), .B(n_547), .C(n_549), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_35), .A2(n_104), .B1(n_115), .B2(n_763), .Y(n_103) );
INVxp67_ASAP7_75t_L g585 ( .A(n_36), .Y(n_585) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_37), .A2(n_47), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_37), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_38), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_39), .A2(n_143), .B(n_194), .C(n_526), .Y(n_525) );
CKINVDCx14_ASAP7_75t_R g545 ( .A(n_40), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_41), .A2(n_46), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_41), .Y(n_752) );
INVx1_ASAP7_75t_L g109 ( .A(n_42), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_43), .A2(n_244), .B(n_486), .C(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_44), .B(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_45), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_46), .Y(n_751) );
INVx1_ASAP7_75t_L g125 ( .A(n_47), .Y(n_125) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_48), .A2(n_122), .A3(n_456), .B1(n_463), .B2(n_464), .C(n_466), .Y(n_121) );
INVx1_ASAP7_75t_L g463 ( .A(n_48), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_49), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_50), .B(n_133), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_51), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_52), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_53), .A2(n_141), .B(n_146), .C(n_156), .Y(n_140) );
INVx1_ASAP7_75t_L g241 ( .A(n_54), .Y(n_241) );
INVx1_ASAP7_75t_L g147 ( .A(n_55), .Y(n_147) );
INVx1_ASAP7_75t_L g516 ( .A(n_56), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_57), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_58), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_59), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g484 ( .A(n_60), .Y(n_484) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_62), .B(n_133), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_63), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_64), .A2(n_174), .B(n_176), .C(n_178), .Y(n_173) );
INVx1_ASAP7_75t_L g161 ( .A(n_65), .Y(n_161) );
INVx1_ASAP7_75t_SL g548 ( .A(n_66), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_68), .B(n_152), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_69), .B(n_180), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_70), .B(n_153), .Y(n_255) );
INVx1_ASAP7_75t_L g538 ( .A(n_71), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_72), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_73), .B(n_149), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_74), .A2(n_143), .B(n_156), .C(n_226), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_75), .Y(n_172) );
INVx1_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_77), .A2(n_133), .B(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_78), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_79), .A2(n_133), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_80), .A2(n_211), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g494 ( .A(n_81), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_82), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_83), .B(n_148), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_84), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_84), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_85), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_86), .A2(n_133), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g497 ( .A(n_87), .Y(n_497) );
INVx2_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
INVx1_ASAP7_75t_L g507 ( .A(n_89), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_90), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_91), .B(n_243), .Y(n_256) );
INVx2_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
OR2x2_ASAP7_75t_L g458 ( .A(n_92), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g746 ( .A(n_92), .B(n_460), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_93), .A2(n_143), .B(n_156), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_94), .B(n_133), .Y(n_200) );
INVx1_ASAP7_75t_L g203 ( .A(n_95), .Y(n_203) );
INVxp67_ASAP7_75t_L g177 ( .A(n_96), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_97), .B(n_168), .Y(n_489) );
INVx2_ASAP7_75t_L g519 ( .A(n_98), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g227 ( .A(n_100), .Y(n_227) );
INVx1_ASAP7_75t_L g251 ( .A(n_101), .Y(n_251) );
AND2x2_ASAP7_75t_L g163 ( .A(n_102), .B(n_158), .Y(n_163) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g764 ( .A(n_107), .Y(n_764) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x2_ASAP7_75t_L g475 ( .A(n_111), .B(n_460), .Y(n_475) );
NOR2x2_ASAP7_75t_L g755 ( .A(n_111), .B(n_459), .Y(n_755) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_468), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g762 ( .A(n_119), .Y(n_762) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_122), .B(n_465), .Y(n_464) );
XOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_126), .A2(n_472), .B1(n_476), .B2(n_743), .Y(n_471) );
INVx4_ASAP7_75t_L g760 ( .A(n_126), .Y(n_760) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR5x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_329), .C(n_407), .D(n_431), .E(n_448), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_195), .B(n_246), .C(n_306), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
AND2x2_ASAP7_75t_L g260 ( .A(n_130), .B(n_166), .Y(n_260) );
INVx5_ASAP7_75t_SL g288 ( .A(n_130), .Y(n_288) );
AND2x2_ASAP7_75t_L g324 ( .A(n_130), .B(n_309), .Y(n_324) );
OR2x2_ASAP7_75t_L g363 ( .A(n_130), .B(n_165), .Y(n_363) );
OR2x2_ASAP7_75t_L g394 ( .A(n_130), .B(n_285), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_130), .B(n_298), .Y(n_430) );
AND2x2_ASAP7_75t_L g442 ( .A(n_130), .B(n_285), .Y(n_442) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_140), .B(n_158), .Y(n_131) );
BUFx2_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_134), .B(n_138), .Y(n_252) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_137), .Y(n_243) );
INVx4_ASAP7_75t_SL g157 ( .A(n_138), .Y(n_157) );
BUFx3_ASAP7_75t_L g194 ( .A(n_138), .Y(n_194) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_157), .B(n_172), .C(n_173), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_142), .A2(n_157), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_142), .A2(n_157), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_142), .A2(n_157), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_142), .A2(n_157), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_142), .A2(n_157), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g580 ( .A1(n_142), .A2(n_157), .B(n_581), .C(n_582), .Y(n_580) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_154), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_148), .A2(n_154), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp5_ASAP7_75t_L g506 ( .A1(n_148), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_148), .A2(n_509), .B(n_538), .C(n_539), .Y(n_537) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_152), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g239 ( .A(n_152), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_152), .A2(n_216), .B(n_527), .C(n_528), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_152), .A2(n_175), .B1(n_584), .B2(n_585), .Y(n_583) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_153), .B(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g244 ( .A(n_155), .Y(n_244) );
INVx1_ASAP7_75t_L g498 ( .A(n_155), .Y(n_498) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_158), .A2(n_482), .B(n_489), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_158), .A2(n_252), .B(n_524), .C(n_525), .Y(n_523) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g169 ( .A(n_159), .B(n_160), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g441 ( .A(n_164), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g304 ( .A(n_165), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_166), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
INVx3_ASAP7_75t_L g312 ( .A(n_166), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_166), .B(n_182), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_166), .B(n_288), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_166), .B(n_309), .Y(n_349) );
AND2x2_ASAP7_75t_L g355 ( .A(n_166), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g392 ( .A(n_166), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_166), .B(n_249), .Y(n_406) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_179), .Y(n_166) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_167), .A2(n_492), .B(n_499), .Y(n_491) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_167), .A2(n_514), .B(n_520), .Y(n_513) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_167), .A2(n_543), .B(n_550), .Y(n_542) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g181 ( .A(n_168), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_168), .A2(n_185), .B(n_186), .Y(n_184) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g259 ( .A(n_169), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_175), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_175), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_178), .B(n_583), .Y(n_582) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_180), .A2(n_235), .B(n_245), .Y(n_234) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_181), .B(n_206), .Y(n_205) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_224), .B(n_232), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_181), .B(n_233), .Y(n_232) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_181), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_181), .B(n_530), .Y(n_529) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_181), .A2(n_534), .B(n_540), .Y(n_533) );
OR2x2_ASAP7_75t_L g298 ( .A(n_182), .B(n_249), .Y(n_298) );
AND2x2_ASAP7_75t_L g309 ( .A(n_182), .B(n_285), .Y(n_309) );
AND2x2_ASAP7_75t_L g321 ( .A(n_182), .B(n_312), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_182), .B(n_249), .Y(n_344) );
INVx1_ASAP7_75t_SL g356 ( .A(n_182), .Y(n_356) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g248 ( .A(n_183), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_183), .B(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B(n_191), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_191), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_207), .Y(n_196) );
AND2x2_ASAP7_75t_L g269 ( .A(n_197), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_197), .B(n_222), .Y(n_273) );
AND2x2_ASAP7_75t_L g276 ( .A(n_197), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g301 ( .A(n_197), .B(n_292), .Y(n_301) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_197), .Y(n_320) );
AND2x2_ASAP7_75t_L g341 ( .A(n_197), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g351 ( .A(n_197), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g397 ( .A(n_197), .B(n_280), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_197), .B(n_303), .Y(n_424) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
AND2x2_ASAP7_75t_L g360 ( .A(n_198), .B(n_292), .Y(n_360) );
AND2x2_ASAP7_75t_L g444 ( .A(n_198), .B(n_312), .Y(n_444) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_205), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_207), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_207), .Y(n_433) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g263 ( .A(n_208), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g272 ( .A(n_208), .B(n_270), .Y(n_272) );
INVx5_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
AND2x2_ASAP7_75t_L g303 ( .A(n_208), .B(n_234), .Y(n_303) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_208), .Y(n_340) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_212), .B(n_217), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_218), .B(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_221), .A2(n_503), .B(n_510), .Y(n_502) );
INVx1_ASAP7_75t_L g381 ( .A(n_222), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_222), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g414 ( .A(n_222), .B(n_280), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_222), .A2(n_337), .B(n_444), .C(n_445), .Y(n_443) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
BUFx2_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
INVx2_ASAP7_75t_L g268 ( .A(n_223), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g549 ( .A(n_230), .Y(n_549) );
INVx2_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_234), .B(n_268), .Y(n_277) );
AND2x2_ASAP7_75t_L g368 ( .A(n_234), .B(n_280), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_242), .B(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g486 ( .A(n_243), .Y(n_486) );
INVx2_ASAP7_75t_L g509 ( .A(n_244), .Y(n_509) );
AOI211x1_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_261), .B(n_274), .C(n_299), .Y(n_246) );
INVx1_ASAP7_75t_L g365 ( .A(n_247), .Y(n_365) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_260), .Y(n_247) );
INVx5_ASAP7_75t_SL g285 ( .A(n_249), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_249), .B(n_355), .Y(n_354) );
AOI311xp33_ASAP7_75t_L g373 ( .A1(n_249), .A2(n_374), .A3(n_376), .B(n_377), .C(n_383), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_249), .A2(n_321), .B(n_409), .C(n_412), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_252), .A2(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_252), .A2(n_535), .B(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g577 ( .A(n_259), .Y(n_577) );
INVxp67_ASAP7_75t_L g328 ( .A(n_260), .Y(n_328) );
NAND4xp25_ASAP7_75t_SL g261 ( .A(n_262), .B(n_265), .C(n_271), .D(n_273), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_262), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g319 ( .A(n_263), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_266), .B(n_272), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_266), .B(n_279), .Y(n_399) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_267), .B(n_280), .Y(n_417) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVxp67_ASAP7_75t_L g327 ( .A(n_269), .Y(n_327) );
AND2x4_ASAP7_75t_L g279 ( .A(n_270), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g353 ( .A(n_270), .B(n_292), .Y(n_353) );
INVx1_ASAP7_75t_L g380 ( .A(n_270), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_270), .B(n_367), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_271), .B(n_341), .Y(n_361) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_272), .B(n_294), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_272), .B(n_341), .Y(n_440) );
INVx1_ASAP7_75t_L g451 ( .A(n_273), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .B(n_281), .C(n_289), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g331 ( .A(n_277), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x2_ASAP7_75t_L g290 ( .A(n_279), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_279), .B(n_341), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_279), .B(n_360), .Y(n_384) );
OR2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_280), .B(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g404 ( .A(n_280), .B(n_360), .Y(n_404) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_282), .A2(n_294), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_415) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g305 ( .A(n_285), .B(n_288), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_285), .B(n_355), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_285), .B(n_312), .Y(n_420) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g405 ( .A(n_287), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g419 ( .A(n_287), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_288), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_309), .Y(n_316) );
AND2x2_ASAP7_75t_L g386 ( .A(n_288), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_288), .B(n_335), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_288), .B(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_295), .Y(n_289) );
INVx2_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
OR2x2_ASAP7_75t_L g346 ( .A(n_294), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g449 ( .A(n_294), .B(n_417), .Y(n_449) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI21xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_304), .Y(n_299) );
INVx1_ASAP7_75t_L g453 ( .A(n_300), .Y(n_453) );
INVx2_ASAP7_75t_SL g367 ( .A(n_301), .Y(n_367) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_304), .A2(n_385), .B(n_449), .C(n_450), .Y(n_448) );
OAI322xp33_ASAP7_75t_SL g317 ( .A1(n_305), .A2(n_318), .A3(n_321), .B1(n_322), .B2(n_323), .C1(n_325), .C2(n_328), .Y(n_317) );
INVx2_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_314), .B2(n_316), .C(n_317), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_SL g383 ( .A1(n_308), .A2(n_384), .B1(n_385), .B2(n_388), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_309), .B(n_312), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_309), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g382 ( .A(n_311), .B(n_344), .Y(n_382) );
INVx1_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_316), .A2(n_426), .B(n_428), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp67_ASAP7_75t_SL g379 ( .A(n_320), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_320), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g436 ( .A(n_321), .Y(n_436) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_330), .B(n_357), .C(n_373), .D(n_389), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_338), .C(n_350), .Y(n_330) );
INVx1_ASAP7_75t_L g422 ( .A(n_331), .Y(n_422) );
AND2x2_ASAP7_75t_L g370 ( .A(n_332), .B(n_353), .Y(n_370) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_337), .B(n_372), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_346), .B2(n_348), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_340), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_341), .A2(n_380), .B(n_403), .C(n_405), .Y(n_402) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g447 ( .A(n_345), .Y(n_447) );
NAND2xp33_ASAP7_75t_SL g437 ( .A(n_346), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g376 ( .A(n_355), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B(n_362), .C(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_369), .B2(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_367), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_372), .B(n_393), .Y(n_455) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI21xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_381), .B(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .B1(n_398), .B2(n_400), .C(n_402), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_415), .C(n_425), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .C(n_443), .Y(n_431) );
INVx1_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_439), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g465 ( .A(n_458), .Y(n_465) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g467 ( .A(n_465), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_466), .B(n_469), .C(n_761), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI22x1_ASAP7_75t_SL g758 ( .A1(n_472), .A2(n_743), .B1(n_759), .B2(n_760), .Y(n_758) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g759 ( .A(n_476), .Y(n_759) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_673), .Y(n_476) );
NAND5xp2_ASAP7_75t_L g477 ( .A(n_478), .B(n_588), .C(n_620), .D(n_637), .E(n_660), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_521), .B1(n_551), .B2(n_555), .C(n_559), .Y(n_478) );
INVx1_ASAP7_75t_L g700 ( .A(n_479), .Y(n_700) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_500), .Y(n_479) );
AND3x2_ASAP7_75t_L g675 ( .A(n_480), .B(n_502), .C(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_481), .B(n_557), .Y(n_556) );
BUFx3_ASAP7_75t_L g566 ( .A(n_481), .Y(n_566) );
AND2x2_ASAP7_75t_L g570 ( .A(n_481), .B(n_512), .Y(n_570) );
INVx2_ASAP7_75t_L g597 ( .A(n_481), .Y(n_597) );
OR2x2_ASAP7_75t_L g608 ( .A(n_481), .B(n_513), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_481), .B(n_501), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_481), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g687 ( .A(n_481), .B(n_513), .Y(n_687) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_490), .Y(n_569) );
AND2x2_ASAP7_75t_L g628 ( .A(n_490), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_490), .B(n_501), .Y(n_647) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_501), .Y(n_558) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_491), .Y(n_565) );
AND2x2_ASAP7_75t_L g614 ( .A(n_491), .B(n_513), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_491), .B(n_500), .C(n_597), .Y(n_639) );
AND2x2_ASAP7_75t_L g704 ( .A(n_491), .B(n_502), .Y(n_704) );
AND2x2_ASAP7_75t_L g738 ( .A(n_491), .B(n_501), .Y(n_738) );
INVxp67_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_501), .B(n_597), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_501), .B(n_628), .Y(n_636) );
AND2x2_ASAP7_75t_L g686 ( .A(n_501), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g714 ( .A(n_501), .Y(n_714) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g621 ( .A(n_502), .B(n_614), .Y(n_621) );
BUFx3_ASAP7_75t_L g653 ( .A(n_502), .Y(n_653) );
INVx2_ASAP7_75t_L g629 ( .A(n_512), .Y(n_629) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_513), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_521), .A2(n_689), .B1(n_691), .B2(n_692), .Y(n_688) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
AND2x2_ASAP7_75t_L g551 ( .A(n_522), .B(n_552), .Y(n_551) );
INVx3_ASAP7_75t_SL g562 ( .A(n_522), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_522), .B(n_592), .Y(n_624) );
OR2x2_ASAP7_75t_L g643 ( .A(n_522), .B(n_532), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_522), .B(n_600), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_522), .B(n_593), .Y(n_651) );
AND2x2_ASAP7_75t_L g663 ( .A(n_522), .B(n_542), .Y(n_663) );
AND2x2_ASAP7_75t_L g679 ( .A(n_522), .B(n_533), .Y(n_679) );
AND2x4_ASAP7_75t_L g682 ( .A(n_522), .B(n_553), .Y(n_682) );
OR2x2_ASAP7_75t_L g699 ( .A(n_522), .B(n_635), .Y(n_699) );
OR2x2_ASAP7_75t_L g730 ( .A(n_522), .B(n_575), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_522), .B(n_658), .Y(n_732) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_529), .Y(n_522) );
AND2x2_ASAP7_75t_L g606 ( .A(n_531), .B(n_573), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_531), .B(n_593), .Y(n_725) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
AND2x2_ASAP7_75t_L g561 ( .A(n_532), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g592 ( .A(n_532), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g600 ( .A(n_532), .B(n_575), .Y(n_600) );
AND2x2_ASAP7_75t_L g618 ( .A(n_532), .B(n_553), .Y(n_618) );
OR2x2_ASAP7_75t_L g635 ( .A(n_532), .B(n_593), .Y(n_635) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g554 ( .A(n_533), .Y(n_554) );
AND2x2_ASAP7_75t_L g658 ( .A(n_533), .B(n_542), .Y(n_658) );
INVx2_ASAP7_75t_L g553 ( .A(n_542), .Y(n_553) );
INVx1_ASAP7_75t_L g670 ( .A(n_542), .Y(n_670) );
AND2x2_ASAP7_75t_L g720 ( .A(n_542), .B(n_562), .Y(n_720) );
AND2x2_ASAP7_75t_L g572 ( .A(n_552), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g604 ( .A(n_552), .B(n_562), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_552), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_L g591 ( .A(n_553), .B(n_562), .Y(n_591) );
OR2x2_ASAP7_75t_L g707 ( .A(n_554), .B(n_681), .Y(n_707) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_557), .B(n_687), .Y(n_693) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
OAI32xp33_ASAP7_75t_L g649 ( .A1(n_558), .A2(n_650), .A3(n_652), .B1(n_654), .B2(n_655), .Y(n_649) );
OR2x2_ASAP7_75t_L g666 ( .A(n_558), .B(n_608), .Y(n_666) );
OAI21xp33_ASAP7_75t_SL g691 ( .A1(n_558), .A2(n_568), .B(n_596), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B1(n_568), .B2(n_571), .Y(n_559) );
INVxp33_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_561), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_562), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g617 ( .A(n_562), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g717 ( .A(n_562), .B(n_658), .Y(n_717) );
OR2x2_ASAP7_75t_L g741 ( .A(n_562), .B(n_635), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g724 ( .A1(n_563), .A2(n_623), .B(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g601 ( .A(n_565), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_565), .B(n_570), .Y(n_619) );
AND2x2_ASAP7_75t_L g641 ( .A(n_566), .B(n_614), .Y(n_641) );
INVx1_ASAP7_75t_L g654 ( .A(n_566), .Y(n_654) );
OR2x2_ASAP7_75t_L g659 ( .A(n_566), .B(n_593), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_569), .B(n_608), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_570), .A2(n_590), .B1(n_595), .B2(n_599), .Y(n_589) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_573), .A2(n_632), .B1(n_639), .B2(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g716 ( .A(n_573), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_575), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g735 ( .A(n_575), .B(n_618), .Y(n_735) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B(n_586), .Y(n_575) );
INVx1_ASAP7_75t_L g594 ( .A(n_576), .Y(n_594) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_579), .A2(n_587), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_601), .B1(n_602), .B2(n_607), .C(n_609), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_591), .B(n_593), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_591), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g610 ( .A(n_592), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_592), .A2(n_698), .B(n_699), .C(n_700), .Y(n_697) );
AND2x2_ASAP7_75t_L g702 ( .A(n_592), .B(n_682), .Y(n_702) );
O2A1O1Ixp33_ASAP7_75t_SL g740 ( .A1(n_592), .A2(n_681), .B(n_741), .C(n_742), .Y(n_740) );
BUFx3_ASAP7_75t_L g632 ( .A(n_593), .Y(n_632) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_596), .B(n_653), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g715 ( .A1(n_596), .A2(n_716), .B(n_718), .C(n_724), .Y(n_715) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVxp67_ASAP7_75t_L g676 ( .A(n_598), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_600), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g620 ( .A1(n_604), .A2(n_621), .B(n_622), .C(n_630), .Y(n_620) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g705 ( .A(n_608), .Y(n_705) );
OR2x2_ASAP7_75t_L g722 ( .A(n_608), .B(n_652), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_616), .B2(n_619), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_611), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
OR2x2_ASAP7_75t_L g709 ( .A(n_613), .B(n_653), .Y(n_709) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g664 ( .A(n_614), .B(n_654), .Y(n_664) );
INVx1_ASAP7_75t_L g672 ( .A(n_615), .Y(n_672) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_618), .B(n_632), .Y(n_680) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_628), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g737 ( .A(n_629), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B(n_636), .Y(n_630) );
INVx1_ASAP7_75t_L g667 ( .A(n_631), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_632), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_632), .B(n_663), .Y(n_662) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_632), .B(n_658), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_632), .B(n_679), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_632), .A2(n_642), .B(n_682), .C(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
AOI221xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_642), .B1(n_644), .B2(n_648), .C(n_649), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_646), .B(n_654), .Y(n_728) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g739 ( .A1(n_648), .A2(n_663), .B(n_665), .C(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_651), .B(n_658), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_652), .B(n_705), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
INVxp33_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_657), .A2(n_669), .B(n_671), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_657), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_658), .B(n_712), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B1(n_665), .B2(n_667), .C(n_668), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_664), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g698 ( .A(n_670), .Y(n_698) );
NAND5xp2_ASAP7_75t_L g673 ( .A(n_674), .B(n_701), .C(n_715), .D(n_726), .E(n_739), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B(n_684), .C(n_697), .Y(n_674) );
INVx2_ASAP7_75t_SL g721 ( .A(n_675), .Y(n_721) );
NAND4xp25_ASAP7_75t_SL g677 ( .A(n_678), .B(n_680), .C(n_681), .D(n_683), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g684 ( .A1(n_683), .A2(n_685), .B(n_688), .C(n_694), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_686), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_686), .A2(n_727), .B1(n_729), .B2(n_731), .C(n_733), .Y(n_726) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_SL g701 ( .A1(n_702), .A2(n_703), .B1(n_706), .B2(n_708), .C(n_710), .Y(n_701) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_709), .A2(n_732), .B1(n_734), .B2(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_718) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_747), .Y(n_756) );
CKINVDCx16_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
endmodule