module fake_ibex_1357_n_4129 (n_151, n_85, n_599, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_4129);

input n_151;
input n_85;
input n_599;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4129;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3674;
wire n_3255;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_3870;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3653;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3904;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3479;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1841;
wire n_1070;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_772;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3225;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_784;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3874;
wire n_1281;
wire n_3094;
wire n_3217;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_4079;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3800;
wire n_3963;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3788;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3529;
wire n_1711;
wire n_3222;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3855;
wire n_3357;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1566;
wire n_1464;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3868;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_1115;
wire n_1395;
wire n_998;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_4047;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_803;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1539;
wire n_1400;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2352;
wire n_2263;
wire n_2716;
wire n_2212;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_3929;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_1815;
wire n_972;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_3314;
wire n_3747;
wire n_1349;
wire n_961;
wire n_1331;
wire n_1223;
wire n_991;
wire n_2127;
wire n_3891;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4116;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_798;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_2180;
wire n_785;
wire n_1952;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3912;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3666;
wire n_3899;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3736;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_3162;
wire n_2732;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_2182;
wire n_1871;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_3044;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3604;
wire n_1838;
wire n_3649;
wire n_833;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_1622;
wire n_897;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_855;
wire n_2367;
wire n_812;
wire n_3576;
wire n_3236;
wire n_3141;
wire n_3491;
wire n_1961;
wire n_3109;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_1547;
wire n_1586;
wire n_1362;
wire n_946;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_790;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_3014;
wire n_1812;
wire n_2703;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3343;
wire n_3163;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3655;
wire n_3543;
wire n_3791;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_2997;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3919;
wire n_3683;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3430;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_3557;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_2302;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_3247;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3933;
wire n_2262;
wire n_3562;
wire n_3516;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1780;
wire n_1678;
wire n_1091;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_478),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_343),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_389),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_635),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_671),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_77),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_94),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_744),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_588),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_179),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_561),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_756),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_137),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_338),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_33),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_62),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_340),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_193),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_643),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_303),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_448),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_71),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_582),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_690),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_431),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_578),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_390),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_451),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_93),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_131),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_605),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_444),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_403),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_739),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_368),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_282),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_142),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_359),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_741),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_382),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_747),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_733),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_751),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_176),
.Y(n_813)
);

BUFx8_ASAP7_75t_SL g814 ( 
.A(n_176),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_81),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_390),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_18),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_464),
.Y(n_818)
);

CKINVDCx16_ASAP7_75t_R g819 ( 
.A(n_172),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_672),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_689),
.Y(n_821)
);

CKINVDCx14_ASAP7_75t_R g822 ( 
.A(n_117),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_598),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_44),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_164),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_728),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_57),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_703),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_546),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_211),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_92),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_357),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_48),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_292),
.Y(n_834)
);

CKINVDCx16_ASAP7_75t_R g835 ( 
.A(n_756),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_675),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_519),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_326),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_754),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_466),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_321),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_187),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_226),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_749),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_203),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_137),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_736),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_95),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_474),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_727),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_708),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_170),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_395),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_372),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_205),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_431),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_286),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_236),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_515),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_215),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_28),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_762),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_43),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_672),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_276),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_482),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_755),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_648),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_432),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_591),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_467),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_469),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_518),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_50),
.Y(n_874)
);

BUFx10_ASAP7_75t_L g875 ( 
.A(n_346),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_194),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_133),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_257),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_267),
.Y(n_879)
);

BUFx2_ASAP7_75t_SL g880 ( 
.A(n_179),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_614),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_174),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_105),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_593),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_645),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_214),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_331),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_608),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_518),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_288),
.Y(n_890)
);

BUFx8_ASAP7_75t_SL g891 ( 
.A(n_196),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_738),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_34),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_71),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_525),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_488),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_337),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_387),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_83),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_473),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_249),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_591),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_642),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_706),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_0),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_274),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_282),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_753),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_628),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_422),
.Y(n_910)
);

INVxp33_ASAP7_75t_SL g911 ( 
.A(n_263),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_375),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_155),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_546),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_395),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_153),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_368),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_184),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_370),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_276),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_269),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_366),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_497),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_735),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_728),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_527),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_730),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_384),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_401),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_407),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_265),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_497),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_263),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_732),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_197),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_286),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_152),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_532),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_609),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_39),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_520),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_583),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_8),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_73),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_191),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_470),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_625),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_79),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_7),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_494),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_330),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_185),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_708),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_48),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_414),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_606),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_343),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_599),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_391),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_29),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_621),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_446),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_174),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_327),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_735),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_768),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_544),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_490),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_143),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_621),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_321),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_540),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_628),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_88),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_614),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_548),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_493),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_404),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_97),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_612),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_145),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_371),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_478),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_316),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_271),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_486),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_766),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_673),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_398),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_161),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_761),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_744),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_366),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_684),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_105),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_477),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_304),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_745),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_683),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_603),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_750),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_729),
.Y(n_1002)
);

BUFx10_ASAP7_75t_L g1003 ( 
.A(n_563),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_438),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_481),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_528),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_104),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_641),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_287),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_723),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_387),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_32),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_461),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_325),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_7),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_141),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_457),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_175),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_656),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_437),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_138),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_605),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_503),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_316),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_590),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_150),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_765),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_224),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_284),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_295),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_362),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_441),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_108),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_592),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_191),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_631),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_17),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_138),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_440),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_70),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_638),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_509),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_602),
.Y(n_1043)
);

BUFx10_ASAP7_75t_L g1044 ( 
.A(n_630),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_75),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_572),
.Y(n_1046)
);

BUFx5_ASAP7_75t_L g1047 ( 
.A(n_159),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_595),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_458),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_455),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_98),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_153),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_257),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_99),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_118),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_742),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_389),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_185),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_202),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_589),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_249),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_454),
.Y(n_1062)
);

BUFx10_ASAP7_75t_L g1063 ( 
.A(n_209),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_459),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_106),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_714),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_311),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_734),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_532),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_726),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_581),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_523),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_329),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_209),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_365),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_353),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_542),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_746),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_603),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_450),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_24),
.Y(n_1081)
);

BUFx8_ASAP7_75t_SL g1082 ( 
.A(n_644),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_438),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_495),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_456),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_3),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_311),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_313),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_566),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_242),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_328),
.Y(n_1091)
);

BUFx5_ASAP7_75t_L g1092 ( 
.A(n_462),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_235),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_718),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_501),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_122),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_318),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_284),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_606),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_303),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_686),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_56),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_73),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_650),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_608),
.Y(n_1105)
);

BUFx10_ASAP7_75t_L g1106 ( 
.A(n_581),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_80),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_189),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_688),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_505),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_302),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_453),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_270),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_71),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_104),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_541),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_273),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_317),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_268),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_204),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_665),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_764),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_740),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_377),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_42),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_200),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_396),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_122),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_332),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_642),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_481),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_295),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_494),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_576),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_261),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_66),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_202),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_139),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_244),
.Y(n_1139)
);

CKINVDCx14_ASAP7_75t_R g1140 ( 
.A(n_340),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_573),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_480),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_684),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_476),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_391),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_475),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_205),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_619),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_459),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_465),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_739),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_743),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_151),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_413),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_471),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_515),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_484),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_442),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_123),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_163),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_103),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_357),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_702),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_235),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_444),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_294),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_678),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_339),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_748),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_737),
.Y(n_1170)
);

BUFx2_ASAP7_75t_SL g1171 ( 
.A(n_4),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_462),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_404),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_217),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_258),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_448),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_635),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_548),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_731),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_45),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_757),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_333),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_69),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_227),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_306),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_242),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_519),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_758),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_468),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_233),
.Y(n_1190)
);

CKINVDCx14_ASAP7_75t_R g1191 ( 
.A(n_236),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_736),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_173),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_172),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_171),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_84),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_298),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_732),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_630),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_47),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_152),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_547),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_429),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_85),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_214),
.Y(n_1205)
);

BUFx10_ASAP7_75t_L g1206 ( 
.A(n_203),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_627),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_491),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_633),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_686),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_190),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_752),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_722),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_741),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_309),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_118),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_759),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_406),
.Y(n_1218)
);

BUFx8_ASAP7_75t_SL g1219 ( 
.A(n_456),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_401),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_121),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_561),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_822),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_877),
.B(n_883),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1136),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_948),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_979),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1122),
.B(n_0),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1122),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_911),
.B(n_0),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_948),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_847),
.B(n_1),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1086),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1012),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1122),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1161),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_1012),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1180),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_775),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_953),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_819),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1140),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_953),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1191),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_959),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_SL g1246 ( 
.A(n_1033),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_775),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_892),
.B(n_1),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_791),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_834),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_835),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_959),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_996),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_996),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_791),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_798),
.Y(n_1256)
);

CKINVDCx16_ASAP7_75t_R g1257 ( 
.A(n_1077),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_798),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1036),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1036),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1090),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1090),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_799),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_776),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1033),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_785),
.Y(n_1266)
);

INVxp33_ASAP7_75t_SL g1267 ( 
.A(n_901),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_799),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_926),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_1118),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_817),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_817),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_815),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_824),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_827),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_833),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1137),
.B(n_1),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_861),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_863),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1160),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_824),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_831),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_831),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1189),
.B(n_980),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_848),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_960),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_894),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_848),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_905),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_874),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_995),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1007),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_874),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1125),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_SL g1295 ( 
.A(n_1040),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1054),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1125),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1102),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1128),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1128),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1171),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1183),
.B(n_2),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1183),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1196),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1196),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1200),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1103),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1049),
.B(n_2),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1107),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1114),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1200),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1204),
.B(n_2),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1040),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1204),
.Y(n_1314)
);

INVxp33_ASAP7_75t_SL g1315 ( 
.A(n_1216),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1159),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1216),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_814),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1159),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_777),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_893),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_893),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1221),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_811),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_SL g1325 ( 
.A(n_779),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1221),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_808),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_808),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_818),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_818),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_899),
.B(n_3),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_855),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_900),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_900),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_913),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_779),
.B(n_3),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_891),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_866),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_913),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1082),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_872),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_909),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_931),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1219),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_931),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1178),
.B(n_4),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_918),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1051),
.B(n_4),
.Y(n_1348)
);

INVxp67_ASAP7_75t_SL g1349 ( 
.A(n_960),
.Y(n_1349)
);

NOR2xp67_ASAP7_75t_L g1350 ( 
.A(n_816),
.B(n_5),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1046),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_940),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1046),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1099),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1099),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1131),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_779),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_929),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1163),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1226),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1256),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1267),
.A2(n_944),
.B1(n_949),
.B2(n_943),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1224),
.B(n_974),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1286),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1353),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1225),
.B(n_1015),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1286),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1238),
.B(n_1163),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1240),
.B(n_1037),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1268),
.B(n_816),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1231),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1353),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1234),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1286),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1315),
.A2(n_1055),
.B1(n_1065),
.B2(n_1045),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1265),
.Y(n_1376)
);

AND2x6_ASAP7_75t_L g1377 ( 
.A(n_1336),
.B(n_960),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1239),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1264),
.A2(n_919),
.B(n_850),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1237),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1247),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1269),
.A2(n_1096),
.B1(n_1115),
.B2(n_1081),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1265),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1299),
.B(n_770),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1243),
.B(n_850),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1321),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1245),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1322),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1252),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1281),
.B(n_1293),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1326),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1323),
.B(n_770),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1253),
.B(n_773),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1254),
.B(n_773),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1229),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1249),
.A2(n_780),
.B1(n_782),
.B2(n_778),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1235),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1255),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1259),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1284),
.B(n_875),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1258),
.B(n_875),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1263),
.B(n_875),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1313),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1260),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1261),
.B(n_881),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1262),
.B(n_778),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1316),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1319),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1282),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1327),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1328),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1266),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1329),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1273),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1330),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1333),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1271),
.B(n_898),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1301),
.B(n_882),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1272),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1334),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1274),
.B(n_780),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1335),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1283),
.B(n_898),
.Y(n_1423)
);

CKINVDCx8_ASAP7_75t_R g1424 ( 
.A(n_1318),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1339),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1285),
.B(n_898),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1343),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1275),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1288),
.B(n_1003),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1345),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1351),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1354),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1355),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1227),
.A2(n_1236),
.B1(n_1233),
.B2(n_1332),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1356),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1359),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1276),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1282),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1349),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1278),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1279),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1287),
.B(n_1047),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1289),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1291),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1297),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1292),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1296),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1300),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1303),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1290),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1298),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1307),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1305),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1309),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1310),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1228),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1352),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1357),
.B(n_919),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1246),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1246),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1290),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1306),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1295),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1295),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1311),
.B(n_1003),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1325),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1348),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1314),
.B(n_782),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1302),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1331),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1223),
.B(n_783),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1312),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1350),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1308),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1346),
.A2(n_950),
.B(n_938),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1248),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1232),
.B(n_783),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1277),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1325),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1230),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1257),
.A2(n_786),
.B1(n_793),
.B2(n_787),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1294),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1270),
.B(n_786),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1294),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1304),
.B(n_787),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1337),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1304),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1317),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1317),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1242),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1244),
.B(n_938),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1340),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1344),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1241),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1241),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1250),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1227),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1250),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_SL g1499 ( 
.A(n_1251),
.B(n_793),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1251),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1280),
.B(n_796),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1280),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1233),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1320),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1236),
.B(n_950),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1324),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1332),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1338),
.B(n_796),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1338),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1341),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1341),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1342),
.B(n_800),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1342),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1347),
.B(n_800),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1347),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1358),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1358),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1226),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1315),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1286),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1226),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1224),
.B(n_801),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1286),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1286),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1286),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1286),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1224),
.B(n_801),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1286),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1264),
.A2(n_988),
.B(n_971),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1256),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1256),
.Y(n_1531)
);

AND2x4_ASAP7_75t_SL g1532 ( 
.A(n_1268),
.B(n_1003),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1224),
.B(n_1044),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1226),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1239),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1353),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1226),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1286),
.Y(n_1538)
);

INVx4_ASAP7_75t_L g1539 ( 
.A(n_1325),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1353),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1353),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1286),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1286),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1226),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1224),
.B(n_1044),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1286),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1226),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_L g1548 ( 
.A(n_1223),
.B(n_1047),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1226),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1286),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1226),
.Y(n_1551)
);

CKINVDCx11_ASAP7_75t_R g1552 ( 
.A(n_1282),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1239),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1286),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1226),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1224),
.B(n_802),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1286),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1226),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1226),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1226),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1226),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1265),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1224),
.B(n_802),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1226),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1286),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1226),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1226),
.Y(n_1567)
);

INVxp33_ASAP7_75t_SL g1568 ( 
.A(n_1239),
.Y(n_1568)
);

BUFx8_ASAP7_75t_L g1569 ( 
.A(n_1325),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1226),
.Y(n_1570)
);

BUFx8_ASAP7_75t_L g1571 ( 
.A(n_1325),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1226),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1226),
.Y(n_1573)
);

AND2x2_ASAP7_75t_SL g1574 ( 
.A(n_1256),
.B(n_960),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1264),
.B(n_1047),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1226),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1239),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1395),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1562),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1469),
.B(n_771),
.Y(n_1580)
);

INVx8_ASAP7_75t_L g1581 ( 
.A(n_1377),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1379),
.Y(n_1582)
);

INVx4_ASAP7_75t_SL g1583 ( 
.A(n_1377),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1472),
.B(n_1047),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1404),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1404),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1387),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1472),
.B(n_960),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1377),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1562),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1467),
.B(n_1047),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1467),
.B(n_1047),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1470),
.A2(n_1092),
.B1(n_1047),
.B2(n_774),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1377),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1377),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1530),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1389),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1365),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1399),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_SL g1600 ( 
.A(n_1457),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1470),
.B(n_1047),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1397),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1395),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1361),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1397),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1385),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1385),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1379),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1395),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1574),
.A2(n_803),
.B1(n_809),
.B2(n_806),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1372),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1476),
.A2(n_1092),
.B1(n_788),
.B2(n_789),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1476),
.A2(n_1092),
.B1(n_790),
.B2(n_792),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1372),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1536),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1532),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1532),
.Y(n_1617)
);

AND2x6_ASAP7_75t_L g1618 ( 
.A(n_1466),
.B(n_971),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1536),
.Y(n_1619)
);

OR2x6_ASAP7_75t_L g1620 ( 
.A(n_1539),
.B(n_880),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1530),
.B(n_1044),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1364),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1364),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1361),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1569),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1540),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1540),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1379),
.A2(n_1092),
.B1(n_794),
.B2(n_797),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1569),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1541),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1474),
.B(n_772),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1444),
.B(n_1092),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1411),
.Y(n_1633)
);

AND2x6_ASAP7_75t_L g1634 ( 
.A(n_1466),
.B(n_988),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1541),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1480),
.B(n_1092),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1363),
.A2(n_784),
.B1(n_954),
.B2(n_806),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1412),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1376),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_1409),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1531),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_L g1642 ( 
.A(n_1480),
.B(n_1092),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1411),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1529),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1459),
.B(n_1080),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1376),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1413),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1531),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1383),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1412),
.B(n_1414),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1539),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1412),
.B(n_1092),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1574),
.Y(n_1653)
);

BUFx4f_ASAP7_75t_L g1654 ( 
.A(n_1486),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1378),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1533),
.B(n_1063),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1529),
.Y(n_1657)
);

AO22x1_ASAP7_75t_L g1658 ( 
.A1(n_1568),
.A2(n_809),
.B1(n_810),
.B2(n_803),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_L g1659 ( 
.A(n_1486),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1383),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1381),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1444),
.B(n_810),
.Y(n_1662)
);

INVxp33_ASAP7_75t_L g1663 ( 
.A(n_1390),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1412),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1414),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1457),
.B(n_804),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1413),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1414),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1449),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1422),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1422),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1425),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1360),
.B(n_807),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1428),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1364),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1453),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1425),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1432),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1432),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1428),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1545),
.B(n_1063),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1462),
.B(n_1080),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1371),
.B(n_812),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1428),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1373),
.B(n_821),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1428),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1400),
.A2(n_823),
.B1(n_825),
.B2(n_820),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1364),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1447),
.B(n_1451),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1409),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1380),
.B(n_826),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1436),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1440),
.Y(n_1693)
);

INVx5_ASAP7_75t_L g1694 ( 
.A(n_1520),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1440),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1535),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_SL g1697 ( 
.A(n_1511),
.Y(n_1697)
);

BUFx4f_ASAP7_75t_L g1698 ( 
.A(n_1479),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1403),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1403),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1392),
.Y(n_1701)
);

INVxp33_ASAP7_75t_L g1702 ( 
.A(n_1398),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1529),
.A2(n_829),
.B1(n_840),
.B2(n_838),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1475),
.A2(n_844),
.B1(n_858),
.B2(n_846),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1520),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1408),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1366),
.A2(n_1382),
.B1(n_1527),
.B2(n_1522),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1440),
.Y(n_1708)
);

BUFx8_ASAP7_75t_SL g1709 ( 
.A(n_1509),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1475),
.A2(n_859),
.B1(n_864),
.B2(n_862),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1447),
.B(n_820),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1518),
.B(n_865),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1520),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1451),
.B(n_823),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1520),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1452),
.B(n_825),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1452),
.B(n_828),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1523),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1523),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1408),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1478),
.A2(n_966),
.B1(n_984),
.B2(n_961),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1556),
.B(n_1063),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1563),
.B(n_1106),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1519),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1552),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1407),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1401),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1523),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1553),
.B(n_1106),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1523),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1526),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1437),
.B(n_828),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1475),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1386),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1386),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1388),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1388),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1519),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1402),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1441),
.B(n_830),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1542),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1478),
.A2(n_832),
.B1(n_836),
.B2(n_830),
.Y(n_1742)
);

INVx5_ASAP7_75t_L g1743 ( 
.A(n_1542),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1542),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1542),
.Y(n_1745)
);

OR2x6_ASAP7_75t_L g1746 ( 
.A(n_1577),
.B(n_1156),
.Y(n_1746)
);

BUFx10_ASAP7_75t_L g1747 ( 
.A(n_1418),
.Y(n_1747)
);

INVx4_ASAP7_75t_L g1748 ( 
.A(n_1543),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1521),
.B(n_1567),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1534),
.B(n_867),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1543),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1391),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1391),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1543),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1568),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1410),
.Y(n_1756)
);

BUFx10_ASAP7_75t_L g1757 ( 
.A(n_1418),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1537),
.B(n_869),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1415),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1416),
.Y(n_1760)
);

OR2x6_ASAP7_75t_L g1761 ( 
.A(n_1419),
.B(n_1156),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1419),
.B(n_1448),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1550),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1544),
.B(n_885),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1547),
.B(n_886),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1508),
.B(n_832),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1460),
.B(n_887),
.Y(n_1767)
);

AO22x2_ASAP7_75t_L g1768 ( 
.A1(n_1505),
.A2(n_896),
.B1(n_908),
.B2(n_890),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1417),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1398),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1443),
.B(n_813),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_SL g1772 ( 
.A(n_1511),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1362),
.A2(n_837),
.B1(n_839),
.B2(n_836),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1550),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1549),
.A2(n_923),
.B1(n_925),
.B2(n_910),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1550),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1375),
.B(n_839),
.C(n_837),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1439),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1420),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1551),
.A2(n_933),
.B1(n_936),
.B2(n_928),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1439),
.Y(n_1781)
);

AND2x6_ASAP7_75t_L g1782 ( 
.A(n_1463),
.B(n_1202),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1427),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1430),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1367),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1576),
.A2(n_956),
.B1(n_958),
.B2(n_952),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1431),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1433),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1448),
.B(n_1202),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1446),
.B(n_813),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1555),
.B(n_963),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1454),
.B(n_841),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1558),
.B(n_967),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1367),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1374),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1435),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1374),
.Y(n_1797)
);

NOR2x1p5_ASAP7_75t_L g1798 ( 
.A(n_1500),
.B(n_841),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1559),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1560),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1561),
.B(n_1573),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1564),
.Y(n_1802)
);

INVx4_ASAP7_75t_L g1803 ( 
.A(n_1370),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1455),
.B(n_842),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1396),
.B(n_843),
.C(n_842),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1566),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1570),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1445),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1524),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1445),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1572),
.B(n_843),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1423),
.B(n_1106),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1368),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_SL g1814 ( 
.A(n_1571),
.B(n_845),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1525),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1552),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1525),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1506),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1442),
.B(n_813),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1370),
.A2(n_968),
.B1(n_981),
.B2(n_976),
.Y(n_1820)
);

BUFx10_ASAP7_75t_L g1821 ( 
.A(n_1491),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1528),
.Y(n_1822)
);

BUFx4f_ASAP7_75t_L g1823 ( 
.A(n_1464),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1456),
.B(n_845),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1368),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1528),
.Y(n_1826)
);

AND3x2_ASAP7_75t_L g1827 ( 
.A(n_1499),
.B(n_1030),
.C(n_989),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1571),
.Y(n_1828)
);

CKINVDCx20_ASAP7_75t_R g1829 ( 
.A(n_1434),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1538),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1426),
.B(n_1205),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1477),
.B(n_983),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1429),
.B(n_1205),
.Y(n_1833)
);

AND3x1_ASAP7_75t_L g1834 ( 
.A(n_1500),
.B(n_993),
.C(n_985),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1393),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1538),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1546),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1458),
.B(n_994),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1394),
.B(n_998),
.Y(n_1839)
);

INVx4_ASAP7_75t_L g1840 ( 
.A(n_1458),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1554),
.Y(n_1841)
);

INVx4_ASAP7_75t_L g1842 ( 
.A(n_1458),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1369),
.B(n_849),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1438),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1369),
.A2(n_1004),
.B1(n_1011),
.B2(n_1005),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1384),
.B(n_849),
.Y(n_1846)
);

INVxp33_ASAP7_75t_L g1847 ( 
.A(n_1485),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1406),
.B(n_1017),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1557),
.Y(n_1849)
);

CKINVDCx6p67_ASAP7_75t_R g1850 ( 
.A(n_1495),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1473),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1557),
.Y(n_1852)
);

OR2x6_ASAP7_75t_L g1853 ( 
.A(n_1495),
.B(n_1020),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1465),
.B(n_1405),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1405),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1438),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1604),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1624),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1663),
.B(n_1501),
.Y(n_1859)
);

OR2x6_ASAP7_75t_L g1860 ( 
.A(n_1762),
.B(n_1495),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1810),
.B(n_1421),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1584),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1596),
.B(n_1450),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1584),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1581),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1835),
.B(n_1468),
.Y(n_1866)
);

O2A1O1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1637),
.A2(n_1481),
.B(n_1483),
.C(n_1471),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1648),
.A2(n_1491),
.B1(n_1548),
.B2(n_1505),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1601),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1704),
.A2(n_1026),
.B1(n_1032),
.B2(n_1021),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1636),
.A2(n_1575),
.B(n_1442),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1663),
.B(n_1575),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1810),
.B(n_1495),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1808),
.B(n_1492),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1648),
.B(n_1493),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1703),
.B(n_1484),
.C(n_1482),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1641),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1656),
.A2(n_1548),
.B1(n_1514),
.B2(n_1512),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1601),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1701),
.B(n_851),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1581),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1702),
.B(n_1565),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1855),
.B(n_851),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1587),
.B(n_852),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1595),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1651),
.B(n_1488),
.Y(n_1886)
);

INVx4_ASAP7_75t_L g1887 ( 
.A(n_1581),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1597),
.B(n_852),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1599),
.B(n_853),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1799),
.B(n_853),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1800),
.B(n_854),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1802),
.B(n_854),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1655),
.B(n_1661),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1806),
.B(n_856),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1807),
.B(n_856),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1847),
.B(n_1494),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1669),
.B(n_1450),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1662),
.B(n_857),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1662),
.B(n_857),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1813),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1825),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1711),
.B(n_860),
.Y(n_1902)
);

INVxp33_ASAP7_75t_L g1903 ( 
.A(n_1724),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1676),
.B(n_1489),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1711),
.B(n_1714),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1714),
.B(n_860),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1716),
.B(n_873),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1716),
.B(n_873),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1717),
.B(n_876),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1606),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1595),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1847),
.B(n_1494),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_L g1913 ( 
.A(n_1721),
.B(n_1487),
.C(n_1461),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1717),
.B(n_876),
.Y(n_1914)
);

OAI22xp33_ASAP7_75t_SL g1915 ( 
.A1(n_1814),
.A2(n_1461),
.B1(n_1487),
.B2(n_879),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1727),
.B(n_1496),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1739),
.B(n_1498),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1769),
.B(n_1502),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1696),
.B(n_1507),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1582),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1704),
.A2(n_1710),
.B1(n_1703),
.B2(n_1612),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1770),
.B(n_1490),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1821),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1732),
.B(n_878),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1854),
.B(n_1490),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1616),
.B(n_1510),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1732),
.B(n_878),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1854),
.B(n_1507),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1651),
.B(n_1517),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1740),
.B(n_879),
.Y(n_1930)
);

INVx8_ASAP7_75t_L g1931 ( 
.A(n_1620),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1617),
.B(n_1637),
.Y(n_1932)
);

OAI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1755),
.A2(n_1513),
.B1(n_1516),
.B2(n_1510),
.Y(n_1933)
);

INVxp67_ASAP7_75t_L g1934 ( 
.A(n_1818),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1803),
.B(n_1513),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1654),
.B(n_1510),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1762),
.B(n_1516),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1796),
.B(n_1116),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1607),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1591),
.A2(n_1042),
.B(n_1041),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1726),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1738),
.B(n_1724),
.Y(n_1942)
);

NOR3xp33_ASAP7_75t_L g1943 ( 
.A(n_1721),
.B(n_1517),
.C(n_1503),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1654),
.B(n_1510),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1796),
.B(n_1749),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1749),
.B(n_1210),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1821),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1801),
.B(n_1211),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1762),
.B(n_1497),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1682),
.B(n_1497),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1756),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1803),
.B(n_1515),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1688),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1759),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1760),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1779),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1707),
.B(n_1504),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1812),
.B(n_1504),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1853),
.Y(n_1959)
);

NOR3xp33_ASAP7_75t_L g1960 ( 
.A(n_1658),
.B(n_1218),
.C(n_1214),
.Y(n_1960)
);

INVx8_ASAP7_75t_L g1961 ( 
.A(n_1620),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1778),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1625),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1659),
.B(n_1116),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1783),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1801),
.B(n_1211),
.Y(n_1966)
);

NOR2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1629),
.B(n_1504),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1781),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1785),
.Y(n_1969)
);

O2A1O1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1811),
.A2(n_1059),
.B(n_1060),
.C(n_1050),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1794),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1831),
.B(n_1504),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1784),
.B(n_1222),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1659),
.B(n_1117),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1828),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1740),
.B(n_1117),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1681),
.A2(n_1124),
.B1(n_1127),
.B2(n_1123),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1682),
.B(n_1123),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1850),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1787),
.B(n_1222),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1792),
.B(n_1124),
.Y(n_1981)
);

INVxp67_ASAP7_75t_SL g1982 ( 
.A(n_1589),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1853),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1582),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1682),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1795),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1792),
.B(n_1127),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1710),
.A2(n_1074),
.B1(n_1079),
.B2(n_1069),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1788),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1840),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1804),
.B(n_1129),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1804),
.B(n_1129),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1840),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1797),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1846),
.B(n_1132),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1589),
.B(n_1132),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_SL g1997 ( 
.A1(n_1600),
.A2(n_1073),
.B1(n_1075),
.B2(n_1035),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1620),
.B(n_1085),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1594),
.B(n_1133),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1842),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1846),
.B(n_1133),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1809),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1842),
.Y(n_2003)
);

O2A1O1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1811),
.A2(n_1095),
.B(n_1098),
.C(n_1089),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1833),
.B(n_1424),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_L g2006 ( 
.A(n_1618),
.B(n_1135),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1709),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1594),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1747),
.B(n_1135),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1815),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1582),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1580),
.B(n_1138),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1766),
.B(n_1138),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1722),
.A2(n_1142),
.B1(n_1143),
.B2(n_1141),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1621),
.B(n_1141),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1580),
.A2(n_1121),
.B(n_1130),
.C(n_1105),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1832),
.B(n_1142),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1653),
.A2(n_1139),
.B1(n_1147),
.B2(n_1134),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1832),
.B(n_1143),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1582),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1612),
.A2(n_1158),
.B1(n_1162),
.B2(n_1150),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1843),
.B(n_1144),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1723),
.A2(n_1145),
.B1(n_1146),
.B2(n_1144),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1843),
.B(n_1839),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1746),
.B(n_1145),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1729),
.B(n_1146),
.Y(n_2026)
);

OAI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1610),
.A2(n_1111),
.B1(n_1119),
.B2(n_1088),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1856),
.B(n_1199),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1817),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1747),
.B(n_1148),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1757),
.B(n_1148),
.Y(n_2031)
);

BUFx5_ASAP7_75t_L g2032 ( 
.A(n_1622),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1746),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1689),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1688),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1757),
.B(n_1149),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1839),
.B(n_1149),
.Y(n_2037)
);

AOI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_1653),
.A2(n_1169),
.B1(n_1188),
.B2(n_1165),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1666),
.B(n_1151),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1822),
.Y(n_2040)
);

INVxp67_ASAP7_75t_SL g2041 ( 
.A(n_1608),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1666),
.B(n_1151),
.Y(n_2042)
);

NOR2xp67_ASAP7_75t_L g2043 ( 
.A(n_1777),
.B(n_5),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1583),
.B(n_1152),
.Y(n_2044)
);

AO22x1_ASAP7_75t_L g2045 ( 
.A1(n_1816),
.A2(n_1153),
.B1(n_1154),
.B2(n_1152),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1689),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1826),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1848),
.B(n_1153),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1830),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1583),
.B(n_1154),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1836),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1585),
.Y(n_2052)
);

INVxp67_ASAP7_75t_L g2053 ( 
.A(n_1746),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1586),
.Y(n_2054)
);

OAI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1853),
.A2(n_1164),
.B1(n_1174),
.B2(n_1120),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1848),
.B(n_1155),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1583),
.B(n_1155),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1687),
.B(n_1805),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1631),
.B(n_1157),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_L g2060 ( 
.A(n_1628),
.B(n_1166),
.C(n_1157),
.Y(n_2060)
);

INVx4_ASAP7_75t_L g2061 ( 
.A(n_1618),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1632),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1768),
.A2(n_1167),
.B1(n_1168),
.B2(n_1166),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1631),
.B(n_1167),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_SL g2065 ( 
.A(n_1761),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1773),
.B(n_1199),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1767),
.B(n_1168),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1632),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1709),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1838),
.Y(n_2070)
);

NOR3xp33_ASAP7_75t_SL g2071 ( 
.A(n_1844),
.B(n_1172),
.C(n_1170),
.Y(n_2071)
);

AOI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_1768),
.A2(n_1195),
.B1(n_1194),
.B2(n_1209),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1761),
.B(n_1170),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_1761),
.B(n_1172),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1837),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1742),
.B(n_1175),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1591),
.A2(n_1212),
.B(n_889),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1673),
.B(n_1175),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1789),
.B(n_1215),
.Y(n_2079)
);

OAI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1789),
.A2(n_1220),
.B1(n_1217),
.B2(n_1177),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1789),
.B(n_1176),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1673),
.B(n_1176),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1683),
.B(n_1177),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1838),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1767),
.B(n_1798),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_1824),
.B(n_1179),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1694),
.B(n_1179),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1683),
.B(n_1181),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1685),
.B(n_1181),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1694),
.B(n_1182),
.Y(n_2090)
);

INVx8_ASAP7_75t_L g2091 ( 
.A(n_1618),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1768),
.B(n_1182),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1613),
.A2(n_1593),
.B1(n_1845),
.B2(n_1820),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1685),
.B(n_1184),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1694),
.B(n_1184),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1640),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1733),
.B(n_1193),
.Y(n_2097)
);

A2O1A1Ixp33_ASAP7_75t_L g2098 ( 
.A1(n_1691),
.A2(n_1186),
.B(n_1187),
.C(n_1185),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1820),
.B(n_1185),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1841),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1823),
.Y(n_2101)
);

INVxp67_ASAP7_75t_SL g2102 ( 
.A(n_1608),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1733),
.B(n_1197),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1849),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1733),
.B(n_1197),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1733),
.B(n_1198),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1613),
.A2(n_1198),
.B1(n_1187),
.B2(n_1190),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1734),
.B(n_1735),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1736),
.B(n_1203),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1737),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1824),
.B(n_1698),
.Y(n_2111)
);

AND2x2_ASAP7_75t_SL g2112 ( 
.A(n_1834),
.B(n_895),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1752),
.B(n_1203),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_1600),
.A2(n_1190),
.B1(n_1192),
.B2(n_1186),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1852),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1827),
.B(n_1192),
.Y(n_2116)
);

O2A1O1Ixp33_ASAP7_75t_L g2117 ( 
.A1(n_1642),
.A2(n_795),
.B(n_805),
.C(n_781),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1753),
.Y(n_2118)
);

OAI221xp5_ASAP7_75t_L g2119 ( 
.A1(n_1845),
.A2(n_1208),
.B1(n_1213),
.B2(n_1201),
.C(n_1193),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_1823),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1602),
.B(n_1201),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_1775),
.B(n_1780),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1694),
.B(n_1731),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1605),
.B(n_1208),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1852),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1645),
.A2(n_1782),
.B1(n_1634),
.B2(n_1712),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1633),
.Y(n_2127)
);

AND2x6_ASAP7_75t_SL g2128 ( 
.A(n_1640),
.B(n_1205),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1608),
.B(n_1213),
.Y(n_2129)
);

O2A1O1Ixp33_ASAP7_75t_L g2130 ( 
.A1(n_1642),
.A2(n_870),
.B(n_871),
.C(n_868),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1608),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1827),
.B(n_1786),
.Y(n_2132)
);

NAND2xp33_ASAP7_75t_L g2133 ( 
.A(n_1634),
.B(n_888),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1644),
.B(n_897),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1644),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1731),
.B(n_902),
.Y(n_2136)
);

AND2x6_ASAP7_75t_L g2137 ( 
.A(n_1644),
.B(n_895),
.Y(n_2137)
);

AO21x2_ASAP7_75t_L g2138 ( 
.A1(n_1592),
.A2(n_1067),
.B(n_895),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_1775),
.B(n_884),
.Y(n_2139)
);

NAND2xp33_ASAP7_75t_L g2140 ( 
.A(n_1634),
.B(n_903),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1644),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_1698),
.B(n_904),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1780),
.B(n_1206),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1728),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_1691),
.A2(n_1207),
.B1(n_1206),
.B2(n_1067),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1657),
.B(n_906),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_1786),
.B(n_1206),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1690),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1657),
.B(n_907),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1643),
.Y(n_2150)
);

NOR3xp33_ASAP7_75t_L g2151 ( 
.A(n_1712),
.B(n_1108),
.C(n_1094),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1647),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1731),
.B(n_912),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1667),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1657),
.B(n_914),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1670),
.B(n_915),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1671),
.B(n_916),
.Y(n_2157)
);

INVxp67_ASAP7_75t_L g2158 ( 
.A(n_1697),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1731),
.B(n_917),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1672),
.B(n_920),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1677),
.B(n_921),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1744),
.Y(n_2162)
);

BUFx2_ASAP7_75t_L g2163 ( 
.A(n_1634),
.Y(n_2163)
);

OAI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_1628),
.A2(n_1126),
.B(n_951),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1678),
.Y(n_2165)
);

NOR3xp33_ASAP7_75t_L g2166 ( 
.A(n_1750),
.B(n_1173),
.C(n_924),
.Y(n_2166)
);

A2O1A1Ixp33_ASAP7_75t_L g2167 ( 
.A1(n_1750),
.A2(n_922),
.B(n_930),
.C(n_927),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_1645),
.A2(n_932),
.B1(n_935),
.B2(n_934),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1758),
.B(n_1207),
.Y(n_2169)
);

INVxp67_ASAP7_75t_L g2170 ( 
.A(n_1697),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1758),
.B(n_1207),
.Y(n_2171)
);

BUFx5_ASAP7_75t_L g2172 ( 
.A(n_1622),
.Y(n_2172)
);

AOI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_1645),
.A2(n_937),
.B1(n_941),
.B2(n_939),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_1772),
.Y(n_2174)
);

NOR2xp67_ASAP7_75t_SL g2175 ( 
.A(n_1743),
.B(n_942),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1744),
.Y(n_2176)
);

INVx2_ASAP7_75t_SL g2177 ( 
.A(n_1634),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1764),
.B(n_945),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1851),
.B(n_946),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1744),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1744),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1764),
.B(n_1765),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1743),
.B(n_1593),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_1791),
.B(n_947),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1623),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1679),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1692),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1793),
.B(n_1619),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1905),
.A2(n_1588),
.B(n_1652),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_2182),
.A2(n_1652),
.B(n_1650),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1877),
.B(n_1934),
.Y(n_2191)
);

BUFx4f_ASAP7_75t_L g2192 ( 
.A(n_1931),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1920),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_1945),
.A2(n_1650),
.B(n_1819),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2034),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_1893),
.A2(n_1772),
.B1(n_1829),
.B2(n_1782),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1866),
.B(n_1645),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1857),
.B(n_1858),
.Y(n_2198)
);

OAI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_1862),
.A2(n_1700),
.B(n_1699),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2055),
.A2(n_1829),
.B1(n_1782),
.B2(n_1645),
.Y(n_2200)
);

INVx1_ASAP7_75t_SL g2201 ( 
.A(n_1942),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1866),
.B(n_1782),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2046),
.B(n_1782),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_SL g2204 ( 
.A(n_2007),
.B(n_1690),
.Y(n_2204)
);

INVx11_ASAP7_75t_L g2205 ( 
.A(n_2137),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_1920),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2099),
.B(n_1706),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1920),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1941),
.Y(n_2209)
);

AOI21xp5_ASAP7_75t_L g2210 ( 
.A1(n_1945),
.A2(n_1819),
.B(n_1720),
.Y(n_2210)
);

A2O1A1Ixp33_ASAP7_75t_L g2211 ( 
.A1(n_2188),
.A2(n_1611),
.B(n_1614),
.C(n_1598),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2122),
.B(n_1615),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_2112),
.B(n_1743),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1984),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1983),
.B(n_1728),
.Y(n_2215)
);

AOI21xp5_ASAP7_75t_L g2216 ( 
.A1(n_1921),
.A2(n_1790),
.B(n_1771),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_1931),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_1921),
.A2(n_1871),
.B(n_2108),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1984),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2080),
.A2(n_1627),
.B1(n_1630),
.B2(n_1626),
.Y(n_2220)
);

OAI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1864),
.A2(n_1879),
.B(n_1869),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2058),
.B(n_1635),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1903),
.B(n_1725),
.Y(n_2223)
);

OAI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2062),
.A2(n_1646),
.B(n_1639),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1951),
.B(n_1579),
.Y(n_2225)
);

NAND3xp33_ASAP7_75t_SL g2226 ( 
.A(n_1913),
.B(n_1725),
.C(n_957),
.Y(n_2226)
);

AO21x1_ASAP7_75t_L g2227 ( 
.A1(n_1957),
.A2(n_1609),
.B(n_1649),
.Y(n_2227)
);

OAI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2068),
.A2(n_1660),
.B(n_1665),
.Y(n_2228)
);

HB1xp67_ASAP7_75t_L g2229 ( 
.A(n_1863),
.Y(n_2229)
);

NAND2xp33_ASAP7_75t_L g2230 ( 
.A(n_2091),
.B(n_1763),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_1985),
.B(n_1748),
.Y(n_2231)
);

AO21x1_ASAP7_75t_L g2232 ( 
.A1(n_2134),
.A2(n_2149),
.B(n_2146),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1954),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2126),
.A2(n_1675),
.B1(n_1705),
.B2(n_1748),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1897),
.A2(n_1590),
.B1(n_955),
.B2(n_964),
.Y(n_2235)
);

AOI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_2156),
.A2(n_1684),
.B(n_1680),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_SL g2237 ( 
.A(n_2069),
.B(n_1751),
.Y(n_2237)
);

AOI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_2156),
.A2(n_1695),
.B(n_1686),
.Y(n_2238)
);

OAI21xp33_ASAP7_75t_L g2239 ( 
.A1(n_2013),
.A2(n_965),
.B(n_962),
.Y(n_2239)
);

A2O1A1Ixp33_ASAP7_75t_L g2240 ( 
.A1(n_1970),
.A2(n_1664),
.B(n_1668),
.C(n_1638),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_2061),
.B(n_1776),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1955),
.B(n_1776),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_2061),
.B(n_1959),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2033),
.B(n_1763),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1956),
.Y(n_2245)
);

INVx3_ASAP7_75t_L g2246 ( 
.A(n_1887),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_1887),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1965),
.B(n_969),
.Y(n_2248)
);

A2O1A1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2004),
.A2(n_1664),
.B(n_1668),
.C(n_1638),
.Y(n_2249)
);

AOI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2041),
.A2(n_1715),
.B(n_1713),
.Y(n_2250)
);

INVx4_ASAP7_75t_L g2251 ( 
.A(n_1931),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2092),
.B(n_970),
.Y(n_2252)
);

AOI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2102),
.A2(n_1719),
.B(n_1718),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2053),
.B(n_1730),
.Y(n_2254)
);

NAND2x1p5_ASAP7_75t_L g2255 ( 
.A(n_1865),
.B(n_1674),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1989),
.Y(n_2256)
);

BUFx4f_ASAP7_75t_L g2257 ( 
.A(n_1961),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2070),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1859),
.B(n_972),
.Y(n_2259)
);

AOI21x1_ASAP7_75t_L g2260 ( 
.A1(n_2183),
.A2(n_1745),
.B(n_1741),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1865),
.Y(n_2261)
);

OR2x6_ASAP7_75t_L g2262 ( 
.A(n_1961),
.B(n_1754),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_1865),
.Y(n_2263)
);

INVxp67_ASAP7_75t_L g2264 ( 
.A(n_2065),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2143),
.B(n_973),
.Y(n_2265)
);

AOI21xp33_ASAP7_75t_L g2266 ( 
.A1(n_1867),
.A2(n_1774),
.B(n_1693),
.Y(n_2266)
);

A2O1A1Ixp33_ASAP7_75t_L g2267 ( 
.A1(n_2117),
.A2(n_1693),
.B(n_1708),
.C(n_1674),
.Y(n_2267)
);

OAI21xp5_ASAP7_75t_L g2268 ( 
.A1(n_2155),
.A2(n_1708),
.B(n_1603),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2147),
.B(n_975),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_2168),
.B(n_1093),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2109),
.B(n_977),
.Y(n_2271)
);

INVxp67_ASAP7_75t_L g2272 ( 
.A(n_2065),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2157),
.A2(n_1603),
.B(n_1578),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2109),
.B(n_978),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_1984),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2093),
.A2(n_982),
.B1(n_987),
.B2(n_986),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_2085),
.B(n_990),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2113),
.B(n_991),
.Y(n_2278)
);

BUFx12f_ASAP7_75t_L g2279 ( 
.A(n_2128),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1962),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_1961),
.Y(n_2281)
);

BUFx2_ASAP7_75t_L g2282 ( 
.A(n_1860),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2113),
.B(n_992),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_2079),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2157),
.A2(n_1578),
.B(n_1067),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2085),
.B(n_997),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2084),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2121),
.B(n_999),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2160),
.A2(n_1067),
.B(n_895),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2173),
.B(n_1076),
.Y(n_2290)
);

OAI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_2129),
.A2(n_1001),
.B(n_1000),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2027),
.A2(n_1002),
.B1(n_1008),
.B2(n_1006),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2121),
.B(n_1009),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1968),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2160),
.A2(n_1067),
.B(n_895),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_R g2296 ( 
.A(n_2096),
.B(n_1010),
.Y(n_2296)
);

AOI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2161),
.A2(n_1109),
.B(n_1084),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1978),
.B(n_2025),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2124),
.B(n_1013),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2124),
.B(n_1014),
.Y(n_2300)
);

OAI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_2129),
.A2(n_1018),
.B(n_1016),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1884),
.B(n_1019),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1884),
.B(n_1022),
.Y(n_2303)
);

AOI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2161),
.A2(n_1932),
.B(n_1940),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_1888),
.B(n_1023),
.Y(n_2305)
);

BUFx4f_ASAP7_75t_L g2306 ( 
.A(n_2091),
.Y(n_2306)
);

NOR2x1_ASAP7_75t_L g2307 ( 
.A(n_1963),
.B(n_1084),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1888),
.B(n_1024),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_1949),
.B(n_1025),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1889),
.B(n_1027),
.Y(n_2310)
);

NOR2x1_ASAP7_75t_L g2311 ( 
.A(n_1975),
.B(n_1084),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_SL g2312 ( 
.A(n_2148),
.B(n_1028),
.Y(n_2312)
);

OAI21xp5_ASAP7_75t_L g2313 ( 
.A1(n_2097),
.A2(n_1031),
.B(n_1029),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2077),
.A2(n_1109),
.B(n_1084),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_SL g2315 ( 
.A(n_2091),
.B(n_1034),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2130),
.A2(n_2111),
.B(n_2086),
.C(n_2043),
.Y(n_2316)
);

BUFx4f_ASAP7_75t_L g2317 ( 
.A(n_1860),
.Y(n_2317)
);

BUFx2_ASAP7_75t_L g2318 ( 
.A(n_1860),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_L g2319 ( 
.A(n_2066),
.B(n_1950),
.Y(n_2319)
);

A2O1A1Ixp33_ASAP7_75t_L g2320 ( 
.A1(n_2164),
.A2(n_1109),
.B(n_1084),
.C(n_1039),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1969),
.Y(n_2321)
);

A2O1A1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2164),
.A2(n_1876),
.B(n_1878),
.C(n_2016),
.Y(n_2322)
);

NOR3xp33_ASAP7_75t_L g2323 ( 
.A(n_1915),
.B(n_1043),
.C(n_1038),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_1938),
.A2(n_1109),
.B(n_1052),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_1938),
.A2(n_1109),
.B(n_1053),
.Y(n_2325)
);

INVx4_ASAP7_75t_L g2326 ( 
.A(n_1979),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_1883),
.A2(n_1056),
.B(n_1048),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1971),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_1883),
.A2(n_1058),
.B(n_1057),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_1881),
.Y(n_2330)
);

OR2x6_ASAP7_75t_L g2331 ( 
.A(n_2158),
.B(n_5),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_1880),
.B(n_1083),
.Y(n_2332)
);

AOI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_2103),
.A2(n_1062),
.B(n_1061),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1986),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2005),
.B(n_1064),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_1889),
.A2(n_1973),
.B1(n_1980),
.B2(n_1868),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_1973),
.A2(n_1068),
.B1(n_1070),
.B2(n_1066),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_2011),
.Y(n_2338)
);

A2O1A1Ixp33_ASAP7_75t_L g2339 ( 
.A1(n_1928),
.A2(n_1072),
.B(n_1078),
.C(n_1071),
.Y(n_2339)
);

O2A1O1Ixp33_ASAP7_75t_L g2340 ( 
.A1(n_2098),
.A2(n_1091),
.B(n_1097),
.C(n_1087),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2103),
.A2(n_1101),
.B(n_1100),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2105),
.A2(n_1110),
.B(n_1104),
.Y(n_2342)
);

NAND2x1_ASAP7_75t_L g2343 ( 
.A(n_2137),
.B(n_6),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_1980),
.A2(n_1890),
.B1(n_1892),
.B2(n_1891),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_1943),
.A2(n_1113),
.B1(n_1112),
.B2(n_8),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1994),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1890),
.B(n_6),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2169),
.B(n_6),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2002),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2010),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1891),
.B(n_7),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_2101),
.B(n_8),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2105),
.A2(n_9),
.B(n_10),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2171),
.B(n_9),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2011),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1892),
.B(n_9),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_1881),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2106),
.A2(n_10),
.B(n_11),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1894),
.B(n_10),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2029),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_1880),
.B(n_12),
.Y(n_2361)
);

AOI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2106),
.A2(n_11),
.B(n_12),
.Y(n_2362)
);

OAI321xp33_ASAP7_75t_L g2363 ( 
.A1(n_2063),
.A2(n_14),
.A3(n_16),
.B1(n_11),
.B2(n_13),
.C(n_15),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1894),
.B(n_13),
.Y(n_2364)
);

A2O1A1Ixp33_ASAP7_75t_L g2365 ( 
.A1(n_2110),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2138),
.A2(n_14),
.B(n_15),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1895),
.B(n_16),
.Y(n_2367)
);

OAI21xp5_ASAP7_75t_L g2368 ( 
.A1(n_2060),
.A2(n_16),
.B(n_17),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2138),
.A2(n_17),
.B(n_18),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_1995),
.A2(n_2001),
.B(n_1899),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2132),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1895),
.B(n_19),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_1898),
.A2(n_19),
.B(n_20),
.Y(n_2373)
);

AOI21xp33_ASAP7_75t_L g2374 ( 
.A1(n_2015),
.A2(n_20),
.B(n_21),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1946),
.B(n_21),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1919),
.B(n_21),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2040),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1946),
.B(n_22),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_1902),
.A2(n_22),
.B(n_23),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1910),
.Y(n_2380)
);

NOR3xp33_ASAP7_75t_L g2381 ( 
.A(n_2045),
.B(n_24),
.C(n_23),
.Y(n_2381)
);

NOR2xp67_ASAP7_75t_L g2382 ( 
.A(n_2170),
.B(n_22),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_1906),
.A2(n_23),
.B(n_24),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1948),
.B(n_25),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_1948),
.B(n_25),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1939),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2047),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_1907),
.A2(n_25),
.B(n_26),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1900),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_1966),
.B(n_26),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2114),
.B(n_27),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_1908),
.A2(n_1914),
.B(n_1909),
.Y(n_2392)
);

AOI33xp33_ASAP7_75t_L g2393 ( 
.A1(n_2018),
.A2(n_28),
.A3(n_30),
.B1(n_26),
.B2(n_27),
.B3(n_29),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1966),
.B(n_27),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_1904),
.B(n_28),
.Y(n_2395)
);

BUFx8_ASAP7_75t_L g2396 ( 
.A(n_1929),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_1881),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2022),
.A2(n_29),
.B(n_30),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2139),
.B(n_30),
.Y(n_2399)
);

BUFx4f_ASAP7_75t_L g2400 ( 
.A(n_1929),
.Y(n_2400)
);

OAI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_1872),
.A2(n_2054),
.B(n_2052),
.Y(n_2401)
);

A2O1A1Ixp33_ASAP7_75t_L g2402 ( 
.A1(n_2118),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1901),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_1924),
.A2(n_31),
.B(n_32),
.Y(n_2404)
);

AOI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_1927),
.A2(n_31),
.B(n_33),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2049),
.Y(n_2406)
);

BUFx3_ASAP7_75t_L g2407 ( 
.A(n_1886),
.Y(n_2407)
);

NOR2xp67_ASAP7_75t_L g2408 ( 
.A(n_2174),
.B(n_34),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_1925),
.B(n_34),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_1930),
.A2(n_35),
.B(n_36),
.Y(n_2410)
);

NOR3xp33_ASAP7_75t_L g2411 ( 
.A(n_1933),
.B(n_37),
.C(n_36),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_1896),
.B(n_35),
.Y(n_2412)
);

OAI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_1872),
.A2(n_35),
.B(n_36),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2028),
.B(n_37),
.Y(n_2414)
);

OAI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2127),
.A2(n_37),
.B(n_38),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2120),
.B(n_38),
.Y(n_2416)
);

AOI21x1_ASAP7_75t_L g2417 ( 
.A1(n_2162),
.A2(n_38),
.B(n_39),
.Y(n_2417)
);

BUFx6f_ASAP7_75t_L g2418 ( 
.A(n_2011),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_1997),
.Y(n_2419)
);

INVx2_ASAP7_75t_SL g2420 ( 
.A(n_1967),
.Y(n_2420)
);

O2A1O1Ixp33_ASAP7_75t_L g2421 ( 
.A1(n_1870),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_2421)
);

AOI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_1981),
.A2(n_40),
.B(n_41),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2014),
.B(n_40),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_1991),
.A2(n_41),
.B(n_42),
.Y(n_2424)
);

AO21x1_ASAP7_75t_L g2425 ( 
.A1(n_1870),
.A2(n_136),
.B(n_135),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_1912),
.B(n_42),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_1874),
.B(n_43),
.Y(n_2427)
);

OAI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2150),
.A2(n_43),
.B(n_44),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1992),
.B(n_44),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_1886),
.B(n_45),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_1976),
.A2(n_45),
.B(n_46),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2051),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2037),
.B(n_46),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2151),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_1987),
.A2(n_47),
.B(n_49),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2075),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_1988),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_1923),
.B(n_50),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2048),
.B(n_49),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2100),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2152),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2104),
.Y(n_2442)
);

AO21x1_ASAP7_75t_L g2443 ( 
.A1(n_1988),
.A2(n_140),
.B(n_139),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2056),
.B(n_51),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_1947),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2107),
.B(n_52),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_1861),
.A2(n_51),
.B(n_52),
.Y(n_2447)
);

OAI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2154),
.A2(n_52),
.B(n_53),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2178),
.A2(n_53),
.B(n_54),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2012),
.A2(n_53),
.B(n_54),
.Y(n_2450)
);

OAI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2072),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2451)
);

O2A1O1Ixp5_ASAP7_75t_SL g2452 ( 
.A1(n_1936),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2107),
.B(n_57),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2017),
.B(n_55),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2165),
.Y(n_2455)
);

AOI22xp5_ASAP7_75t_L g2456 ( 
.A1(n_2026),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_1998),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2163),
.B(n_59),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2019),
.B(n_58),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_1998),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_1937),
.B(n_58),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2073),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_2186),
.A2(n_59),
.B(n_60),
.Y(n_2463)
);

OAI21xp33_ASAP7_75t_L g2464 ( 
.A1(n_1916),
.A2(n_60),
.B(n_61),
.Y(n_2464)
);

OAI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2187),
.A2(n_61),
.B(n_62),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2023),
.B(n_62),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_1922),
.B(n_61),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2059),
.A2(n_63),
.B(n_64),
.Y(n_2468)
);

AOI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2064),
.A2(n_63),
.B(n_64),
.Y(n_2469)
);

OAI22xp5_ASAP7_75t_L g2470 ( 
.A1(n_2184),
.A2(n_2177),
.B1(n_2082),
.B2(n_2083),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2020),
.Y(n_2471)
);

AOI21x1_ASAP7_75t_L g2472 ( 
.A1(n_2176),
.A2(n_2181),
.B(n_2180),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2074),
.B(n_64),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_1882),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2078),
.B(n_63),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2088),
.B(n_65),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2081),
.B(n_65),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2032),
.B(n_66),
.Y(n_2478)
);

AOI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2089),
.A2(n_65),
.B(n_66),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2094),
.B(n_2038),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2032),
.B(n_68),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1977),
.B(n_1958),
.Y(n_2482)
);

AOI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2006),
.A2(n_67),
.B(n_68),
.Y(n_2483)
);

INVx2_ASAP7_75t_SL g2484 ( 
.A(n_1873),
.Y(n_2484)
);

A2O1A1Ixp33_ASAP7_75t_L g2485 ( 
.A1(n_1935),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_2485)
);

INVxp67_ASAP7_75t_L g2486 ( 
.A(n_2039),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1990),
.Y(n_2487)
);

INVx3_ASAP7_75t_L g2488 ( 
.A(n_1953),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_1972),
.B(n_70),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2116),
.B(n_70),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2042),
.B(n_72),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2067),
.B(n_72),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2166),
.B(n_72),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2167),
.B(n_73),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2032),
.B(n_75),
.Y(n_2495)
);

OAI22xp5_ASAP7_75t_L g2496 ( 
.A1(n_2021),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_2496)
);

A2O1A1Ixp33_ASAP7_75t_L g2497 ( 
.A1(n_1952),
.A2(n_77),
.B(n_74),
.C(n_76),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2115),
.A2(n_2125),
.B(n_1875),
.Y(n_2498)
);

OAI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2021),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2020),
.A2(n_78),
.B(n_79),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2076),
.B(n_80),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_1993),
.B(n_81),
.Y(n_2502)
);

OR2x2_ASAP7_75t_L g2503 ( 
.A(n_2119),
.B(n_81),
.Y(n_2503)
);

O2A1O1Ixp5_ASAP7_75t_L g2504 ( 
.A1(n_1944),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2000),
.B(n_2003),
.Y(n_2505)
);

NOR2x1p5_ASAP7_75t_L g2506 ( 
.A(n_2071),
.B(n_82),
.Y(n_2506)
);

AOI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_2020),
.A2(n_82),
.B(n_83),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2131),
.A2(n_84),
.B(n_85),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2145),
.B(n_85),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2133),
.A2(n_86),
.B(n_87),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2140),
.A2(n_86),
.B(n_87),
.Y(n_2511)
);

AOI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2131),
.A2(n_86),
.B(n_87),
.Y(n_2512)
);

CKINVDCx10_ASAP7_75t_R g2513 ( 
.A(n_1960),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_1917),
.B(n_88),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_1918),
.B(n_88),
.Y(n_2515)
);

AOI22xp5_ASAP7_75t_L g2516 ( 
.A1(n_2179),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2516)
);

HB1xp67_ASAP7_75t_L g2517 ( 
.A(n_1953),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2009),
.B(n_89),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2030),
.B(n_89),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_SL g2520 ( 
.A(n_2142),
.B(n_90),
.C(n_91),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2031),
.B(n_90),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2036),
.B(n_1964),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2032),
.B(n_92),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2131),
.A2(n_91),
.B(n_92),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1974),
.B(n_93),
.Y(n_2525)
);

NOR2xp67_ASAP7_75t_L g2526 ( 
.A(n_1926),
.B(n_2035),
.Y(n_2526)
);

NOR2xp67_ASAP7_75t_L g2527 ( 
.A(n_2035),
.B(n_93),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2087),
.Y(n_2528)
);

OAI21xp5_ASAP7_75t_L g2529 ( 
.A1(n_2185),
.A2(n_94),
.B(n_95),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2144),
.B(n_94),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2090),
.Y(n_2531)
);

AOI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2141),
.A2(n_95),
.B(n_96),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2095),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2144),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2136),
.B(n_2153),
.Y(n_2535)
);

OAI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2141),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2159),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_1996),
.Y(n_2538)
);

OAI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2044),
.A2(n_96),
.B(n_97),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_1999),
.B(n_99),
.Y(n_2540)
);

NOR2x1_ASAP7_75t_L g2541 ( 
.A(n_2123),
.B(n_100),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2137),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2175),
.B(n_100),
.Y(n_2543)
);

AOI21xp5_ASAP7_75t_L g2544 ( 
.A1(n_2141),
.A2(n_100),
.B(n_101),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_L g2545 ( 
.A(n_2050),
.B(n_101),
.Y(n_2545)
);

BUFx3_ASAP7_75t_L g2546 ( 
.A(n_2137),
.Y(n_2546)
);

AOI21xp5_ASAP7_75t_L g2547 ( 
.A1(n_2057),
.A2(n_101),
.B(n_102),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2032),
.B(n_102),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2172),
.B(n_102),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2172),
.B(n_103),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2172),
.B(n_104),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2172),
.B(n_103),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2172),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_1885),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_1911),
.Y(n_2555)
);

HB1xp67_ASAP7_75t_L g2556 ( 
.A(n_1911),
.Y(n_2556)
);

AOI21x1_ASAP7_75t_L g2557 ( 
.A1(n_1982),
.A2(n_106),
.B(n_107),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2008),
.B(n_106),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_1866),
.B(n_107),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_1866),
.B(n_107),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_1941),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_1877),
.B(n_108),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_1866),
.B(n_108),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1941),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_1903),
.B(n_109),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_1877),
.B(n_110),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_1866),
.B(n_109),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2024),
.A2(n_110),
.B(n_111),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_1893),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2569)
);

O2A1O1Ixp33_ASAP7_75t_L g2570 ( 
.A1(n_2024),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1941),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2024),
.A2(n_112),
.B(n_113),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_1893),
.B(n_114),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2024),
.A2(n_114),
.B(n_115),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_1903),
.B(n_114),
.Y(n_2575)
);

OAI321xp33_ASAP7_75t_L g2576 ( 
.A1(n_2093),
.A2(n_117),
.A3(n_119),
.B1(n_115),
.B2(n_116),
.C(n_118),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_1877),
.B(n_116),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_1877),
.B(n_116),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2024),
.A2(n_115),
.B(n_117),
.Y(n_2579)
);

AOI21xp5_ASAP7_75t_L g2580 ( 
.A1(n_2024),
.A2(n_119),
.B(n_120),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2034),
.Y(n_2581)
);

INVxp67_ASAP7_75t_L g2582 ( 
.A(n_1893),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1941),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_1893),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_1866),
.B(n_119),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_1866),
.B(n_120),
.Y(n_2586)
);

OAI21xp33_ASAP7_75t_L g2587 ( 
.A1(n_2013),
.A2(n_120),
.B(n_121),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_1866),
.B(n_121),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_1893),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2589)
);

NAND2x1_ASAP7_75t_L g2590 ( 
.A(n_2137),
.B(n_123),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_1893),
.B(n_124),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_1893),
.B(n_124),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_1866),
.B(n_125),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_1903),
.B(n_125),
.Y(n_2594)
);

CKINVDCx10_ASAP7_75t_R g2595 ( 
.A(n_2065),
.Y(n_2595)
);

AOI21x1_ASAP7_75t_L g2596 ( 
.A1(n_2135),
.A2(n_125),
.B(n_126),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2007),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2024),
.A2(n_126),
.B(n_127),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_1866),
.B(n_126),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_1941),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2034),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_1941),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_1866),
.B(n_127),
.Y(n_2603)
);

NAND2x1p5_ASAP7_75t_L g2604 ( 
.A(n_2061),
.B(n_127),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_1866),
.B(n_128),
.Y(n_2605)
);

AOI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2024),
.A2(n_128),
.B(n_129),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2024),
.A2(n_128),
.B(n_129),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_1941),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2034),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2034),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2024),
.A2(n_130),
.B(n_132),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1941),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_1941),
.Y(n_2613)
);

A2O1A1Ixp33_ASAP7_75t_L g2614 ( 
.A1(n_2024),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2024),
.A2(n_132),
.B(n_133),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_1941),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_1866),
.B(n_134),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_1893),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2209),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2218),
.A2(n_134),
.B(n_144),
.Y(n_2620)
);

O2A1O1Ixp33_ASAP7_75t_L g2621 ( 
.A1(n_2344),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2317),
.B(n_146),
.Y(n_2622)
);

CKINVDCx14_ASAP7_75t_R g2623 ( 
.A(n_2296),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2233),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_L g2625 ( 
.A(n_2284),
.B(n_147),
.Y(n_2625)
);

OAI22x1_ASAP7_75t_L g2626 ( 
.A1(n_2562),
.A2(n_150),
.B1(n_151),
.B2(n_149),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2195),
.B(n_148),
.Y(n_2627)
);

A2O1A1Ixp33_ASAP7_75t_L g2628 ( 
.A1(n_2370),
.A2(n_155),
.B(n_149),
.C(n_154),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2581),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2317),
.B(n_154),
.Y(n_2630)
);

A2O1A1Ixp33_ASAP7_75t_L g2631 ( 
.A1(n_2370),
.A2(n_2392),
.B(n_2316),
.C(n_2221),
.Y(n_2631)
);

OAI221xp5_ASAP7_75t_L g2632 ( 
.A1(n_2319),
.A2(n_766),
.B1(n_767),
.B2(n_765),
.C(n_764),
.Y(n_2632)
);

NAND2x1p5_ASAP7_75t_L g2633 ( 
.A(n_2306),
.B(n_156),
.Y(n_2633)
);

AOI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2218),
.A2(n_156),
.B(n_157),
.Y(n_2634)
);

AOI21xp5_ASAP7_75t_L g2635 ( 
.A1(n_2392),
.A2(n_157),
.B(n_158),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_L g2636 ( 
.A(n_2462),
.B(n_158),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2601),
.B(n_2609),
.Y(n_2637)
);

O2A1O1Ixp33_ASAP7_75t_L g2638 ( 
.A1(n_2336),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2610),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2201),
.B(n_160),
.Y(n_2640)
);

NOR2xp67_ASAP7_75t_SL g2641 ( 
.A(n_2279),
.B(n_162),
.Y(n_2641)
);

A2O1A1Ixp33_ASAP7_75t_L g2642 ( 
.A1(n_2587),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_2642)
);

INVx2_ASAP7_75t_SL g2643 ( 
.A(n_2595),
.Y(n_2643)
);

OAI22xp33_ASAP7_75t_L g2644 ( 
.A1(n_2200),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2644)
);

HB1xp67_ASAP7_75t_L g2645 ( 
.A(n_2584),
.Y(n_2645)
);

AOI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2252),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2646)
);

AOI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2304),
.A2(n_168),
.B(n_169),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_SL g2648 ( 
.A(n_2315),
.B(n_168),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2245),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2256),
.Y(n_2650)
);

OAI21x1_ASAP7_75t_L g2651 ( 
.A1(n_2260),
.A2(n_169),
.B(n_170),
.Y(n_2651)
);

OAI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2197),
.A2(n_175),
.B1(n_171),
.B2(n_173),
.Y(n_2652)
);

INVx5_ASAP7_75t_L g2653 ( 
.A(n_2331),
.Y(n_2653)
);

OR2x6_ASAP7_75t_SL g2654 ( 
.A(n_2419),
.B(n_769),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_SL g2655 ( 
.A1(n_2562),
.A2(n_2430),
.B1(n_2331),
.B2(n_2416),
.Y(n_2655)
);

HB1xp67_ASAP7_75t_L g2656 ( 
.A(n_2618),
.Y(n_2656)
);

OAI22x1_ASAP7_75t_L g2657 ( 
.A1(n_2430),
.A2(n_180),
.B1(n_181),
.B2(n_178),
.Y(n_2657)
);

O2A1O1Ixp33_ASAP7_75t_L g2658 ( 
.A1(n_2470),
.A2(n_180),
.B(n_177),
.C(n_178),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_2396),
.Y(n_2659)
);

INVx1_ASAP7_75t_SL g2660 ( 
.A(n_2604),
.Y(n_2660)
);

OR2x6_ASAP7_75t_L g2661 ( 
.A(n_2251),
.B(n_177),
.Y(n_2661)
);

OA21x2_ASAP7_75t_L g2662 ( 
.A1(n_2227),
.A2(n_181),
.B(n_182),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2193),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2312),
.B(n_182),
.Y(n_2664)
);

O2A1O1Ixp33_ASAP7_75t_SL g2665 ( 
.A1(n_2213),
.A2(n_186),
.B(n_183),
.C(n_184),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2205),
.Y(n_2666)
);

OAI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2202),
.A2(n_187),
.B1(n_183),
.B2(n_186),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2455),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2246),
.Y(n_2669)
);

AO32x1_ASAP7_75t_L g2670 ( 
.A1(n_2437),
.A2(n_190),
.A3(n_188),
.B1(n_189),
.B2(n_192),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_2246),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2192),
.Y(n_2672)
);

AND2x6_ASAP7_75t_L g2673 ( 
.A(n_2546),
.B(n_2247),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2400),
.B(n_188),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2304),
.A2(n_192),
.B(n_193),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_2582),
.B(n_2226),
.Y(n_2676)
);

O2A1O1Ixp33_ASAP7_75t_SL g2677 ( 
.A1(n_2343),
.A2(n_2590),
.B(n_2322),
.C(n_2267),
.Y(n_2677)
);

INVx3_ASAP7_75t_L g2678 ( 
.A(n_2247),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2561),
.Y(n_2679)
);

OAI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2207),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_2680)
);

CKINVDCx20_ASAP7_75t_R g2681 ( 
.A(n_2597),
.Y(n_2681)
);

HB1xp67_ASAP7_75t_L g2682 ( 
.A(n_2229),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2564),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2298),
.B(n_195),
.Y(n_2684)
);

NOR2xp67_ASAP7_75t_SL g2685 ( 
.A(n_2251),
.B(n_197),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2407),
.B(n_198),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2571),
.B(n_198),
.Y(n_2687)
);

OAI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2559),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2399),
.B(n_199),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2573),
.B(n_201),
.Y(n_2690)
);

O2A1O1Ixp33_ASAP7_75t_L g2691 ( 
.A1(n_2480),
.A2(n_2473),
.B(n_2497),
.C(n_2566),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2457),
.B(n_204),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2591),
.B(n_206),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2583),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2592),
.B(n_206),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2600),
.B(n_2602),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2285),
.A2(n_207),
.B(n_208),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2608),
.B(n_207),
.Y(n_2698)
);

CKINVDCx14_ASAP7_75t_R g2699 ( 
.A(n_2331),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2612),
.Y(n_2700)
);

A2O1A1Ixp33_ASAP7_75t_SL g2701 ( 
.A1(n_2477),
.A2(n_211),
.B(n_208),
.C(n_210),
.Y(n_2701)
);

O2A1O1Ixp33_ASAP7_75t_L g2702 ( 
.A1(n_2577),
.A2(n_213),
.B(n_210),
.C(n_212),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_L g2703 ( 
.A(n_2460),
.B(n_212),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2613),
.B(n_213),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2414),
.B(n_215),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2306),
.Y(n_2706)
);

BUFx6f_ASAP7_75t_L g2707 ( 
.A(n_2193),
.Y(n_2707)
);

CKINVDCx6p67_ASAP7_75t_R g2708 ( 
.A(n_2326),
.Y(n_2708)
);

BUFx6f_ASAP7_75t_L g2709 ( 
.A(n_2193),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2616),
.B(n_216),
.Y(n_2710)
);

NOR2xp33_ASAP7_75t_SL g2711 ( 
.A(n_2542),
.B(n_216),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2486),
.B(n_217),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2309),
.B(n_218),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2236),
.A2(n_218),
.B(n_219),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2482),
.B(n_219),
.Y(n_2715)
);

O2A1O1Ixp5_ASAP7_75t_L g2716 ( 
.A1(n_2232),
.A2(n_2289),
.B(n_2297),
.C(n_2295),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2259),
.B(n_220),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_L g2718 ( 
.A1(n_2238),
.A2(n_220),
.B(n_221),
.Y(n_2718)
);

NOR2x1_ASAP7_75t_L g2719 ( 
.A(n_2326),
.B(n_221),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2261),
.Y(n_2720)
);

BUFx4f_ASAP7_75t_L g2721 ( 
.A(n_2604),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2423),
.B(n_222),
.Y(n_2722)
);

BUFx3_ASAP7_75t_L g2723 ( 
.A(n_2396),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2513),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2210),
.A2(n_222),
.B(n_223),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_2411),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2560),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_2727)
);

OR2x2_ASAP7_75t_L g2728 ( 
.A(n_2191),
.B(n_2198),
.Y(n_2728)
);

INVxp67_ASAP7_75t_SL g2729 ( 
.A(n_2192),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2223),
.B(n_228),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2441),
.Y(n_2731)
);

INVx3_ASAP7_75t_L g2732 ( 
.A(n_2261),
.Y(n_2732)
);

CKINVDCx11_ASAP7_75t_R g2733 ( 
.A(n_2262),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2348),
.B(n_228),
.Y(n_2734)
);

OAI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2196),
.A2(n_2204),
.B1(n_2292),
.B2(n_2503),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2257),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2380),
.Y(n_2737)
);

HB1xp67_ASAP7_75t_L g2738 ( 
.A(n_2352),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2386),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2354),
.B(n_229),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2389),
.B(n_229),
.Y(n_2741)
);

OAI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2563),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_2742)
);

AO22x1_ASAP7_75t_L g2743 ( 
.A1(n_2352),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_2743)
);

OAI21xp5_ASAP7_75t_L g2744 ( 
.A1(n_2327),
.A2(n_233),
.B(n_234),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2403),
.Y(n_2745)
);

AND3x2_ASAP7_75t_L g2746 ( 
.A(n_2264),
.B(n_234),
.C(n_237),
.Y(n_2746)
);

O2A1O1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2578),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2400),
.B(n_238),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2257),
.B(n_240),
.Y(n_2749)
);

AOI21xp5_ASAP7_75t_L g2750 ( 
.A1(n_2190),
.A2(n_241),
.B(n_243),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2416),
.B(n_241),
.Y(n_2751)
);

BUFx3_ASAP7_75t_L g2752 ( 
.A(n_2445),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2527),
.Y(n_2753)
);

A2O1A1Ixp33_ASAP7_75t_L g2754 ( 
.A1(n_2510),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_L g2755 ( 
.A1(n_2190),
.A2(n_2216),
.B(n_2194),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2567),
.B(n_245),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2451),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2280),
.Y(n_2758)
);

O2A1O1Ixp33_ASAP7_75t_L g2759 ( 
.A1(n_2374),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2585),
.B(n_250),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2586),
.B(n_250),
.Y(n_2761)
);

AO22x1_ASAP7_75t_L g2762 ( 
.A1(n_2381),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_SL g2763 ( 
.A(n_2199),
.B(n_251),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2294),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2502),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2382),
.B(n_2408),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2321),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2588),
.B(n_252),
.Y(n_2768)
);

OAI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2593),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2769)
);

BUFx2_ASAP7_75t_SL g2770 ( 
.A(n_2217),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2599),
.B(n_254),
.Y(n_2771)
);

OR2x6_ASAP7_75t_SL g2772 ( 
.A(n_2496),
.B(n_255),
.Y(n_2772)
);

A2O1A1Ixp33_ASAP7_75t_SL g2773 ( 
.A1(n_2368),
.A2(n_259),
.B(n_256),
.C(n_258),
.Y(n_2773)
);

OAI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2603),
.A2(n_260),
.B1(n_256),
.B2(n_259),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2335),
.B(n_260),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_2323),
.A2(n_264),
.B1(n_261),
.B2(n_262),
.Y(n_2776)
);

AO32x2_ASAP7_75t_L g2777 ( 
.A1(n_2536),
.A2(n_265),
.A3(n_262),
.B1(n_264),
.B2(n_266),
.Y(n_2777)
);

A2O1A1Ixp33_ASAP7_75t_L g2778 ( 
.A1(n_2510),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2376),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2263),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2328),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2393),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_2272),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2511),
.A2(n_271),
.B(n_269),
.C(n_270),
.Y(n_2784)
);

AOI21xp5_ASAP7_75t_L g2785 ( 
.A1(n_2216),
.A2(n_272),
.B(n_273),
.Y(n_2785)
);

INVxp67_ASAP7_75t_SL g2786 ( 
.A(n_2242),
.Y(n_2786)
);

INVx4_ASAP7_75t_L g2787 ( 
.A(n_2262),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2605),
.A2(n_275),
.B1(n_272),
.B2(n_274),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2258),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2194),
.A2(n_275),
.B(n_277),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2334),
.Y(n_2791)
);

OR2x6_ASAP7_75t_L g2792 ( 
.A(n_2262),
.B(n_277),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2617),
.B(n_2461),
.Y(n_2793)
);

AO32x2_ASAP7_75t_L g2794 ( 
.A1(n_2499),
.A2(n_280),
.A3(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2265),
.B(n_278),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2269),
.B(n_279),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2327),
.B(n_280),
.Y(n_2797)
);

O2A1O1Ixp5_ASAP7_75t_L g2798 ( 
.A1(n_2289),
.A2(n_285),
.B(n_281),
.C(n_283),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2493),
.B(n_283),
.Y(n_2799)
);

NAND2x1p5_ASAP7_75t_L g2800 ( 
.A(n_2282),
.B(n_285),
.Y(n_2800)
);

HB1xp67_ASAP7_75t_L g2801 ( 
.A(n_2346),
.Y(n_2801)
);

NOR3xp33_ASAP7_75t_L g2802 ( 
.A(n_2520),
.B(n_2391),
.C(n_2363),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2329),
.B(n_287),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2277),
.B(n_2286),
.Y(n_2804)
);

O2A1O1Ixp33_ASAP7_75t_SL g2805 ( 
.A1(n_2320),
.A2(n_2249),
.B(n_2240),
.C(n_2478),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2329),
.B(n_288),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2345),
.B(n_289),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_SL g2808 ( 
.A(n_2206),
.B(n_289),
.Y(n_2808)
);

INVxp67_ASAP7_75t_SL g2809 ( 
.A(n_2206),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2287),
.B(n_290),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2347),
.B(n_291),
.Y(n_2811)
);

A2O1A1Ixp33_ASAP7_75t_L g2812 ( 
.A1(n_2483),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_2812)
);

AND2x4_ASAP7_75t_L g2813 ( 
.A(n_2281),
.B(n_293),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_2506),
.Y(n_2814)
);

O2A1O1Ixp33_ASAP7_75t_L g2815 ( 
.A1(n_2466),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_2815)
);

A2O1A1Ixp33_ASAP7_75t_L g2816 ( 
.A1(n_2404),
.A2(n_299),
.B(n_296),
.C(n_297),
.Y(n_2816)
);

NAND3xp33_ASAP7_75t_L g2817 ( 
.A(n_2452),
.B(n_299),
.C(n_300),
.Y(n_2817)
);

NOR2x1_ASAP7_75t_SL g2818 ( 
.A(n_2206),
.B(n_300),
.Y(n_2818)
);

NAND2x1p5_ASAP7_75t_L g2819 ( 
.A(n_2318),
.B(n_301),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2351),
.A2(n_304),
.B1(n_301),
.B2(n_302),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2565),
.B(n_305),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2487),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2356),
.B(n_305),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2530),
.Y(n_2824)
);

A2O1A1Ixp33_ASAP7_75t_L g2825 ( 
.A1(n_2405),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_2825)
);

A2O1A1Ixp33_ASAP7_75t_L g2826 ( 
.A1(n_2405),
.A2(n_2410),
.B(n_2424),
.C(n_2422),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2189),
.A2(n_307),
.B(n_308),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2349),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2350),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2360),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2420),
.Y(n_2831)
);

OAI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2359),
.A2(n_312),
.B1(n_309),
.B2(n_310),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2377),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_2276),
.B(n_310),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2575),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2273),
.A2(n_312),
.B(n_313),
.Y(n_2836)
);

NOR2xp67_ASAP7_75t_L g2837 ( 
.A(n_2594),
.B(n_314),
.Y(n_2837)
);

NAND2xp33_ASAP7_75t_SL g2838 ( 
.A(n_2446),
.B(n_314),
.Y(n_2838)
);

INVx3_ASAP7_75t_L g2839 ( 
.A(n_2263),
.Y(n_2839)
);

INVx4_ASAP7_75t_L g2840 ( 
.A(n_2330),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2225),
.Y(n_2841)
);

HB1xp67_ASAP7_75t_L g2842 ( 
.A(n_2387),
.Y(n_2842)
);

O2A1O1Ixp5_ASAP7_75t_SL g2843 ( 
.A1(n_2481),
.A2(n_318),
.B(n_315),
.C(n_317),
.Y(n_2843)
);

NAND2xp33_ASAP7_75t_SL g2844 ( 
.A(n_2453),
.B(n_315),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_SL g2845 ( 
.A(n_2208),
.B(n_319),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2332),
.B(n_319),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2364),
.B(n_320),
.Y(n_2847)
);

INVx1_ASAP7_75t_SL g2848 ( 
.A(n_2237),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2367),
.B(n_320),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2372),
.B(n_322),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2514),
.B(n_322),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2406),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2515),
.B(n_323),
.Y(n_2853)
);

BUFx2_ASAP7_75t_L g2854 ( 
.A(n_2330),
.Y(n_2854)
);

HB1xp67_ASAP7_75t_L g2855 ( 
.A(n_2432),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2291),
.B(n_323),
.Y(n_2856)
);

INVx2_ASAP7_75t_SL g2857 ( 
.A(n_2535),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2427),
.Y(n_2858)
);

INVx3_ASAP7_75t_L g2859 ( 
.A(n_2357),
.Y(n_2859)
);

BUFx6f_ASAP7_75t_L g2860 ( 
.A(n_2208),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2301),
.B(n_324),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2313),
.B(n_2203),
.Y(n_2862)
);

AOI21xp33_ASAP7_75t_L g2863 ( 
.A1(n_2375),
.A2(n_2384),
.B(n_2378),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2401),
.B(n_324),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2266),
.A2(n_325),
.B(n_326),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2494),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_2517),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2456),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2208),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2436),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2222),
.A2(n_330),
.B(n_331),
.Y(n_2871)
);

OR2x6_ASAP7_75t_L g2872 ( 
.A(n_2421),
.B(n_332),
.Y(n_2872)
);

INVx3_ASAP7_75t_L g2873 ( 
.A(n_2357),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2385),
.B(n_333),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2525),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2440),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2235),
.B(n_334),
.Y(n_2877)
);

OAI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2390),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_L g2879 ( 
.A1(n_2492),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_2879)
);

OR2x2_ASAP7_75t_L g2880 ( 
.A(n_2337),
.B(n_338),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2302),
.B(n_339),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2394),
.B(n_341),
.Y(n_2882)
);

AOI21xp33_ASAP7_75t_L g2883 ( 
.A1(n_2412),
.A2(n_341),
.B(n_342),
.Y(n_2883)
);

AND2x4_ASAP7_75t_L g2884 ( 
.A(n_2537),
.B(n_342),
.Y(n_2884)
);

AOI22xp33_ASAP7_75t_L g2885 ( 
.A1(n_2491),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2464),
.A2(n_347),
.B1(n_344),
.B2(n_345),
.Y(n_2886)
);

O2A1O1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_2485),
.A2(n_350),
.B(n_348),
.C(n_349),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2395),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2397),
.Y(n_2889)
);

NOR3xp33_ASAP7_75t_SL g2890 ( 
.A(n_2576),
.B(n_351),
.C(n_352),
.Y(n_2890)
);

NOR3xp33_ASAP7_75t_SL g2891 ( 
.A(n_2467),
.B(n_351),
.C(n_352),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2303),
.B(n_353),
.Y(n_2892)
);

O2A1O1Ixp33_ASAP7_75t_L g2893 ( 
.A1(n_2361),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_2893)
);

HB1xp67_ASAP7_75t_L g2894 ( 
.A(n_2442),
.Y(n_2894)
);

OAI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2426),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2409),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_2896)
);

HB1xp67_ASAP7_75t_L g2897 ( 
.A(n_2548),
.Y(n_2897)
);

INVx3_ASAP7_75t_SL g2898 ( 
.A(n_2397),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_R g2899 ( 
.A(n_2557),
.B(n_358),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_2314),
.A2(n_360),
.B(n_361),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2305),
.B(n_361),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2569),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2308),
.B(n_2310),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_L g2904 ( 
.A(n_2214),
.Y(n_2904)
);

INVx4_ASAP7_75t_L g2905 ( 
.A(n_2214),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2413),
.B(n_363),
.Y(n_2906)
);

CKINVDCx14_ASAP7_75t_R g2907 ( 
.A(n_2490),
.Y(n_2907)
);

HB1xp67_ASAP7_75t_L g2908 ( 
.A(n_2549),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2540),
.A2(n_367),
.B1(n_364),
.B2(n_365),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2522),
.B(n_367),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2214),
.B(n_369),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2314),
.A2(n_369),
.B(n_370),
.Y(n_2912)
);

OA22x2_ASAP7_75t_L g2913 ( 
.A1(n_2589),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2324),
.A2(n_373),
.B(n_374),
.Y(n_2914)
);

CKINVDCx20_ASAP7_75t_R g2915 ( 
.A(n_2516),
.Y(n_2915)
);

INVx4_ASAP7_75t_L g2916 ( 
.A(n_2219),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2434),
.B(n_374),
.Y(n_2917)
);

OR2x6_ASAP7_75t_L g2918 ( 
.A(n_2431),
.B(n_375),
.Y(n_2918)
);

NAND3xp33_ASAP7_75t_L g2919 ( 
.A(n_2570),
.B(n_376),
.C(n_377),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2271),
.B(n_2274),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_SL g2921 ( 
.A1(n_2415),
.A2(n_379),
.B1(n_376),
.B2(n_378),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2278),
.B(n_378),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2324),
.A2(n_379),
.B(n_380),
.Y(n_2923)
);

AOI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2325),
.A2(n_2268),
.B(n_2498),
.Y(n_2924)
);

BUFx2_ASAP7_75t_L g2925 ( 
.A(n_2488),
.Y(n_2925)
);

OR2x6_ASAP7_75t_L g2926 ( 
.A(n_2431),
.B(n_380),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2325),
.A2(n_381),
.B(n_382),
.Y(n_2927)
);

NOR2xp33_ASAP7_75t_L g2928 ( 
.A(n_2283),
.B(n_381),
.Y(n_2928)
);

BUFx6f_ASAP7_75t_SL g2929 ( 
.A(n_2528),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2307),
.Y(n_2930)
);

OAI21xp5_ASAP7_75t_L g2931 ( 
.A1(n_2333),
.A2(n_2342),
.B(n_2341),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2288),
.B(n_383),
.Y(n_2932)
);

A2O1A1Ixp33_ASAP7_75t_L g2933 ( 
.A1(n_2410),
.A2(n_388),
.B(n_385),
.C(n_386),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2505),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2293),
.B(n_385),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2488),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2447),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_SL g2938 ( 
.A(n_2531),
.Y(n_2938)
);

NOR2xp33_ASAP7_75t_L g2939 ( 
.A(n_2299),
.B(n_388),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_SL g2940 ( 
.A(n_2219),
.B(n_392),
.Y(n_2940)
);

OAI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2333),
.A2(n_392),
.B(n_393),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_L g2942 ( 
.A(n_2300),
.B(n_393),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2429),
.B(n_394),
.Y(n_2943)
);

HB1xp67_ASAP7_75t_L g2944 ( 
.A(n_2550),
.Y(n_2944)
);

INVx4_ASAP7_75t_L g2945 ( 
.A(n_2219),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2250),
.A2(n_394),
.B(n_396),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2275),
.B(n_397),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2518),
.Y(n_2948)
);

CKINVDCx20_ASAP7_75t_R g2949 ( 
.A(n_2438),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2433),
.B(n_397),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2255),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2253),
.A2(n_398),
.B(n_399),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2239),
.B(n_399),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2275),
.B(n_400),
.Y(n_2954)
);

NOR2xp33_ASAP7_75t_R g2955 ( 
.A(n_2230),
.B(n_400),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2596),
.Y(n_2956)
);

OAI22xp5_ASAP7_75t_SL g2957 ( 
.A1(n_2371),
.A2(n_405),
.B1(n_402),
.B2(n_403),
.Y(n_2957)
);

AOI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2425),
.A2(n_406),
.B1(n_402),
.B2(n_405),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2275),
.B(n_407),
.Y(n_2959)
);

A2O1A1Ixp33_ASAP7_75t_SL g2960 ( 
.A1(n_2545),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_2960)
);

AOI22xp5_ASAP7_75t_L g2961 ( 
.A1(n_2443),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_2961)
);

O2A1O1Ixp33_ASAP7_75t_L g2962 ( 
.A1(n_2339),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2439),
.B(n_411),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2444),
.B(n_412),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2454),
.B(n_414),
.Y(n_2965)
);

OAI21xp33_ASAP7_75t_SL g2966 ( 
.A1(n_2428),
.A2(n_415),
.B(n_416),
.Y(n_2966)
);

AOI21x1_ASAP7_75t_L g2967 ( 
.A1(n_2472),
.A2(n_415),
.B(n_416),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2519),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2270),
.B(n_417),
.Y(n_2969)
);

NOR2xp33_ASAP7_75t_L g2970 ( 
.A(n_2290),
.B(n_417),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2459),
.B(n_418),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2338),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_SL g2973 ( 
.A(n_2338),
.B(n_418),
.Y(n_2973)
);

OR2x2_ASAP7_75t_L g2974 ( 
.A(n_2248),
.B(n_419),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2417),
.Y(n_2975)
);

INVx4_ASAP7_75t_L g2976 ( 
.A(n_2338),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2538),
.B(n_419),
.Y(n_2977)
);

O2A1O1Ixp33_ASAP7_75t_L g2978 ( 
.A1(n_2340),
.A2(n_422),
.B(n_420),
.C(n_421),
.Y(n_2978)
);

O2A1O1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2614),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_2979)
);

BUFx2_ASAP7_75t_L g2980 ( 
.A(n_2534),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2475),
.B(n_423),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2649),
.Y(n_2982)
);

AOI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_2631),
.A2(n_2418),
.B(n_2355),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2694),
.Y(n_2984)
);

O2A1O1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2793),
.A2(n_2402),
.B(n_2365),
.C(n_2521),
.Y(n_2985)
);

OAI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2691),
.A2(n_2802),
.B(n_2826),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2700),
.Y(n_2987)
);

INVxp67_ASAP7_75t_SL g2988 ( 
.A(n_2721),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2737),
.Y(n_2989)
);

NAND2x1p5_ASAP7_75t_L g2990 ( 
.A(n_2659),
.B(n_2541),
.Y(n_2990)
);

A2O1A1Ixp33_ASAP7_75t_L g2991 ( 
.A1(n_2721),
.A2(n_2448),
.B(n_2465),
.C(n_2568),
.Y(n_2991)
);

OA21x2_ASAP7_75t_L g2992 ( 
.A1(n_2755),
.A2(n_2369),
.B(n_2366),
.Y(n_2992)
);

NOR2xp33_ASAP7_75t_L g2993 ( 
.A(n_2907),
.B(n_2231),
.Y(n_2993)
);

AOI221x1_ASAP7_75t_L g2994 ( 
.A1(n_2626),
.A2(n_2657),
.B1(n_2785),
.B2(n_2634),
.C(n_2675),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2782),
.B(n_2422),
.Y(n_2995)
);

INVx2_ASAP7_75t_SL g2996 ( 
.A(n_2708),
.Y(n_2996)
);

A2O1A1Ixp33_ASAP7_75t_L g2997 ( 
.A1(n_2658),
.A2(n_2572),
.B(n_2574),
.C(n_2568),
.Y(n_2997)
);

INVx5_ASAP7_75t_L g2998 ( 
.A(n_2661),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2934),
.B(n_2424),
.Y(n_2999)
);

NAND2x1p5_ASAP7_75t_L g3000 ( 
.A(n_2723),
.B(n_2243),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2739),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2920),
.B(n_2373),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2841),
.B(n_2373),
.Y(n_3003)
);

AOI221x1_ASAP7_75t_L g3004 ( 
.A1(n_2647),
.A2(n_2362),
.B1(n_2358),
.B2(n_2353),
.C(n_2512),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2677),
.A2(n_2418),
.B(n_2355),
.Y(n_3005)
);

OA21x2_ASAP7_75t_L g3006 ( 
.A1(n_2716),
.A2(n_2529),
.B(n_2524),
.Y(n_3006)
);

BUFx2_ASAP7_75t_L g3007 ( 
.A(n_2653),
.Y(n_3007)
);

NAND3xp33_ASAP7_75t_SL g3008 ( 
.A(n_2955),
.B(n_2574),
.C(n_2572),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_L g3009 ( 
.A(n_2663),
.Y(n_3009)
);

AO31x2_ASAP7_75t_L g3010 ( 
.A1(n_2956),
.A2(n_2975),
.A3(n_2924),
.B(n_2937),
.Y(n_3010)
);

A2O1A1Ixp33_ASAP7_75t_L g3011 ( 
.A1(n_2638),
.A2(n_2580),
.B(n_2598),
.C(n_2579),
.Y(n_3011)
);

BUFx10_ASAP7_75t_L g3012 ( 
.A(n_2643),
.Y(n_3012)
);

AOI221xp5_ASAP7_75t_SL g3013 ( 
.A1(n_2735),
.A2(n_2398),
.B1(n_2388),
.B2(n_2383),
.C(n_2379),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2668),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2805),
.A2(n_2471),
.B(n_2212),
.Y(n_3015)
);

HB1xp67_ASAP7_75t_L g3016 ( 
.A(n_2682),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2655),
.B(n_2379),
.Y(n_3017)
);

AOI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2863),
.A2(n_2471),
.B(n_2552),
.Y(n_3018)
);

OAI21xp5_ASAP7_75t_L g3019 ( 
.A1(n_2858),
.A2(n_2504),
.B(n_2358),
.Y(n_3019)
);

A2O1A1Ixp33_ASAP7_75t_L g3020 ( 
.A1(n_2621),
.A2(n_2580),
.B(n_2598),
.C(n_2579),
.Y(n_3020)
);

OAI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2661),
.A2(n_2463),
.B1(n_2615),
.B2(n_2607),
.Y(n_3021)
);

NOR2xp67_ASAP7_75t_L g3022 ( 
.A(n_2653),
.B(n_2435),
.Y(n_3022)
);

BUFx8_ASAP7_75t_L g3023 ( 
.A(n_2929),
.Y(n_3023)
);

AOI21x1_ASAP7_75t_SL g3024 ( 
.A1(n_2864),
.A2(n_2543),
.B(n_2489),
.Y(n_3024)
);

AND2x6_ASAP7_75t_L g3025 ( 
.A(n_2660),
.B(n_2471),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2792),
.A2(n_2607),
.B1(n_2611),
.B2(n_2606),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2705),
.B(n_2606),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2745),
.B(n_2696),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2804),
.B(n_2509),
.Y(n_3029)
);

NOR2x1p5_ASAP7_75t_L g3030 ( 
.A(n_2672),
.B(n_2501),
.Y(n_3030)
);

INVx1_ASAP7_75t_SL g3031 ( 
.A(n_2752),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2679),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2786),
.A2(n_2234),
.B(n_2228),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2862),
.A2(n_2553),
.B(n_2476),
.Y(n_3034)
);

A2O1A1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2978),
.A2(n_2611),
.B(n_2615),
.C(n_2449),
.Y(n_3035)
);

BUFx12f_ASAP7_75t_L g3036 ( 
.A(n_2724),
.Y(n_3036)
);

A2O1A1Ixp33_ASAP7_75t_L g3037 ( 
.A1(n_2966),
.A2(n_2775),
.B(n_2887),
.C(n_2979),
.Y(n_3037)
);

INVx2_ASAP7_75t_SL g3038 ( 
.A(n_2736),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2683),
.B(n_2383),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2731),
.B(n_2388),
.Y(n_3040)
);

INVx5_ASAP7_75t_L g3041 ( 
.A(n_2661),
.Y(n_3041)
);

A2O1A1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_2962),
.A2(n_2449),
.B(n_2468),
.C(n_2450),
.Y(n_3042)
);

BUFx10_ASAP7_75t_L g3043 ( 
.A(n_2792),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2866),
.A2(n_2224),
.B(n_2495),
.Y(n_3044)
);

AOI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2808),
.A2(n_2551),
.B(n_2523),
.Y(n_3045)
);

AND2x4_ASAP7_75t_L g3046 ( 
.A(n_2653),
.B(n_2474),
.Y(n_3046)
);

BUFx2_ASAP7_75t_L g3047 ( 
.A(n_2729),
.Y(n_3047)
);

A2O1A1Ixp33_ASAP7_75t_L g3048 ( 
.A1(n_2744),
.A2(n_2450),
.B(n_2469),
.C(n_2468),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2857),
.B(n_2915),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2949),
.B(n_2533),
.Y(n_3050)
);

NAND2x1_ASAP7_75t_L g3051 ( 
.A(n_2673),
.B(n_2311),
.Y(n_3051)
);

OAI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2881),
.A2(n_2362),
.B(n_2353),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2779),
.B(n_2398),
.Y(n_3053)
);

NAND2xp33_ASAP7_75t_L g3054 ( 
.A(n_2673),
.B(n_2539),
.Y(n_3054)
);

OAI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2928),
.A2(n_2342),
.B(n_2341),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2808),
.A2(n_2211),
.B(n_2558),
.Y(n_3056)
);

AOI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2845),
.A2(n_2458),
.B(n_2532),
.Y(n_3057)
);

AOI22xp33_ASAP7_75t_L g3058 ( 
.A1(n_2872),
.A2(n_2469),
.B1(n_2479),
.B2(n_2435),
.Y(n_3058)
);

OAI21x1_ASAP7_75t_L g3059 ( 
.A1(n_2651),
.A2(n_2544),
.B(n_2507),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2629),
.Y(n_3060)
);

NOR2x1_ASAP7_75t_L g3061 ( 
.A(n_2792),
.B(n_2463),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2903),
.B(n_2479),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2822),
.Y(n_3063)
);

AOI22x1_ASAP7_75t_L g3064 ( 
.A1(n_2633),
.A2(n_2508),
.B1(n_2500),
.B2(n_2547),
.Y(n_3064)
);

OAI22xp5_ASAP7_75t_L g3065 ( 
.A1(n_2699),
.A2(n_2220),
.B1(n_2484),
.B2(n_2556),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2845),
.A2(n_2241),
.B(n_2215),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2663),
.Y(n_3067)
);

AO32x2_ASAP7_75t_L g3068 ( 
.A1(n_2957),
.A2(n_2526),
.A3(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_3068)
);

INVx4_ASAP7_75t_L g3069 ( 
.A(n_2672),
.Y(n_3069)
);

OAI22xp5_ASAP7_75t_L g3070 ( 
.A1(n_2772),
.A2(n_2534),
.B1(n_2254),
.B2(n_2554),
.Y(n_3070)
);

OAI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2939),
.A2(n_2244),
.B(n_2555),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2639),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2789),
.B(n_769),
.Y(n_3073)
);

OA22x2_ASAP7_75t_L g3074 ( 
.A1(n_2746),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_3074)
);

OAI21x1_ASAP7_75t_L g3075 ( 
.A1(n_2967),
.A2(n_427),
.B(n_428),
.Y(n_3075)
);

OAI21x1_ASAP7_75t_L g3076 ( 
.A1(n_2931),
.A2(n_2843),
.B(n_2809),
.Y(n_3076)
);

NAND2x1p5_ASAP7_75t_L g3077 ( 
.A(n_2706),
.B(n_768),
.Y(n_3077)
);

OAI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2942),
.A2(n_429),
.B(n_430),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2973),
.A2(n_430),
.B(n_432),
.Y(n_3079)
);

OAI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2906),
.A2(n_433),
.B(n_434),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2619),
.Y(n_3081)
);

CKINVDCx11_ASAP7_75t_R g3082 ( 
.A(n_2681),
.Y(n_3082)
);

INVx3_ASAP7_75t_L g3083 ( 
.A(n_2666),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2948),
.B(n_767),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2684),
.B(n_433),
.Y(n_3085)
);

A2O1A1Ixp33_ASAP7_75t_L g3086 ( 
.A1(n_2864),
.A2(n_436),
.B(n_434),
.C(n_435),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2624),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2835),
.B(n_435),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2919),
.A2(n_2763),
.B(n_2715),
.Y(n_3089)
);

OAI22x1_ASAP7_75t_L g3090 ( 
.A1(n_2800),
.A2(n_439),
.B1(n_436),
.B2(n_437),
.Y(n_3090)
);

INVx3_ASAP7_75t_L g3091 ( 
.A(n_2666),
.Y(n_3091)
);

BUFx3_ASAP7_75t_L g3092 ( 
.A(n_2733),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2676),
.B(n_2814),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2690),
.B(n_2693),
.Y(n_3094)
);

AOI21x1_ASAP7_75t_L g3095 ( 
.A1(n_2662),
.A2(n_439),
.B(n_440),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2973),
.A2(n_441),
.B(n_442),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2660),
.A2(n_443),
.B(n_445),
.Y(n_3097)
);

OAI22x1_ASAP7_75t_L g3098 ( 
.A1(n_2800),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_3098)
);

AO31x2_ASAP7_75t_L g3099 ( 
.A1(n_2628),
.A2(n_450),
.A3(n_447),
.B(n_449),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2650),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2713),
.B(n_447),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2637),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2791),
.Y(n_3103)
);

O2A1O1Ixp5_ASAP7_75t_SL g3104 ( 
.A1(n_2766),
.A2(n_452),
.B(n_449),
.C(n_451),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2695),
.B(n_2717),
.Y(n_3105)
);

INVxp67_ASAP7_75t_SL g3106 ( 
.A(n_2738),
.Y(n_3106)
);

NAND2x1p5_ASAP7_75t_L g3107 ( 
.A(n_2706),
.B(n_452),
.Y(n_3107)
);

BUFx6f_ASAP7_75t_L g3108 ( 
.A(n_2663),
.Y(n_3108)
);

OAI21x1_ASAP7_75t_L g3109 ( 
.A1(n_2865),
.A2(n_453),
.B(n_454),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2801),
.Y(n_3110)
);

AOI21xp5_ASAP7_75t_SL g3111 ( 
.A1(n_2687),
.A2(n_455),
.B(n_457),
.Y(n_3111)
);

OAI21x1_ASAP7_75t_L g3112 ( 
.A1(n_2662),
.A2(n_458),
.B(n_460),
.Y(n_3112)
);

O2A1O1Ixp33_ASAP7_75t_L g3113 ( 
.A1(n_2701),
.A2(n_2960),
.B(n_2751),
.C(n_2632),
.Y(n_3113)
);

AO31x2_ASAP7_75t_L g3114 ( 
.A1(n_2642),
.A2(n_463),
.A3(n_460),
.B(n_461),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_SL g3115 ( 
.A1(n_2687),
.A2(n_463),
.B(n_464),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_SL g3116 ( 
.A(n_2787),
.B(n_465),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2773),
.A2(n_466),
.B(n_467),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2824),
.A2(n_468),
.B(n_469),
.Y(n_3118)
);

OR2x6_ASAP7_75t_L g3119 ( 
.A(n_2633),
.B(n_470),
.Y(n_3119)
);

AND2x4_ASAP7_75t_L g3120 ( 
.A(n_2787),
.B(n_471),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2730),
.B(n_472),
.Y(n_3121)
);

BUFx2_ASAP7_75t_R g3122 ( 
.A(n_2654),
.Y(n_3122)
);

AOI221xp5_ASAP7_75t_SL g3123 ( 
.A1(n_2776),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.C(n_475),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2968),
.B(n_763),
.Y(n_3124)
);

AND2x4_ASAP7_75t_L g3125 ( 
.A(n_2669),
.B(n_476),
.Y(n_3125)
);

OAI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2635),
.A2(n_477),
.B(n_479),
.Y(n_3126)
);

INVxp67_ASAP7_75t_SL g3127 ( 
.A(n_2828),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2875),
.B(n_763),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2756),
.A2(n_479),
.B(n_480),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2760),
.A2(n_482),
.B(n_483),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_2842),
.B(n_483),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_2855),
.B(n_2894),
.Y(n_3132)
);

OAI22xp5_ASAP7_75t_L g3133 ( 
.A1(n_2872),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2761),
.A2(n_485),
.B(n_487),
.Y(n_3134)
);

AOI21xp33_ASAP7_75t_L g3135 ( 
.A1(n_2753),
.A2(n_487),
.B(n_488),
.Y(n_3135)
);

INVx1_ASAP7_75t_SL g3136 ( 
.A(n_2770),
.Y(n_3136)
);

A2O1A1Ixp33_ASAP7_75t_L g3137 ( 
.A1(n_2941),
.A2(n_491),
.B(n_489),
.C(n_490),
.Y(n_3137)
);

CKINVDCx8_ASAP7_75t_R g3138 ( 
.A(n_2783),
.Y(n_3138)
);

AO32x2_ASAP7_75t_L g3139 ( 
.A1(n_2957),
.A2(n_493),
.A3(n_489),
.B1(n_492),
.B2(n_495),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2758),
.Y(n_3140)
);

A2O1A1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_2815),
.A2(n_498),
.B(n_492),
.C(n_496),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2698),
.Y(n_3142)
);

BUFx3_ASAP7_75t_L g3143 ( 
.A(n_2898),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2698),
.Y(n_3144)
);

OAI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2919),
.A2(n_496),
.B(n_498),
.Y(n_3145)
);

BUFx3_ASAP7_75t_L g3146 ( 
.A(n_2831),
.Y(n_3146)
);

OAI21xp5_ASAP7_75t_L g3147 ( 
.A1(n_2856),
.A2(n_499),
.B(n_500),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2764),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2765),
.B(n_762),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2767),
.Y(n_3150)
);

O2A1O1Ixp5_ASAP7_75t_SL g3151 ( 
.A1(n_2664),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_3151)
);

OAI21x1_ASAP7_75t_L g3152 ( 
.A1(n_2620),
.A2(n_502),
.B(n_503),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2722),
.B(n_502),
.Y(n_3153)
);

CKINVDCx5p33_ASAP7_75t_R g3154 ( 
.A(n_2623),
.Y(n_3154)
);

O2A1O1Ixp33_ASAP7_75t_L g3155 ( 
.A1(n_2834),
.A2(n_506),
.B(n_504),
.C(n_505),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2781),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_2877),
.A2(n_507),
.B1(n_504),
.B2(n_506),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2799),
.B(n_507),
.Y(n_3158)
);

O2A1O1Ixp33_ASAP7_75t_SL g3159 ( 
.A1(n_2754),
.A2(n_510),
.B(n_508),
.C(n_509),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2645),
.B(n_2656),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2861),
.A2(n_508),
.B(n_510),
.Y(n_3161)
);

INVxp67_ASAP7_75t_SL g3162 ( 
.A(n_2813),
.Y(n_3162)
);

O2A1O1Ixp33_ASAP7_75t_L g3163 ( 
.A1(n_2795),
.A2(n_513),
.B(n_511),
.C(n_512),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_2872),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_3164)
);

AND2x4_ASAP7_75t_L g3165 ( 
.A(n_2669),
.B(n_514),
.Y(n_3165)
);

O2A1O1Ixp33_ASAP7_75t_SL g3166 ( 
.A1(n_2778),
.A2(n_517),
.B(n_514),
.C(n_516),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2768),
.A2(n_516),
.B(n_517),
.Y(n_3167)
);

OAI22x1_ASAP7_75t_L g3168 ( 
.A1(n_2819),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2636),
.B(n_761),
.Y(n_3169)
);

OAI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2892),
.A2(n_521),
.B(n_522),
.Y(n_3170)
);

OAI21x1_ASAP7_75t_L g3171 ( 
.A1(n_2798),
.A2(n_523),
.B(n_524),
.Y(n_3171)
);

AOI211x1_ASAP7_75t_L g3172 ( 
.A1(n_2743),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_3172)
);

AOI31xp67_ASAP7_75t_L g3173 ( 
.A1(n_2958),
.A2(n_530),
.A3(n_528),
.B(n_529),
.Y(n_3173)
);

AOI221xp5_ASAP7_75t_L g3174 ( 
.A1(n_2625),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.C(n_533),
.Y(n_3174)
);

AOI21x1_ASAP7_75t_L g3175 ( 
.A1(n_2897),
.A2(n_531),
.B(n_533),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_2728),
.B(n_534),
.Y(n_3176)
);

AO21x2_ASAP7_75t_L g3177 ( 
.A1(n_2899),
.A2(n_2817),
.B(n_2644),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2771),
.A2(n_534),
.B(n_535),
.Y(n_3178)
);

AOI21xp5_ASAP7_75t_L g3179 ( 
.A1(n_2874),
.A2(n_2882),
.B(n_2823),
.Y(n_3179)
);

A2O1A1Ixp33_ASAP7_75t_L g3180 ( 
.A1(n_2958),
.A2(n_537),
.B(n_535),
.C(n_536),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_2811),
.A2(n_2849),
.B(n_2847),
.Y(n_3181)
);

INVx1_ASAP7_75t_SL g3182 ( 
.A(n_2848),
.Y(n_3182)
);

INVx4_ASAP7_75t_L g3183 ( 
.A(n_2673),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2829),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2850),
.A2(n_536),
.B(n_537),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2830),
.Y(n_3186)
);

OAI21x1_ASAP7_75t_L g3187 ( 
.A1(n_2951),
.A2(n_538),
.B(n_539),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2833),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2851),
.A2(n_538),
.B(n_539),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2852),
.Y(n_3190)
);

AOI22xp33_ASAP7_75t_L g3191 ( 
.A1(n_2913),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2870),
.Y(n_3192)
);

O2A1O1Ixp5_ASAP7_75t_L g3193 ( 
.A1(n_2838),
.A2(n_545),
.B(n_543),
.C(n_544),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2876),
.Y(n_3194)
);

OAI21x1_ASAP7_75t_L g3195 ( 
.A1(n_2725),
.A2(n_543),
.B(n_545),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2704),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2689),
.B(n_547),
.Y(n_3197)
);

BUFx6f_ASAP7_75t_L g3198 ( 
.A(n_2707),
.Y(n_3198)
);

O2A1O1Ixp33_ASAP7_75t_SL g3199 ( 
.A1(n_2784),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_3199)
);

O2A1O1Ixp33_ASAP7_75t_SL g3200 ( 
.A1(n_2812),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2853),
.A2(n_552),
.B(n_553),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2813),
.B(n_2821),
.Y(n_3202)
);

AOI221x1_ASAP7_75t_L g3203 ( 
.A1(n_2817),
.A2(n_552),
.B1(n_553),
.B2(n_554),
.C(n_555),
.Y(n_3203)
);

OAI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2901),
.A2(n_554),
.B(n_555),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2710),
.Y(n_3205)
);

O2A1O1Ixp33_ASAP7_75t_SL g3206 ( 
.A1(n_2816),
.A2(n_558),
.B(n_556),
.C(n_557),
.Y(n_3206)
);

O2A1O1Ixp33_ASAP7_75t_L g3207 ( 
.A1(n_2796),
.A2(n_558),
.B(n_556),
.C(n_557),
.Y(n_3207)
);

AOI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2950),
.A2(n_559),
.B(n_560),
.Y(n_3208)
);

NAND2x1p5_ASAP7_75t_L g3209 ( 
.A(n_2685),
.B(n_760),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_2974),
.B(n_559),
.Y(n_3210)
);

AOI221x1_ASAP7_75t_L g3211 ( 
.A1(n_2714),
.A2(n_560),
.B1(n_562),
.B2(n_563),
.C(n_564),
.Y(n_3211)
);

AOI22xp5_ASAP7_75t_L g3212 ( 
.A1(n_2917),
.A2(n_565),
.B1(n_562),
.B2(n_564),
.Y(n_3212)
);

A2O1A1Ixp33_ASAP7_75t_L g3213 ( 
.A1(n_2961),
.A2(n_567),
.B(n_565),
.C(n_566),
.Y(n_3213)
);

A2O1A1Ixp33_ASAP7_75t_L g3214 ( 
.A1(n_2961),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_3214)
);

AOI221xp5_ASAP7_75t_SL g3215 ( 
.A1(n_2702),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.C(n_571),
.Y(n_3215)
);

AOI21x1_ASAP7_75t_L g3216 ( 
.A1(n_2908),
.A2(n_570),
.B(n_571),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2963),
.A2(n_572),
.B(n_573),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2929),
.B(n_574),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_2964),
.A2(n_574),
.B(n_575),
.Y(n_3219)
);

CKINVDCx5p33_ASAP7_75t_R g3220 ( 
.A(n_2938),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2910),
.B(n_575),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2965),
.A2(n_576),
.B(n_577),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2938),
.B(n_577),
.Y(n_3223)
);

AO21x1_ASAP7_75t_L g3224 ( 
.A1(n_2711),
.A2(n_578),
.B(n_579),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_2971),
.A2(n_579),
.B(n_580),
.Y(n_3225)
);

AO32x2_ASAP7_75t_L g3226 ( 
.A1(n_2878),
.A2(n_580),
.A3(n_582),
.B1(n_583),
.B2(n_584),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2918),
.Y(n_3227)
);

OAI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2922),
.A2(n_584),
.B(n_585),
.Y(n_3228)
);

AO31x2_ASAP7_75t_L g3229 ( 
.A1(n_2718),
.A2(n_585),
.A3(n_586),
.B(n_587),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2918),
.Y(n_3230)
);

NAND3x1_ASAP7_75t_L g3231 ( 
.A(n_2719),
.B(n_586),
.C(n_587),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_2790),
.A2(n_588),
.B(n_589),
.Y(n_3232)
);

A2O1A1Ixp33_ASAP7_75t_L g3233 ( 
.A1(n_2844),
.A2(n_590),
.B(n_592),
.C(n_593),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2692),
.B(n_760),
.Y(n_3234)
);

A2O1A1Ixp33_ASAP7_75t_L g3235 ( 
.A1(n_2868),
.A2(n_594),
.B(n_595),
.C(n_596),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_2981),
.A2(n_594),
.B(n_596),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2918),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_2943),
.A2(n_597),
.B(n_598),
.Y(n_3238)
);

OAI22x1_ASAP7_75t_L g3239 ( 
.A1(n_2819),
.A2(n_597),
.B1(n_599),
.B2(n_600),
.Y(n_3239)
);

AND2x4_ASAP7_75t_L g3240 ( 
.A(n_2671),
.B(n_600),
.Y(n_3240)
);

OAI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2932),
.A2(n_601),
.B(n_602),
.Y(n_3241)
);

AOI221xp5_ASAP7_75t_L g3242 ( 
.A1(n_2640),
.A2(n_601),
.B1(n_604),
.B2(n_607),
.C(n_609),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_2944),
.A2(n_610),
.B(n_611),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2741),
.Y(n_3244)
);

OA21x2_ASAP7_75t_L g3245 ( 
.A1(n_2827),
.A2(n_611),
.B(n_612),
.Y(n_3245)
);

OAI21x1_ASAP7_75t_L g3246 ( 
.A1(n_2697),
.A2(n_613),
.B(n_615),
.Y(n_3246)
);

INVx3_ASAP7_75t_L g3247 ( 
.A(n_2673),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_2750),
.A2(n_613),
.B(n_615),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2627),
.Y(n_3249)
);

O2A1O1Ixp33_ASAP7_75t_SL g3250 ( 
.A1(n_2825),
.A2(n_616),
.B(n_617),
.C(n_618),
.Y(n_3250)
);

AO31x2_ASAP7_75t_L g3251 ( 
.A1(n_2836),
.A2(n_616),
.A3(n_617),
.B(n_618),
.Y(n_3251)
);

AO31x2_ASAP7_75t_L g3252 ( 
.A1(n_2933),
.A2(n_620),
.A3(n_622),
.B(n_623),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2911),
.A2(n_622),
.B(n_623),
.Y(n_3253)
);

INVx3_ASAP7_75t_L g3254 ( 
.A(n_2840),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_2940),
.A2(n_624),
.B(n_625),
.Y(n_3255)
);

INVx5_ASAP7_75t_L g3256 ( 
.A(n_2707),
.Y(n_3256)
);

INVxp67_ASAP7_75t_L g3257 ( 
.A(n_2686),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3094),
.B(n_3105),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2982),
.Y(n_3259)
);

CKINVDCx6p67_ASAP7_75t_R g3260 ( 
.A(n_3082),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3014),
.Y(n_3261)
);

AOI22xp33_ASAP7_75t_L g3262 ( 
.A1(n_3029),
.A2(n_2926),
.B1(n_2977),
.B2(n_2884),
.Y(n_3262)
);

INVx6_ASAP7_75t_L g3263 ( 
.A(n_3069),
.Y(n_3263)
);

CKINVDCx11_ASAP7_75t_R g3264 ( 
.A(n_3012),
.Y(n_3264)
);

BUFx6f_ASAP7_75t_L g3265 ( 
.A(n_3143),
.Y(n_3265)
);

OAI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_3119),
.A2(n_2711),
.B1(n_2902),
.B2(n_2888),
.Y(n_3266)
);

INVx5_ASAP7_75t_L g3267 ( 
.A(n_3119),
.Y(n_3267)
);

INVx6_ASAP7_75t_L g3268 ( 
.A(n_3012),
.Y(n_3268)
);

INVx8_ASAP7_75t_L g3269 ( 
.A(n_2998),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2984),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2987),
.Y(n_3271)
);

BUFx6f_ASAP7_75t_L g3272 ( 
.A(n_3009),
.Y(n_3272)
);

INVx1_ASAP7_75t_SL g3273 ( 
.A(n_3136),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3061),
.A2(n_2926),
.B1(n_2977),
.B2(n_2884),
.Y(n_3274)
);

CKINVDCx20_ASAP7_75t_R g3275 ( 
.A(n_3138),
.Y(n_3275)
);

CKINVDCx11_ASAP7_75t_R g3276 ( 
.A(n_3036),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_SL g3277 ( 
.A1(n_3070),
.A2(n_2818),
.B1(n_2926),
.B2(n_2925),
.Y(n_3277)
);

BUFx10_ASAP7_75t_L g3278 ( 
.A(n_2996),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3060),
.Y(n_3279)
);

BUFx12f_ASAP7_75t_L g3280 ( 
.A(n_3023),
.Y(n_3280)
);

BUFx2_ASAP7_75t_L g3281 ( 
.A(n_3127),
.Y(n_3281)
);

INVx6_ASAP7_75t_L g3282 ( 
.A(n_3023),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2989),
.Y(n_3283)
);

CKINVDCx14_ASAP7_75t_R g3284 ( 
.A(n_3154),
.Y(n_3284)
);

INVx1_ASAP7_75t_SL g3285 ( 
.A(n_3031),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3102),
.B(n_2891),
.Y(n_3286)
);

INVx2_ASAP7_75t_SL g3287 ( 
.A(n_3146),
.Y(n_3287)
);

OAI22xp33_ASAP7_75t_L g3288 ( 
.A1(n_3116),
.A2(n_2902),
.B1(n_2888),
.B2(n_2868),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3072),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_2998),
.A2(n_2757),
.B1(n_2921),
.B2(n_2886),
.Y(n_3290)
);

NAND2x1p5_ASAP7_75t_L g3291 ( 
.A(n_2998),
.B(n_2641),
.Y(n_3291)
);

INVx6_ASAP7_75t_L g3292 ( 
.A(n_3041),
.Y(n_3292)
);

OAI21xp33_ASAP7_75t_L g3293 ( 
.A1(n_3122),
.A2(n_2890),
.B(n_2712),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3001),
.Y(n_3294)
);

INVx6_ASAP7_75t_L g3295 ( 
.A(n_3041),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_SL g3296 ( 
.A1(n_3041),
.A2(n_2936),
.B1(n_2980),
.B2(n_2680),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3063),
.Y(n_3297)
);

OAI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3162),
.A2(n_2757),
.B1(n_2886),
.B2(n_2880),
.Y(n_3298)
);

CKINVDCx20_ASAP7_75t_R g3299 ( 
.A(n_3092),
.Y(n_3299)
);

BUFx3_ASAP7_75t_L g3300 ( 
.A(n_3038),
.Y(n_3300)
);

NAND2x1p5_ASAP7_75t_L g3301 ( 
.A(n_3183),
.B(n_2840),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3008),
.A2(n_2837),
.B1(n_2970),
.B2(n_2969),
.Y(n_3302)
);

BUFx3_ASAP7_75t_L g3303 ( 
.A(n_3132),
.Y(n_3303)
);

INVx6_ASAP7_75t_L g3304 ( 
.A(n_3043),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3010),
.Y(n_3305)
);

INVx1_ASAP7_75t_SL g3306 ( 
.A(n_3182),
.Y(n_3306)
);

AOI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_3121),
.A2(n_2807),
.B1(n_2846),
.B2(n_2630),
.Y(n_3307)
);

BUFx8_ASAP7_75t_L g3308 ( 
.A(n_3047),
.Y(n_3308)
);

INVx1_ASAP7_75t_SL g3309 ( 
.A(n_3160),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3081),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3087),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_SL g3312 ( 
.A1(n_3065),
.A2(n_2678),
.B1(n_2671),
.B2(n_2688),
.Y(n_3312)
);

OAI22x1_ASAP7_75t_L g3313 ( 
.A1(n_3120),
.A2(n_2648),
.B1(n_2622),
.B2(n_2749),
.Y(n_3313)
);

BUFx2_ASAP7_75t_L g3314 ( 
.A(n_2988),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3100),
.Y(n_3315)
);

AOI22xp33_ASAP7_75t_L g3316 ( 
.A1(n_3017),
.A2(n_2726),
.B1(n_2953),
.B2(n_2646),
.Y(n_3316)
);

INVx6_ASAP7_75t_L g3317 ( 
.A(n_3256),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3010),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_3164),
.A2(n_2885),
.B1(n_2879),
.B2(n_2909),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_3227),
.A2(n_2883),
.B1(n_2727),
.B2(n_2769),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3230),
.A2(n_2742),
.B1(n_2788),
.B2(n_2774),
.Y(n_3321)
);

INVx4_ASAP7_75t_L g3322 ( 
.A(n_3025),
.Y(n_3322)
);

CKINVDCx5p33_ASAP7_75t_R g3323 ( 
.A(n_3220),
.Y(n_3323)
);

CKINVDCx11_ASAP7_75t_R g3324 ( 
.A(n_3120),
.Y(n_3324)
);

CKINVDCx11_ASAP7_75t_R g3325 ( 
.A(n_3007),
.Y(n_3325)
);

OAI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3074),
.A2(n_2748),
.B1(n_2674),
.B2(n_2797),
.Y(n_3326)
);

INVx4_ASAP7_75t_L g3327 ( 
.A(n_3025),
.Y(n_3327)
);

AOI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_3101),
.A2(n_2703),
.B1(n_2832),
.B2(n_2820),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3140),
.Y(n_3329)
);

NAND2x1p5_ASAP7_75t_L g3330 ( 
.A(n_3256),
.B(n_2889),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_SL g3331 ( 
.A1(n_3026),
.A2(n_2678),
.B1(n_2896),
.B2(n_2895),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_3237),
.A2(n_2806),
.B1(n_2803),
.B2(n_2935),
.Y(n_3332)
);

OAI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_2991),
.A2(n_2740),
.B1(n_2734),
.B2(n_2867),
.Y(n_3333)
);

CKINVDCx6p67_ASAP7_75t_R g3334 ( 
.A(n_3090),
.Y(n_3334)
);

OAI22xp5_ASAP7_75t_L g3335 ( 
.A1(n_3191),
.A2(n_2652),
.B1(n_2667),
.B2(n_2959),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3032),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_SL g3337 ( 
.A1(n_3133),
.A2(n_2854),
.B1(n_2930),
.B2(n_2873),
.Y(n_3337)
);

INVx8_ASAP7_75t_L g3338 ( 
.A(n_3025),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3156),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_SL g3340 ( 
.A1(n_3054),
.A2(n_2839),
.B1(n_2859),
.B2(n_2873),
.Y(n_3340)
);

OAI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_3209),
.A2(n_2954),
.B1(n_2947),
.B2(n_2747),
.Y(n_3341)
);

BUFx12f_ASAP7_75t_L g3342 ( 
.A(n_3030),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3103),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_3083),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3184),
.Y(n_3345)
);

CKINVDCx5p33_ASAP7_75t_R g3346 ( 
.A(n_3093),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3186),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3039),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3190),
.Y(n_3349)
);

BUFx2_ASAP7_75t_L g3350 ( 
.A(n_3254),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3202),
.A2(n_2871),
.B1(n_2914),
.B2(n_2927),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3192),
.Y(n_3352)
);

CKINVDCx20_ASAP7_75t_R g3353 ( 
.A(n_3049),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3194),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_SL g3355 ( 
.A1(n_3145),
.A2(n_2859),
.B1(n_2720),
.B2(n_2732),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3085),
.B(n_2794),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3002),
.A2(n_2923),
.B1(n_2952),
.B2(n_2946),
.Y(n_3357)
);

OAI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3086),
.A2(n_2810),
.B1(n_2759),
.B2(n_2893),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_SL g3359 ( 
.A1(n_3077),
.A2(n_2839),
.B1(n_2732),
.B2(n_2780),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3148),
.Y(n_3360)
);

OAI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_3107),
.A2(n_2912),
.B1(n_2900),
.B2(n_2780),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3150),
.Y(n_3362)
);

OAI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_3235),
.A2(n_2976),
.B1(n_2945),
.B2(n_2916),
.Y(n_3363)
);

CKINVDCx11_ASAP7_75t_R g3364 ( 
.A(n_3110),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3028),
.Y(n_3365)
);

BUFx3_ASAP7_75t_L g3366 ( 
.A(n_3016),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3257),
.A2(n_2762),
.B1(n_2665),
.B2(n_2945),
.Y(n_3367)
);

AOI21xp33_ASAP7_75t_L g3368 ( 
.A1(n_3113),
.A2(n_2916),
.B(n_2905),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3188),
.Y(n_3369)
);

INVx4_ASAP7_75t_L g3370 ( 
.A(n_3256),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3131),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3125),
.Y(n_3372)
);

AOI22xp33_ASAP7_75t_L g3373 ( 
.A1(n_3055),
.A2(n_2976),
.B1(n_2905),
.B2(n_2972),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3062),
.B(n_2707),
.Y(n_3374)
);

NAND2x1p5_ASAP7_75t_L g3375 ( 
.A(n_3247),
.B(n_2709),
.Y(n_3375)
);

OAI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_3193),
.A2(n_2670),
.B(n_2794),
.Y(n_3376)
);

BUFx3_ASAP7_75t_L g3377 ( 
.A(n_3091),
.Y(n_3377)
);

BUFx8_ASAP7_75t_L g3378 ( 
.A(n_3139),
.Y(n_3378)
);

INVx2_ASAP7_75t_SL g3379 ( 
.A(n_3000),
.Y(n_3379)
);

BUFx3_ASAP7_75t_L g3380 ( 
.A(n_2993),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_3125),
.Y(n_3381)
);

OAI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_3058),
.A2(n_3212),
.B1(n_3027),
.B2(n_3137),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3073),
.Y(n_3383)
);

BUFx3_ASAP7_75t_L g3384 ( 
.A(n_3165),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3142),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3158),
.B(n_2794),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3165),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3144),
.Y(n_3388)
);

NAND2x1p5_ASAP7_75t_L g3389 ( 
.A(n_3240),
.B(n_2709),
.Y(n_3389)
);

BUFx6f_ASAP7_75t_L g3390 ( 
.A(n_3009),
.Y(n_3390)
);

CKINVDCx11_ASAP7_75t_R g3391 ( 
.A(n_3009),
.Y(n_3391)
);

AOI22xp5_ASAP7_75t_SL g3392 ( 
.A1(n_3218),
.A2(n_2777),
.B1(n_2670),
.B2(n_2869),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3040),
.Y(n_3393)
);

OAI22xp5_ASAP7_75t_SL g3394 ( 
.A1(n_3223),
.A2(n_2777),
.B1(n_2670),
.B2(n_2869),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3078),
.A2(n_2972),
.B1(n_2904),
.B2(n_2869),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_3021),
.A2(n_2972),
.B1(n_2904),
.B2(n_2860),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_SL g3397 ( 
.A1(n_3177),
.A2(n_2904),
.B1(n_2860),
.B2(n_2709),
.Y(n_3397)
);

BUFx12f_ASAP7_75t_L g3398 ( 
.A(n_2990),
.Y(n_3398)
);

OAI22xp33_ASAP7_75t_L g3399 ( 
.A1(n_3098),
.A2(n_2860),
.B1(n_2777),
.B2(n_627),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_3051),
.Y(n_3400)
);

INVx6_ASAP7_75t_L g3401 ( 
.A(n_3240),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3175),
.Y(n_3402)
);

AOI22xp33_ASAP7_75t_SL g3403 ( 
.A1(n_3106),
.A2(n_624),
.B1(n_626),
.B2(n_629),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3216),
.Y(n_3404)
);

INVx1_ASAP7_75t_SL g3405 ( 
.A(n_3067),
.Y(n_3405)
);

HB1xp67_ASAP7_75t_SL g3406 ( 
.A(n_3168),
.Y(n_3406)
);

AOI22xp33_ASAP7_75t_L g3407 ( 
.A1(n_3176),
.A2(n_626),
.B1(n_629),
.B2(n_631),
.Y(n_3407)
);

OAI21xp5_ASAP7_75t_SL g3408 ( 
.A1(n_3157),
.A2(n_632),
.B(n_633),
.Y(n_3408)
);

CKINVDCx11_ASAP7_75t_R g3409 ( 
.A(n_3067),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3196),
.B(n_632),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_2999),
.Y(n_3411)
);

INVx6_ASAP7_75t_L g3412 ( 
.A(n_3046),
.Y(n_3412)
);

INVx1_ASAP7_75t_SL g3413 ( 
.A(n_3067),
.Y(n_3413)
);

BUFx4_ASAP7_75t_R g3414 ( 
.A(n_3111),
.Y(n_3414)
);

CKINVDCx5p33_ASAP7_75t_R g3415 ( 
.A(n_3088),
.Y(n_3415)
);

AOI22xp33_ASAP7_75t_L g3416 ( 
.A1(n_3210),
.A2(n_634),
.B1(n_636),
.B2(n_637),
.Y(n_3416)
);

BUFx2_ASAP7_75t_L g3417 ( 
.A(n_3108),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3053),
.Y(n_3418)
);

BUFx10_ASAP7_75t_L g3419 ( 
.A(n_3050),
.Y(n_3419)
);

AOI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3221),
.A2(n_634),
.B1(n_636),
.B2(n_637),
.Y(n_3420)
);

INVx3_ASAP7_75t_L g3421 ( 
.A(n_3108),
.Y(n_3421)
);

OR2x2_ASAP7_75t_L g3422 ( 
.A(n_3003),
.B(n_638),
.Y(n_3422)
);

INVx5_ASAP7_75t_L g3423 ( 
.A(n_3108),
.Y(n_3423)
);

BUFx2_ASAP7_75t_SL g3424 ( 
.A(n_3022),
.Y(n_3424)
);

BUFx12f_ASAP7_75t_L g3425 ( 
.A(n_3046),
.Y(n_3425)
);

OAI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_3115),
.A2(n_639),
.B1(n_640),
.B2(n_641),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3052),
.A2(n_639),
.B1(n_640),
.B2(n_643),
.Y(n_3427)
);

BUFx2_ASAP7_75t_SL g3428 ( 
.A(n_3224),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3174),
.A2(n_644),
.B1(n_645),
.B2(n_646),
.Y(n_3429)
);

OAI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3239),
.A2(n_646),
.B1(n_647),
.B2(n_648),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3229),
.Y(n_3431)
);

BUFx3_ASAP7_75t_L g3432 ( 
.A(n_3198),
.Y(n_3432)
);

CKINVDCx14_ASAP7_75t_R g3433 ( 
.A(n_3198),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3251),
.Y(n_3434)
);

AOI22xp5_ASAP7_75t_L g3435 ( 
.A1(n_3205),
.A2(n_647),
.B1(n_649),
.B2(n_650),
.Y(n_3435)
);

INVx6_ASAP7_75t_L g3436 ( 
.A(n_3198),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3242),
.A2(n_649),
.B1(n_651),
.B2(n_652),
.Y(n_3437)
);

CKINVDCx11_ASAP7_75t_R g3438 ( 
.A(n_3244),
.Y(n_3438)
);

BUFx2_ASAP7_75t_SL g3439 ( 
.A(n_3231),
.Y(n_3439)
);

BUFx3_ASAP7_75t_L g3440 ( 
.A(n_3187),
.Y(n_3440)
);

AOI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_3169),
.A2(n_651),
.B1(n_652),
.B2(n_653),
.Y(n_3441)
);

BUFx2_ASAP7_75t_L g3442 ( 
.A(n_3068),
.Y(n_3442)
);

CKINVDCx11_ASAP7_75t_R g3443 ( 
.A(n_3249),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2995),
.B(n_3149),
.Y(n_3444)
);

AOI22xp33_ASAP7_75t_L g3445 ( 
.A1(n_3170),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3251),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3251),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3179),
.B(n_654),
.Y(n_3448)
);

OAI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3204),
.A2(n_655),
.B1(n_656),
.B2(n_657),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3112),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3095),
.Y(n_3451)
);

CKINVDCx20_ASAP7_75t_R g3452 ( 
.A(n_3084),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_L g3453 ( 
.A1(n_3228),
.A2(n_657),
.B1(n_658),
.B2(n_659),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3241),
.A2(n_658),
.B1(n_659),
.B2(n_660),
.Y(n_3454)
);

BUFx2_ASAP7_75t_L g3455 ( 
.A(n_3068),
.Y(n_3455)
);

INVx6_ASAP7_75t_L g3456 ( 
.A(n_3024),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3173),
.Y(n_3457)
);

BUFx8_ASAP7_75t_SL g3458 ( 
.A(n_3124),
.Y(n_3458)
);

INVx6_ASAP7_75t_L g3459 ( 
.A(n_3172),
.Y(n_3459)
);

INVx6_ASAP7_75t_L g3460 ( 
.A(n_3135),
.Y(n_3460)
);

BUFx10_ASAP7_75t_L g3461 ( 
.A(n_3139),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2986),
.Y(n_3462)
);

BUFx2_ASAP7_75t_L g3463 ( 
.A(n_3068),
.Y(n_3463)
);

CKINVDCx11_ASAP7_75t_R g3464 ( 
.A(n_3139),
.Y(n_3464)
);

INVx4_ASAP7_75t_L g3465 ( 
.A(n_3245),
.Y(n_3465)
);

BUFx3_ASAP7_75t_L g3466 ( 
.A(n_3128),
.Y(n_3466)
);

INVx3_ASAP7_75t_L g3467 ( 
.A(n_3152),
.Y(n_3467)
);

NOR2xp33_ASAP7_75t_L g3468 ( 
.A(n_3234),
.B(n_660),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3064),
.A2(n_661),
.B1(n_662),
.B2(n_663),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3252),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_L g3471 ( 
.A1(n_3019),
.A2(n_661),
.B1(n_662),
.B2(n_663),
.Y(n_3471)
);

INVx2_ASAP7_75t_SL g3472 ( 
.A(n_3269),
.Y(n_3472)
);

INVx3_ASAP7_75t_L g3473 ( 
.A(n_3400),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3365),
.B(n_3013),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_3400),
.Y(n_3475)
);

INVx3_ASAP7_75t_L g3476 ( 
.A(n_3465),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3309),
.B(n_3181),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3303),
.B(n_3252),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3270),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3271),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3283),
.Y(n_3481)
);

AND2x4_ASAP7_75t_L g3482 ( 
.A(n_3348),
.B(n_3076),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3294),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_L g3484 ( 
.A(n_3460),
.B(n_3197),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3460),
.B(n_3153),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3297),
.Y(n_3486)
);

AOI21x1_ASAP7_75t_L g3487 ( 
.A1(n_3402),
.A2(n_2994),
.B(n_3203),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3310),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3305),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3311),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_3322),
.Y(n_3491)
);

HB1xp67_ASAP7_75t_L g3492 ( 
.A(n_3281),
.Y(n_3492)
);

CKINVDCx11_ASAP7_75t_R g3493 ( 
.A(n_3280),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3315),
.Y(n_3494)
);

OR2x2_ASAP7_75t_L g3495 ( 
.A(n_3366),
.B(n_3252),
.Y(n_3495)
);

INVx3_ASAP7_75t_L g3496 ( 
.A(n_3322),
.Y(n_3496)
);

INVx3_ASAP7_75t_L g3497 ( 
.A(n_3465),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3343),
.Y(n_3498)
);

OR2x6_ASAP7_75t_L g3499 ( 
.A(n_3338),
.B(n_3269),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3258),
.B(n_2992),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3462),
.B(n_3048),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3318),
.Y(n_3502)
);

BUFx4f_ASAP7_75t_SL g3503 ( 
.A(n_3342),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3336),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3369),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3360),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3371),
.B(n_2992),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3362),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3462),
.B(n_3226),
.Y(n_3509)
);

OR2x2_ASAP7_75t_L g3510 ( 
.A(n_3306),
.B(n_3099),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3318),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3385),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3411),
.Y(n_3513)
);

BUFx2_ASAP7_75t_L g3514 ( 
.A(n_3308),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3388),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3259),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3348),
.Y(n_3517)
);

OAI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3408),
.A2(n_3213),
.B(n_3180),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3393),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3350),
.B(n_3226),
.Y(n_3520)
);

INVx3_ASAP7_75t_L g3521 ( 
.A(n_3327),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3261),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3279),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3289),
.Y(n_3524)
);

OR2x2_ASAP7_75t_L g3525 ( 
.A(n_3285),
.B(n_3099),
.Y(n_3525)
);

HB1xp67_ASAP7_75t_L g3526 ( 
.A(n_3374),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3329),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3339),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3393),
.Y(n_3529)
);

BUFx2_ASAP7_75t_L g3530 ( 
.A(n_3308),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3418),
.Y(n_3531)
);

NAND2x1p5_ASAP7_75t_L g3532 ( 
.A(n_3267),
.B(n_3079),
.Y(n_3532)
);

AO31x2_ASAP7_75t_L g3533 ( 
.A1(n_3457),
.A2(n_3004),
.A3(n_3033),
.B(n_3035),
.Y(n_3533)
);

BUFx2_ASAP7_75t_L g3534 ( 
.A(n_3433),
.Y(n_3534)
);

OAI21x1_ASAP7_75t_L g3535 ( 
.A1(n_3467),
.A2(n_2983),
.B(n_3005),
.Y(n_3535)
);

CKINVDCx5p33_ASAP7_75t_R g3536 ( 
.A(n_3264),
.Y(n_3536)
);

HB1xp67_ASAP7_75t_L g3537 ( 
.A(n_3450),
.Y(n_3537)
);

INVx6_ASAP7_75t_L g3538 ( 
.A(n_3278),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3345),
.Y(n_3539)
);

INVx3_ASAP7_75t_L g3540 ( 
.A(n_3327),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3347),
.Y(n_3541)
);

BUFx6f_ASAP7_75t_L g3542 ( 
.A(n_3272),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3467),
.A2(n_3015),
.B(n_3018),
.Y(n_3543)
);

BUFx3_ASAP7_75t_L g3544 ( 
.A(n_3317),
.Y(n_3544)
);

BUFx2_ASAP7_75t_L g3545 ( 
.A(n_3425),
.Y(n_3545)
);

BUFx4f_ASAP7_75t_SL g3546 ( 
.A(n_3398),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3349),
.B(n_3226),
.Y(n_3547)
);

INVx2_ASAP7_75t_SL g3548 ( 
.A(n_3338),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3352),
.Y(n_3549)
);

CKINVDCx20_ASAP7_75t_R g3550 ( 
.A(n_3275),
.Y(n_3550)
);

BUFx2_ASAP7_75t_L g3551 ( 
.A(n_3314),
.Y(n_3551)
);

INVx11_ASAP7_75t_L g3552 ( 
.A(n_3282),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3354),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3356),
.Y(n_3554)
);

OAI21x1_ASAP7_75t_L g3555 ( 
.A1(n_3451),
.A2(n_3059),
.B(n_3075),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3431),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3386),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3434),
.Y(n_3558)
);

OR2x6_ASAP7_75t_L g3559 ( 
.A(n_3424),
.B(n_3096),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3446),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3447),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3422),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3372),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3381),
.Y(n_3564)
);

AOI22xp5_ASAP7_75t_L g3565 ( 
.A1(n_3266),
.A2(n_3123),
.B1(n_3215),
.B2(n_3243),
.Y(n_3565)
);

AOI22xp33_ASAP7_75t_L g3566 ( 
.A1(n_3334),
.A2(n_3089),
.B1(n_3080),
.B2(n_3161),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3387),
.B(n_3099),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3383),
.Y(n_3568)
);

INVx2_ASAP7_75t_SL g3569 ( 
.A(n_3412),
.Y(n_3569)
);

HB1xp67_ASAP7_75t_L g3570 ( 
.A(n_3470),
.Y(n_3570)
);

OAI21xp33_ASAP7_75t_SL g3571 ( 
.A1(n_3274),
.A2(n_3147),
.B(n_3246),
.Y(n_3571)
);

INVx3_ASAP7_75t_L g3572 ( 
.A(n_3370),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3461),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3442),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3455),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3461),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3404),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3463),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3272),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3410),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3444),
.Y(n_3581)
);

HB1xp67_ASAP7_75t_L g3582 ( 
.A(n_3417),
.Y(n_3582)
);

BUFx6f_ASAP7_75t_L g3583 ( 
.A(n_3272),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3384),
.B(n_3114),
.Y(n_3584)
);

INVx3_ASAP7_75t_L g3585 ( 
.A(n_3370),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3273),
.B(n_3114),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3364),
.Y(n_3587)
);

INVx3_ASAP7_75t_L g3588 ( 
.A(n_3440),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3390),
.Y(n_3589)
);

AND2x4_ASAP7_75t_L g3590 ( 
.A(n_3396),
.B(n_3421),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3286),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3448),
.Y(n_3592)
);

NAND2x1_ASAP7_75t_L g3593 ( 
.A(n_3401),
.B(n_3245),
.Y(n_3593)
);

BUFx3_ASAP7_75t_L g3594 ( 
.A(n_3317),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3379),
.Y(n_3595)
);

OR2x2_ASAP7_75t_L g3596 ( 
.A(n_3380),
.B(n_3114),
.Y(n_3596)
);

AND2x6_ASAP7_75t_L g3597 ( 
.A(n_3390),
.B(n_3159),
.Y(n_3597)
);

OAI21x1_ASAP7_75t_L g3598 ( 
.A1(n_3373),
.A2(n_3171),
.B(n_3056),
.Y(n_3598)
);

AO21x2_ASAP7_75t_L g3599 ( 
.A1(n_3376),
.A2(n_3117),
.B(n_3034),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3401),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3456),
.Y(n_3601)
);

INVx3_ASAP7_75t_L g3602 ( 
.A(n_3292),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3456),
.Y(n_3603)
);

HB1xp67_ASAP7_75t_L g3604 ( 
.A(n_3405),
.Y(n_3604)
);

OAI211xp5_ASAP7_75t_L g3605 ( 
.A1(n_3566),
.A2(n_3293),
.B(n_3324),
.C(n_3267),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_L g3606 ( 
.A(n_3587),
.B(n_3265),
.Y(n_3606)
);

OR2x6_ASAP7_75t_L g3607 ( 
.A(n_3499),
.B(n_3439),
.Y(n_3607)
);

NAND2xp33_ASAP7_75t_L g3608 ( 
.A(n_3536),
.B(n_3267),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3571),
.A2(n_3288),
.B(n_3333),
.Y(n_3609)
);

INVx3_ASAP7_75t_L g3610 ( 
.A(n_3572),
.Y(n_3610)
);

BUFx3_ASAP7_75t_L g3611 ( 
.A(n_3546),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3581),
.B(n_3298),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3492),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_3573),
.B(n_3265),
.Y(n_3614)
);

AND2x2_ASAP7_75t_L g3615 ( 
.A(n_3500),
.B(n_3419),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3551),
.B(n_3419),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3492),
.B(n_3526),
.Y(n_3617)
);

INVx4_ASAP7_75t_L g3618 ( 
.A(n_3499),
.Y(n_3618)
);

OAI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_3565),
.A2(n_3403),
.B(n_3290),
.Y(n_3619)
);

OAI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3566),
.A2(n_3214),
.B(n_3430),
.Y(n_3620)
);

INVx4_ASAP7_75t_L g3621 ( 
.A(n_3499),
.Y(n_3621)
);

OAI211xp5_ASAP7_75t_L g3622 ( 
.A1(n_3514),
.A2(n_3464),
.B(n_3277),
.C(n_3312),
.Y(n_3622)
);

AOI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_3591),
.A2(n_3406),
.B1(n_3326),
.B2(n_3382),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3526),
.B(n_3265),
.Y(n_3624)
);

AOI221xp5_ASAP7_75t_L g3625 ( 
.A1(n_3592),
.A2(n_3468),
.B1(n_3426),
.B2(n_3449),
.C(n_3399),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3554),
.B(n_3443),
.Y(n_3626)
);

OAI211xp5_ASAP7_75t_L g3627 ( 
.A1(n_3530),
.A2(n_3262),
.B(n_3325),
.C(n_3438),
.Y(n_3627)
);

OA21x2_ASAP7_75t_L g3628 ( 
.A1(n_3501),
.A2(n_3368),
.B(n_3302),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3498),
.Y(n_3629)
);

OR2x2_ASAP7_75t_L g3630 ( 
.A(n_3557),
.B(n_3287),
.Y(n_3630)
);

OAI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3538),
.A2(n_3337),
.B1(n_3296),
.B2(n_3359),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3582),
.B(n_3300),
.Y(n_3632)
);

OR2x2_ASAP7_75t_L g3633 ( 
.A(n_3477),
.B(n_3344),
.Y(n_3633)
);

OR2x2_ASAP7_75t_L g3634 ( 
.A(n_3513),
.B(n_3466),
.Y(n_3634)
);

A2O1A1Ixp33_ASAP7_75t_L g3635 ( 
.A1(n_3472),
.A2(n_3534),
.B(n_3548),
.C(n_3545),
.Y(n_3635)
);

AND2x4_ASAP7_75t_L g3636 ( 
.A(n_3573),
.B(n_3432),
.Y(n_3636)
);

INVx4_ASAP7_75t_L g3637 ( 
.A(n_3538),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3562),
.B(n_3378),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3582),
.B(n_3413),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3568),
.B(n_3378),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3507),
.B(n_3332),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3604),
.Y(n_3642)
);

A2O1A1Ixp33_ASAP7_75t_L g3643 ( 
.A1(n_3472),
.A2(n_3414),
.B(n_3377),
.C(n_3392),
.Y(n_3643)
);

NOR3xp33_ASAP7_75t_SL g3644 ( 
.A(n_3536),
.B(n_3323),
.C(n_3346),
.Y(n_3644)
);

NOR4xp25_ASAP7_75t_SL g3645 ( 
.A(n_3601),
.B(n_3415),
.C(n_3199),
.D(n_3200),
.Y(n_3645)
);

BUFx12f_ASAP7_75t_L g3646 ( 
.A(n_3493),
.Y(n_3646)
);

AO22x2_ASAP7_75t_L g3647 ( 
.A1(n_3576),
.A2(n_3428),
.B1(n_3341),
.B2(n_3363),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3604),
.B(n_3412),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3595),
.B(n_3421),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3479),
.Y(n_3650)
);

INVx4_ASAP7_75t_L g3651 ( 
.A(n_3538),
.Y(n_3651)
);

INVx4_ASAP7_75t_L g3652 ( 
.A(n_3572),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3480),
.B(n_3278),
.Y(n_3653)
);

AOI22xp5_ASAP7_75t_SL g3654 ( 
.A1(n_3548),
.A2(n_3299),
.B1(n_3284),
.B2(n_3291),
.Y(n_3654)
);

OAI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_3518),
.A2(n_3233),
.B(n_3420),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3546),
.A2(n_3331),
.B1(n_3355),
.B2(n_3367),
.Y(n_3656)
);

HB1xp67_ASAP7_75t_L g3657 ( 
.A(n_3506),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3481),
.B(n_3391),
.Y(n_3658)
);

OAI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3521),
.A2(n_3340),
.B1(n_3395),
.B2(n_3452),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3485),
.A2(n_3459),
.B1(n_3319),
.B2(n_3328),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3517),
.Y(n_3661)
);

NOR2xp33_ASAP7_75t_L g3662 ( 
.A(n_3552),
.B(n_3268),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3517),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3503),
.B(n_3268),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3519),
.Y(n_3665)
);

AOI21xp5_ASAP7_75t_SL g3666 ( 
.A1(n_3559),
.A2(n_3313),
.B(n_3389),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3483),
.B(n_3409),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3486),
.B(n_3304),
.Y(n_3668)
);

AND2x4_ASAP7_75t_L g3669 ( 
.A(n_3576),
.B(n_3423),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3513),
.B(n_3260),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_3473),
.B(n_3423),
.Y(n_3671)
);

OAI211xp5_ASAP7_75t_SL g3672 ( 
.A1(n_3484),
.A2(n_3307),
.B(n_3276),
.C(n_3441),
.Y(n_3672)
);

NOR2x1_ASAP7_75t_SL g3673 ( 
.A(n_3559),
.B(n_3423),
.Y(n_3673)
);

OAI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3474),
.A2(n_3037),
.B(n_3445),
.Y(n_3674)
);

NOR2x1_ASAP7_75t_SL g3675 ( 
.A(n_3559),
.B(n_3603),
.Y(n_3675)
);

OR2x6_ASAP7_75t_L g3676 ( 
.A(n_3521),
.B(n_3292),
.Y(n_3676)
);

A2O1A1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3585),
.A2(n_3163),
.B(n_3207),
.C(n_3155),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3531),
.B(n_3316),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3488),
.B(n_3304),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3657),
.Y(n_3680)
);

OR2x2_ASAP7_75t_L g3681 ( 
.A(n_3617),
.B(n_3574),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3661),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3663),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3665),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3607),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3629),
.Y(n_3686)
);

BUFx2_ASAP7_75t_L g3687 ( 
.A(n_3607),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3650),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3615),
.B(n_3586),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3641),
.B(n_3575),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3642),
.B(n_3578),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3652),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3613),
.B(n_3482),
.Y(n_3693)
);

BUFx2_ASAP7_75t_L g3694 ( 
.A(n_3607),
.Y(n_3694)
);

OR2x2_ASAP7_75t_L g3695 ( 
.A(n_3633),
.B(n_3510),
.Y(n_3695)
);

INVx2_ASAP7_75t_SL g3696 ( 
.A(n_3652),
.Y(n_3696)
);

AND2x2_ASAP7_75t_SL g3697 ( 
.A(n_3618),
.B(n_3478),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3678),
.B(n_3509),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3630),
.Y(n_3699)
);

OR2x2_ASAP7_75t_L g3700 ( 
.A(n_3634),
.B(n_3525),
.Y(n_3700)
);

AND2x4_ASAP7_75t_L g3701 ( 
.A(n_3675),
.B(n_3476),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3624),
.B(n_3482),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3610),
.Y(n_3703)
);

AOI22xp33_ASAP7_75t_L g3704 ( 
.A1(n_3619),
.A2(n_3459),
.B1(n_3484),
.B2(n_3485),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3653),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3639),
.B(n_3482),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3614),
.B(n_3584),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3610),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3612),
.Y(n_3709)
);

AOI22xp33_ASAP7_75t_L g3710 ( 
.A1(n_3619),
.A2(n_3394),
.B1(n_3597),
.B2(n_3600),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3640),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3660),
.B(n_3520),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3649),
.Y(n_3713)
);

AOI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3631),
.A2(n_3597),
.B1(n_3596),
.B2(n_3580),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3636),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3614),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3648),
.B(n_3567),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3668),
.Y(n_3718)
);

INVxp67_ASAP7_75t_L g3719 ( 
.A(n_3632),
.Y(n_3719)
);

INVxp67_ASAP7_75t_SL g3720 ( 
.A(n_3673),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3636),
.B(n_3476),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3669),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3669),
.Y(n_3723)
);

AND2x4_ASAP7_75t_L g3724 ( 
.A(n_3618),
.B(n_3476),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3660),
.B(n_3531),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3638),
.B(n_3497),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3679),
.B(n_3497),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3670),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3647),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3647),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3609),
.B(n_3508),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3628),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3628),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3671),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3671),
.Y(n_3735)
);

OR2x2_ASAP7_75t_L g3736 ( 
.A(n_3616),
.B(n_3495),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_3701),
.Y(n_3737)
);

BUFx2_ASAP7_75t_L g3738 ( 
.A(n_3720),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3689),
.B(n_3626),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3689),
.B(n_3497),
.Y(n_3740)
);

AND2x4_ASAP7_75t_L g3741 ( 
.A(n_3685),
.B(n_3621),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3682),
.Y(n_3742)
);

AND2x4_ASAP7_75t_L g3743 ( 
.A(n_3685),
.B(n_3621),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_L g3744 ( 
.A1(n_3710),
.A2(n_3656),
.B1(n_3672),
.B2(n_3659),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3711),
.B(n_3658),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3709),
.B(n_3490),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3684),
.Y(n_3747)
);

AOI22xp33_ASAP7_75t_L g3748 ( 
.A1(n_3714),
.A2(n_3620),
.B1(n_3623),
.B2(n_3655),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3711),
.B(n_3667),
.Y(n_3749)
);

OAI221xp5_ASAP7_75t_L g3750 ( 
.A1(n_3704),
.A2(n_3623),
.B1(n_3605),
.B2(n_3622),
.C(n_3635),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_SL g3751 ( 
.A1(n_3687),
.A2(n_3654),
.B1(n_3637),
.B2(n_3651),
.Y(n_3751)
);

INVxp67_ASAP7_75t_SL g3752 ( 
.A(n_3696),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3682),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3684),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3683),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3687),
.A2(n_3620),
.B1(n_3655),
.B2(n_3625),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3693),
.B(n_3570),
.Y(n_3757)
);

AOI221xp5_ASAP7_75t_L g3758 ( 
.A1(n_3709),
.A2(n_3674),
.B1(n_3666),
.B2(n_3627),
.C(n_3643),
.Y(n_3758)
);

OAI22xp5_ASAP7_75t_L g3759 ( 
.A1(n_3694),
.A2(n_3696),
.B1(n_3654),
.B2(n_3731),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3712),
.B(n_3494),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3701),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3693),
.B(n_3570),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3683),
.Y(n_3763)
);

NAND2xp33_ASAP7_75t_R g3764 ( 
.A(n_3694),
.B(n_3644),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3728),
.B(n_3537),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3725),
.B(n_3504),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3701),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3686),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3686),
.Y(n_3769)
);

AO21x2_ASAP7_75t_L g3770 ( 
.A1(n_3732),
.A2(n_3487),
.B(n_3674),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3688),
.Y(n_3771)
);

AND2x4_ASAP7_75t_L g3772 ( 
.A(n_3729),
.B(n_3588),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3691),
.B(n_3505),
.Y(n_3773)
);

AOI221xp5_ASAP7_75t_L g3774 ( 
.A1(n_3729),
.A2(n_3608),
.B1(n_3512),
.B2(n_3515),
.C(n_3606),
.Y(n_3774)
);

OA21x2_ASAP7_75t_L g3775 ( 
.A1(n_3730),
.A2(n_3535),
.B(n_3543),
.Y(n_3775)
);

HB1xp67_ASAP7_75t_L g3776 ( 
.A(n_3680),
.Y(n_3776)
);

HB1xp67_ASAP7_75t_L g3777 ( 
.A(n_3680),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3688),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3700),
.Y(n_3779)
);

AND4x1_ASAP7_75t_L g3780 ( 
.A(n_3730),
.B(n_3664),
.C(n_3662),
.D(n_3646),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3691),
.B(n_3519),
.Y(n_3781)
);

AO221x2_ASAP7_75t_L g3782 ( 
.A1(n_3692),
.A2(n_3503),
.B1(n_3493),
.B2(n_3611),
.C(n_3282),
.Y(n_3782)
);

AO21x2_ASAP7_75t_L g3783 ( 
.A1(n_3732),
.A2(n_3555),
.B(n_3677),
.Y(n_3783)
);

OR2x2_ASAP7_75t_L g3784 ( 
.A(n_3681),
.B(n_3533),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3719),
.B(n_3637),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3700),
.Y(n_3786)
);

AND2x4_ASAP7_75t_L g3787 ( 
.A(n_3724),
.B(n_3588),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3690),
.B(n_3529),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3681),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3728),
.B(n_3537),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3738),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3738),
.B(n_3740),
.Y(n_3792)
);

HB1xp67_ASAP7_75t_L g3793 ( 
.A(n_3752),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3776),
.Y(n_3794)
);

AND2x4_ASAP7_75t_L g3795 ( 
.A(n_3741),
.B(n_3733),
.Y(n_3795)
);

OR2x2_ASAP7_75t_L g3796 ( 
.A(n_3784),
.B(n_3733),
.Y(n_3796)
);

OR2x6_ASAP7_75t_L g3797 ( 
.A(n_3759),
.B(n_3651),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3740),
.B(n_3706),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3777),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3779),
.B(n_3706),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3779),
.B(n_3718),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3769),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3786),
.B(n_3718),
.Y(n_3803)
);

OR2x2_ASAP7_75t_L g3804 ( 
.A(n_3784),
.B(n_3695),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3769),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3786),
.B(n_3702),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3757),
.B(n_3702),
.Y(n_3807)
);

OR2x6_ASAP7_75t_L g3808 ( 
.A(n_3759),
.B(n_3676),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3757),
.B(n_3699),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3765),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3765),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3762),
.B(n_3699),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3756),
.B(n_3698),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3790),
.Y(n_3814)
);

BUFx2_ASAP7_75t_L g3815 ( 
.A(n_3737),
.Y(n_3815)
);

AND2x2_ASAP7_75t_SL g3816 ( 
.A(n_3780),
.B(n_3697),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3762),
.B(n_3717),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3770),
.B(n_3789),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_L g3819 ( 
.A(n_3780),
.B(n_3705),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3790),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3782),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3770),
.B(n_3713),
.Y(n_3822)
);

HB1xp67_ASAP7_75t_L g3823 ( 
.A(n_3782),
.Y(n_3823)
);

AND2x4_ASAP7_75t_L g3824 ( 
.A(n_3741),
.B(n_3724),
.Y(n_3824)
);

NOR2x1_ASAP7_75t_SL g3825 ( 
.A(n_3782),
.B(n_3676),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3797),
.B(n_3772),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3797),
.B(n_3772),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3793),
.Y(n_3828)
);

INVxp67_ASAP7_75t_L g3829 ( 
.A(n_3821),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3797),
.B(n_3772),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_L g3831 ( 
.A(n_3823),
.B(n_3750),
.Y(n_3831)
);

NOR3xp33_ASAP7_75t_L g3832 ( 
.A(n_3791),
.B(n_3758),
.C(n_3751),
.Y(n_3832)
);

OAI21xp33_ASAP7_75t_L g3833 ( 
.A1(n_3808),
.A2(n_3744),
.B(n_3748),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3825),
.B(n_3741),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3792),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3792),
.Y(n_3836)
);

HB1xp67_ASAP7_75t_L g3837 ( 
.A(n_3794),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3809),
.Y(n_3838)
);

OR2x2_ASAP7_75t_L g3839 ( 
.A(n_3804),
.B(n_3760),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3809),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3804),
.Y(n_3841)
);

NOR2xp67_ASAP7_75t_L g3842 ( 
.A(n_3824),
.B(n_3737),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3812),
.Y(n_3843)
);

AND2x4_ASAP7_75t_SL g3844 ( 
.A(n_3797),
.B(n_3782),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3813),
.B(n_3770),
.Y(n_3845)
);

NOR2xp67_ASAP7_75t_L g3846 ( 
.A(n_3824),
.B(n_3737),
.Y(n_3846)
);

NAND3xp33_ASAP7_75t_L g3847 ( 
.A(n_3808),
.B(n_3818),
.C(n_3822),
.Y(n_3847)
);

INVx1_ASAP7_75t_SL g3848 ( 
.A(n_3816),
.Y(n_3848)
);

OR2x2_ASAP7_75t_L g3849 ( 
.A(n_3796),
.B(n_3766),
.Y(n_3849)
);

AND2x4_ASAP7_75t_SL g3850 ( 
.A(n_3808),
.B(n_3741),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3812),
.Y(n_3851)
);

INVx2_ASAP7_75t_SL g3852 ( 
.A(n_3816),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3799),
.B(n_3774),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3796),
.Y(n_3854)
);

OR2x2_ASAP7_75t_L g3855 ( 
.A(n_3808),
.B(n_3789),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3795),
.B(n_3817),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3810),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3795),
.B(n_3817),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3828),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3854),
.Y(n_3860)
);

OR2x2_ASAP7_75t_L g3861 ( 
.A(n_3841),
.B(n_3811),
.Y(n_3861)
);

NAND2xp33_ASAP7_75t_SL g3862 ( 
.A(n_3834),
.B(n_3764),
.Y(n_3862)
);

INVx4_ASAP7_75t_L g3863 ( 
.A(n_3844),
.Y(n_3863)
);

OAI31xp33_ASAP7_75t_L g3864 ( 
.A1(n_3833),
.A2(n_3815),
.A3(n_3819),
.B(n_3795),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3831),
.B(n_3814),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3837),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3841),
.Y(n_3867)
);

OR2x2_ASAP7_75t_L g3868 ( 
.A(n_3849),
.B(n_3820),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3835),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3831),
.B(n_3783),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3849),
.B(n_3839),
.Y(n_3871)
);

INVxp67_ASAP7_75t_L g3872 ( 
.A(n_3845),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_3834),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3854),
.Y(n_3874)
);

NAND2x1p5_ASAP7_75t_L g3875 ( 
.A(n_3834),
.B(n_3743),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3835),
.Y(n_3876)
);

INVxp67_ASAP7_75t_L g3877 ( 
.A(n_3853),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3836),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3829),
.B(n_3783),
.Y(n_3879)
);

OR2x2_ASAP7_75t_L g3880 ( 
.A(n_3839),
.B(n_3788),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3836),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3838),
.Y(n_3882)
);

OAI21xp33_ASAP7_75t_L g3883 ( 
.A1(n_3848),
.A2(n_3743),
.B(n_3824),
.Y(n_3883)
);

A2O1A1O1Ixp25_ASAP7_75t_L g3884 ( 
.A1(n_3883),
.A2(n_3852),
.B(n_3844),
.C(n_3850),
.D(n_3847),
.Y(n_3884)
);

OAI21xp33_ASAP7_75t_L g3885 ( 
.A1(n_3877),
.A2(n_3852),
.B(n_3832),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3871),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3873),
.B(n_3850),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3863),
.B(n_3855),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3867),
.Y(n_3889)
);

OR2x2_ASAP7_75t_L g3890 ( 
.A(n_3865),
.B(n_3840),
.Y(n_3890)
);

AND2x4_ASAP7_75t_L g3891 ( 
.A(n_3863),
.B(n_3825),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3877),
.B(n_3843),
.Y(n_3892)
);

OAI221xp5_ASAP7_75t_L g3893 ( 
.A1(n_3864),
.A2(n_3846),
.B1(n_3842),
.B2(n_3815),
.C(n_3826),
.Y(n_3893)
);

NAND4xp75_ASAP7_75t_L g3894 ( 
.A(n_3870),
.B(n_3827),
.C(n_3830),
.D(n_3826),
.Y(n_3894)
);

AOI221xp5_ASAP7_75t_L g3895 ( 
.A1(n_3862),
.A2(n_3866),
.B1(n_3872),
.B2(n_3859),
.C(n_3879),
.Y(n_3895)
);

OAI32xp33_ASAP7_75t_L g3896 ( 
.A1(n_3862),
.A2(n_3827),
.A3(n_3830),
.B1(n_3858),
.B2(n_3856),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3860),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3872),
.A2(n_3858),
.B(n_3856),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3860),
.Y(n_3899)
);

OAI22xp5_ASAP7_75t_L g3900 ( 
.A1(n_3875),
.A2(n_3851),
.B1(n_3743),
.B2(n_3857),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3874),
.Y(n_3901)
);

INVxp67_ASAP7_75t_L g3902 ( 
.A(n_3874),
.Y(n_3902)
);

AOI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_3882),
.A2(n_3743),
.B1(n_3353),
.B2(n_3783),
.Y(n_3903)
);

AOI21xp33_ASAP7_75t_L g3904 ( 
.A1(n_3878),
.A2(n_3775),
.B(n_3772),
.Y(n_3904)
);

AOI222xp33_ASAP7_75t_L g3905 ( 
.A1(n_3885),
.A2(n_3869),
.B1(n_3876),
.B2(n_3881),
.C1(n_3878),
.C2(n_3550),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3898),
.B(n_3881),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3887),
.B(n_3875),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3886),
.B(n_3880),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3889),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3891),
.A2(n_3868),
.B1(n_3861),
.B2(n_3785),
.Y(n_3910)
);

CKINVDCx14_ASAP7_75t_R g3911 ( 
.A(n_3888),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3897),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3899),
.Y(n_3913)
);

AOI322xp5_ASAP7_75t_L g3914 ( 
.A1(n_3891),
.A2(n_3745),
.A3(n_3749),
.B1(n_3739),
.B2(n_3803),
.C1(n_3801),
.C2(n_3800),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3896),
.B(n_3550),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3901),
.Y(n_3916)
);

OAI22xp33_ASAP7_75t_L g3917 ( 
.A1(n_3884),
.A2(n_3767),
.B1(n_3761),
.B2(n_3692),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3895),
.A2(n_3749),
.B(n_3745),
.Y(n_3918)
);

AOI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3893),
.A2(n_3746),
.B(n_3739),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3902),
.Y(n_3920)
);

NAND4xp25_ASAP7_75t_L g3921 ( 
.A(n_3892),
.B(n_3416),
.C(n_3407),
.D(n_3453),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3890),
.Y(n_3922)
);

OAI21xp33_ASAP7_75t_L g3923 ( 
.A1(n_3900),
.A2(n_3767),
.B(n_3761),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3904),
.A2(n_3805),
.B(n_3802),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3894),
.Y(n_3925)
);

OAI21xp33_ASAP7_75t_L g3926 ( 
.A1(n_3903),
.A2(n_3773),
.B(n_3801),
.Y(n_3926)
);

AOI211x1_ASAP7_75t_L g3927 ( 
.A1(n_3903),
.A2(n_3803),
.B(n_3798),
.C(n_3807),
.Y(n_3927)
);

OAI21xp5_ASAP7_75t_SL g3928 ( 
.A1(n_3911),
.A2(n_3435),
.B(n_3454),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3906),
.Y(n_3929)
);

OR2x2_ASAP7_75t_L g3930 ( 
.A(n_3908),
.B(n_3806),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3909),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3907),
.B(n_3798),
.Y(n_3932)
);

BUFx3_ASAP7_75t_L g3933 ( 
.A(n_3920),
.Y(n_3933)
);

OAI221xp5_ASAP7_75t_L g3934 ( 
.A1(n_3915),
.A2(n_3263),
.B1(n_3532),
.B2(n_3397),
.C(n_3544),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3905),
.B(n_3802),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3922),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3912),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3913),
.B(n_3805),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3925),
.A2(n_3645),
.B(n_3807),
.Y(n_3939)
);

OAI222xp33_ASAP7_75t_L g3940 ( 
.A1(n_3916),
.A2(n_3532),
.B1(n_3676),
.B2(n_3736),
.C1(n_3735),
.C2(n_3734),
.Y(n_3940)
);

OAI22xp33_ASAP7_75t_SL g3941 ( 
.A1(n_3910),
.A2(n_3263),
.B1(n_3295),
.B2(n_3544),
.Y(n_3941)
);

OAI21xp33_ASAP7_75t_L g3942 ( 
.A1(n_3905),
.A2(n_3726),
.B(n_3594),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3914),
.B(n_3806),
.Y(n_3943)
);

NAND4xp25_ASAP7_75t_SL g3944 ( 
.A(n_3918),
.B(n_3800),
.C(n_3736),
.D(n_3734),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3917),
.A2(n_3923),
.B1(n_3919),
.B2(n_3926),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3924),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3927),
.B(n_3771),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3921),
.Y(n_3948)
);

AOI322xp5_ASAP7_75t_L g3949 ( 
.A1(n_3921),
.A2(n_3726),
.A3(n_3713),
.B1(n_3735),
.B2(n_3697),
.C1(n_3781),
.C2(n_3787),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3906),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3933),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3931),
.Y(n_3952)
);

NAND2xp33_ASAP7_75t_SL g3953 ( 
.A(n_3948),
.B(n_3645),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3932),
.B(n_3771),
.Y(n_3954)
);

AOI211xp5_ASAP7_75t_SL g3955 ( 
.A1(n_3929),
.A2(n_3201),
.B(n_3189),
.C(n_3208),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3936),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3950),
.Y(n_3957)
);

O2A1O1Ixp33_ASAP7_75t_L g3958 ( 
.A1(n_3937),
.A2(n_3219),
.B(n_3222),
.C(n_3217),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3946),
.B(n_3778),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3941),
.B(n_3787),
.Y(n_3960)
);

NAND3xp33_ASAP7_75t_L g3961 ( 
.A(n_3945),
.B(n_3427),
.C(n_3236),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3930),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3938),
.Y(n_3963)
);

OAI211xp5_ASAP7_75t_L g3964 ( 
.A1(n_3928),
.A2(n_3429),
.B(n_3437),
.C(n_3471),
.Y(n_3964)
);

AND2x4_ASAP7_75t_L g3965 ( 
.A(n_3943),
.B(n_3787),
.Y(n_3965)
);

OAI211xp5_ASAP7_75t_L g3966 ( 
.A1(n_3928),
.A2(n_3939),
.B(n_3935),
.C(n_3942),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3938),
.Y(n_3967)
);

NOR2xp67_ASAP7_75t_L g3968 ( 
.A(n_3934),
.B(n_664),
.Y(n_3968)
);

AND2x4_ASAP7_75t_L g3969 ( 
.A(n_3947),
.B(n_3787),
.Y(n_3969)
);

NAND4xp25_ASAP7_75t_L g3970 ( 
.A(n_3949),
.B(n_3211),
.C(n_3238),
.D(n_3225),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3947),
.Y(n_3971)
);

BUFx2_ASAP7_75t_L g3972 ( 
.A(n_3940),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_SL g3973 ( 
.A(n_3944),
.B(n_3724),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3946),
.A2(n_3130),
.B(n_3129),
.Y(n_3974)
);

NOR2x1_ASAP7_75t_L g3975 ( 
.A(n_3933),
.B(n_3134),
.Y(n_3975)
);

INVx2_ASAP7_75t_SL g3976 ( 
.A(n_3933),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3948),
.B(n_3778),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3929),
.B(n_3458),
.Y(n_3978)
);

OAI22xp33_ASAP7_75t_L g3979 ( 
.A1(n_3948),
.A2(n_3594),
.B1(n_3295),
.B2(n_3496),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3948),
.B(n_3602),
.Y(n_3980)
);

OAI211xp5_ASAP7_75t_L g3981 ( 
.A1(n_3951),
.A2(n_3167),
.B(n_3185),
.C(n_3178),
.Y(n_3981)
);

OAI221xp5_ASAP7_75t_L g3982 ( 
.A1(n_3953),
.A2(n_3469),
.B1(n_3320),
.B2(n_3141),
.C(n_3321),
.Y(n_3982)
);

AOI221xp5_ASAP7_75t_L g3983 ( 
.A1(n_3976),
.A2(n_3361),
.B1(n_3250),
.B2(n_3206),
.C(n_3358),
.Y(n_3983)
);

AOI31xp33_ASAP7_75t_L g3984 ( 
.A1(n_3957),
.A2(n_3097),
.A3(n_3330),
.B(n_3118),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_L g3985 ( 
.A1(n_3972),
.A2(n_3775),
.B1(n_3602),
.B2(n_3585),
.Y(n_3985)
);

OAI222xp33_ASAP7_75t_L g3986 ( 
.A1(n_3956),
.A2(n_3301),
.B1(n_3496),
.B2(n_3491),
.C1(n_3540),
.C2(n_3521),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3978),
.A2(n_3491),
.B1(n_3716),
.B2(n_3569),
.Y(n_3987)
);

NAND4xp25_ASAP7_75t_L g3988 ( 
.A(n_3968),
.B(n_3248),
.C(n_3255),
.D(n_3253),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3965),
.A2(n_3775),
.B1(n_3569),
.B2(n_3716),
.Y(n_3989)
);

NOR3xp33_ASAP7_75t_L g3990 ( 
.A(n_3966),
.B(n_3071),
.C(n_3166),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_L g3991 ( 
.A(n_3952),
.B(n_3962),
.Y(n_3991)
);

NAND3xp33_ASAP7_75t_L g3992 ( 
.A(n_3963),
.B(n_3151),
.C(n_3104),
.Y(n_3992)
);

AO221x1_ASAP7_75t_L g3993 ( 
.A1(n_3979),
.A2(n_3540),
.B1(n_3335),
.B2(n_3475),
.C(n_3473),
.Y(n_3993)
);

AOI322xp5_ASAP7_75t_L g3994 ( 
.A1(n_3967),
.A2(n_3697),
.A3(n_3727),
.B1(n_3593),
.B2(n_3703),
.C1(n_3708),
.C2(n_3763),
.Y(n_3994)
);

AOI221xp5_ASAP7_75t_L g3995 ( 
.A1(n_3980),
.A2(n_2985),
.B1(n_3763),
.B2(n_3755),
.C(n_3753),
.Y(n_3995)
);

OAI321xp33_ASAP7_75t_L g3996 ( 
.A1(n_3971),
.A2(n_3703),
.A3(n_3708),
.B1(n_3695),
.B2(n_3753),
.C(n_3755),
.Y(n_3996)
);

OAI322xp33_ASAP7_75t_L g3997 ( 
.A1(n_3959),
.A2(n_3742),
.A3(n_3768),
.B1(n_3754),
.B2(n_3747),
.C1(n_3722),
.C2(n_3723),
.Y(n_3997)
);

NOR4xp75_ASAP7_75t_L g3998 ( 
.A(n_3977),
.B(n_3540),
.C(n_3727),
.D(n_3721),
.Y(n_3998)
);

A2O1A1Ixp33_ASAP7_75t_L g3999 ( 
.A1(n_3961),
.A2(n_2997),
.B(n_3011),
.C(n_3020),
.Y(n_3999)
);

NOR4xp25_ASAP7_75t_L g4000 ( 
.A(n_3973),
.B(n_3742),
.C(n_3042),
.D(n_3768),
.Y(n_4000)
);

AOI211xp5_ASAP7_75t_SL g4001 ( 
.A1(n_3964),
.A2(n_3721),
.B(n_666),
.C(n_664),
.Y(n_4001)
);

AOI32xp33_ASAP7_75t_L g4002 ( 
.A1(n_3975),
.A2(n_3590),
.A3(n_3723),
.B1(n_3722),
.B2(n_3126),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3965),
.B(n_3969),
.Y(n_4003)
);

A2O1A1Ixp33_ASAP7_75t_SL g4004 ( 
.A1(n_3974),
.A2(n_667),
.B(n_665),
.C(n_666),
.Y(n_4004)
);

AOI221xp5_ASAP7_75t_L g4005 ( 
.A1(n_3970),
.A2(n_3351),
.B1(n_3747),
.B2(n_3754),
.C(n_3057),
.Y(n_4005)
);

HB1xp67_ASAP7_75t_L g4006 ( 
.A(n_3991),
.Y(n_4006)
);

OAI211xp5_ASAP7_75t_SL g4007 ( 
.A1(n_4001),
.A2(n_3960),
.B(n_3954),
.C(n_3955),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_4003),
.Y(n_4008)
);

AND4x1_ASAP7_75t_L g4009 ( 
.A(n_3985),
.B(n_3958),
.C(n_3969),
.D(n_669),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3989),
.A2(n_3715),
.B1(n_3775),
.B2(n_3475),
.Y(n_4010)
);

AOI322xp5_ASAP7_75t_L g4011 ( 
.A1(n_3990),
.A2(n_3715),
.A3(n_3707),
.B1(n_3590),
.B2(n_3717),
.C1(n_3357),
.C2(n_3473),
.Y(n_4011)
);

NAND3xp33_ASAP7_75t_SL g4012 ( 
.A(n_4004),
.B(n_667),
.C(n_668),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3984),
.Y(n_4013)
);

AOI22xp5_ASAP7_75t_L g4014 ( 
.A1(n_3993),
.A2(n_3597),
.B1(n_3707),
.B2(n_3590),
.Y(n_4014)
);

AOI211xp5_ASAP7_75t_L g4015 ( 
.A1(n_4000),
.A2(n_3232),
.B(n_3195),
.C(n_3109),
.Y(n_4015)
);

NOR3xp33_ASAP7_75t_L g4016 ( 
.A(n_3988),
.B(n_668),
.C(n_669),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_4005),
.Y(n_4017)
);

NAND4xp25_ASAP7_75t_L g4018 ( 
.A(n_3995),
.B(n_670),
.C(n_671),
.D(n_673),
.Y(n_4018)
);

AOI211xp5_ASAP7_75t_L g4019 ( 
.A1(n_3986),
.A2(n_670),
.B(n_674),
.C(n_675),
.Y(n_4019)
);

NAND3xp33_ASAP7_75t_L g4020 ( 
.A(n_4002),
.B(n_674),
.C(n_676),
.Y(n_4020)
);

NAND3xp33_ASAP7_75t_L g4021 ( 
.A(n_3981),
.B(n_676),
.C(n_677),
.Y(n_4021)
);

OAI221xp5_ASAP7_75t_L g4022 ( 
.A1(n_3982),
.A2(n_3436),
.B1(n_3375),
.B2(n_3475),
.C(n_3045),
.Y(n_4022)
);

BUFx6f_ASAP7_75t_L g4023 ( 
.A(n_3992),
.Y(n_4023)
);

OAI211xp5_ASAP7_75t_SL g4024 ( 
.A1(n_3994),
.A2(n_677),
.B(n_678),
.C(n_679),
.Y(n_4024)
);

AOI211xp5_ASAP7_75t_L g4025 ( 
.A1(n_3987),
.A2(n_679),
.B(n_680),
.C(n_681),
.Y(n_4025)
);

AOI221xp5_ASAP7_75t_L g4026 ( 
.A1(n_3996),
.A2(n_3066),
.B1(n_3588),
.B2(n_3563),
.C(n_3564),
.Y(n_4026)
);

AOI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3983),
.A2(n_3597),
.B1(n_3599),
.B2(n_3436),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3997),
.Y(n_4028)
);

XNOR2xp5_ASAP7_75t_L g4029 ( 
.A(n_4019),
.B(n_3998),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_4006),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_4008),
.Y(n_4031)
);

BUFx2_ASAP7_75t_L g4032 ( 
.A(n_4013),
.Y(n_4032)
);

INVx1_ASAP7_75t_SL g4033 ( 
.A(n_4017),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_4023),
.Y(n_4034)
);

NOR2x1_ASAP7_75t_L g4035 ( 
.A(n_4012),
.B(n_3999),
.Y(n_4035)
);

NOR2x1_ASAP7_75t_L g4036 ( 
.A(n_4018),
.B(n_680),
.Y(n_4036)
);

NAND4xp75_ASAP7_75t_L g4037 ( 
.A(n_4028),
.B(n_681),
.C(n_682),
.D(n_683),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_4021),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_4025),
.B(n_682),
.Y(n_4039)
);

AND4x1_ASAP7_75t_L g4040 ( 
.A(n_4016),
.B(n_685),
.C(n_687),
.D(n_688),
.Y(n_4040)
);

OR2x2_ASAP7_75t_L g4041 ( 
.A(n_4020),
.B(n_685),
.Y(n_4041)
);

INVxp33_ASAP7_75t_L g4042 ( 
.A(n_4022),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_4009),
.Y(n_4043)
);

AOI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_4007),
.A2(n_3597),
.B1(n_3599),
.B2(n_3542),
.Y(n_4044)
);

NOR4xp75_ASAP7_75t_L g4045 ( 
.A(n_4010),
.B(n_687),
.C(n_689),
.D(n_690),
.Y(n_4045)
);

AND2x4_ASAP7_75t_L g4046 ( 
.A(n_4014),
.B(n_3579),
.Y(n_4046)
);

INVxp67_ASAP7_75t_L g4047 ( 
.A(n_4023),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_4024),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_4027),
.Y(n_4049)
);

OAI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_4026),
.A2(n_3589),
.B1(n_3579),
.B2(n_3583),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_4015),
.Y(n_4051)
);

XNOR2xp5_ASAP7_75t_L g4052 ( 
.A(n_4040),
.B(n_4011),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_4037),
.B(n_4030),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_4033),
.B(n_4031),
.Y(n_4054)
);

OAI211xp5_ASAP7_75t_L g4055 ( 
.A1(n_4036),
.A2(n_691),
.B(n_692),
.C(n_693),
.Y(n_4055)
);

NAND4xp25_ASAP7_75t_L g4056 ( 
.A(n_4035),
.B(n_691),
.C(n_692),
.D(n_693),
.Y(n_4056)
);

AOI221x1_ASAP7_75t_L g4057 ( 
.A1(n_4034),
.A2(n_694),
.B1(n_695),
.B2(n_696),
.C(n_697),
.Y(n_4057)
);

A2O1A1O1Ixp25_ASAP7_75t_L g4058 ( 
.A1(n_4048),
.A2(n_3044),
.B(n_3549),
.C(n_3541),
.D(n_3539),
.Y(n_4058)
);

NAND3xp33_ASAP7_75t_L g4059 ( 
.A(n_4047),
.B(n_694),
.C(n_695),
.Y(n_4059)
);

NOR3xp33_ASAP7_75t_L g4060 ( 
.A(n_4032),
.B(n_696),
.C(n_697),
.Y(n_4060)
);

NOR2xp67_ASAP7_75t_L g4061 ( 
.A(n_4041),
.B(n_698),
.Y(n_4061)
);

AOI221xp5_ASAP7_75t_L g4062 ( 
.A1(n_4042),
.A2(n_3527),
.B1(n_3524),
.B2(n_3516),
.C(n_3553),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_4046),
.Y(n_4063)
);

OAI211xp5_ASAP7_75t_L g4064 ( 
.A1(n_4036),
.A2(n_698),
.B(n_699),
.C(n_700),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_4043),
.B(n_4038),
.Y(n_4065)
);

HB1xp67_ASAP7_75t_L g4066 ( 
.A(n_4045),
.Y(n_4066)
);

AOI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_4029),
.A2(n_3542),
.B1(n_3583),
.B2(n_3390),
.Y(n_4067)
);

NOR2x1_ASAP7_75t_L g4068 ( 
.A(n_4039),
.B(n_699),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_4051),
.B(n_700),
.Y(n_4069)
);

OR2x2_ASAP7_75t_L g4070 ( 
.A(n_4049),
.B(n_701),
.Y(n_4070)
);

AND4x1_ASAP7_75t_L g4071 ( 
.A(n_4044),
.B(n_701),
.C(n_702),
.D(n_703),
.Y(n_4071)
);

AND3x2_ASAP7_75t_L g4072 ( 
.A(n_4046),
.B(n_704),
.C(n_705),
.Y(n_4072)
);

INVx2_ASAP7_75t_L g4073 ( 
.A(n_4065),
.Y(n_4073)
);

XOR2xp5_ASAP7_75t_L g4074 ( 
.A(n_4052),
.B(n_4050),
.Y(n_4074)
);

AOI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_4061),
.A2(n_3583),
.B1(n_3542),
.B2(n_3589),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4054),
.Y(n_4076)
);

HB1xp67_ASAP7_75t_L g4077 ( 
.A(n_4066),
.Y(n_4077)
);

OAI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_4069),
.A2(n_4070),
.B1(n_4053),
.B2(n_4063),
.Y(n_4078)
);

NOR2xp33_ASAP7_75t_L g4079 ( 
.A(n_4055),
.B(n_705),
.Y(n_4079)
);

O2A1O1Ixp5_ASAP7_75t_L g4080 ( 
.A1(n_4064),
.A2(n_4059),
.B(n_4071),
.C(n_4072),
.Y(n_4080)
);

INVx2_ASAP7_75t_SL g4081 ( 
.A(n_4068),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_4067),
.Y(n_4082)
);

OAI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_4060),
.A2(n_3598),
.B(n_3543),
.Y(n_4083)
);

OAI311xp33_ASAP7_75t_L g4084 ( 
.A1(n_4056),
.A2(n_706),
.A3(n_707),
.B1(n_709),
.C1(n_710),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_4057),
.B(n_3522),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_4062),
.B(n_707),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_4058),
.A2(n_3583),
.B1(n_3542),
.B2(n_3577),
.Y(n_4087)
);

OR2x6_ASAP7_75t_L g4088 ( 
.A(n_4065),
.B(n_709),
.Y(n_4088)
);

INVxp67_ASAP7_75t_SL g4089 ( 
.A(n_4073),
.Y(n_4089)
);

AOI22xp5_ASAP7_75t_L g4090 ( 
.A1(n_4076),
.A2(n_3006),
.B1(n_3523),
.B2(n_3528),
.Y(n_4090)
);

AO22x1_ASAP7_75t_L g4091 ( 
.A1(n_4079),
.A2(n_4082),
.B1(n_4077),
.B2(n_4086),
.Y(n_4091)
);

AOI22xp5_ASAP7_75t_L g4092 ( 
.A1(n_4074),
.A2(n_3006),
.B1(n_3577),
.B2(n_3547),
.Y(n_4092)
);

BUFx6f_ASAP7_75t_L g4093 ( 
.A(n_4088),
.Y(n_4093)
);

AO22x2_ASAP7_75t_L g4094 ( 
.A1(n_4078),
.A2(n_3529),
.B1(n_3560),
.B2(n_3558),
.Y(n_4094)
);

AO22x2_ASAP7_75t_L g4095 ( 
.A1(n_4087),
.A2(n_4081),
.B1(n_4085),
.B2(n_4084),
.Y(n_4095)
);

AOI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_4088),
.A2(n_3598),
.B1(n_3556),
.B2(n_3561),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_4080),
.Y(n_4097)
);

AO22x2_ASAP7_75t_L g4098 ( 
.A1(n_4083),
.A2(n_3561),
.B1(n_3560),
.B2(n_3558),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4075),
.Y(n_4099)
);

AO22x2_ASAP7_75t_SL g4100 ( 
.A1(n_4073),
.A2(n_710),
.B1(n_711),
.B2(n_712),
.Y(n_4100)
);

NOR2xp67_ASAP7_75t_L g4101 ( 
.A(n_4073),
.B(n_711),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_4097),
.Y(n_4102)
);

XNOR2xp5_ASAP7_75t_L g4103 ( 
.A(n_4100),
.B(n_712),
.Y(n_4103)
);

HB1xp67_ASAP7_75t_L g4104 ( 
.A(n_4089),
.Y(n_4104)
);

AO21x2_ASAP7_75t_L g4105 ( 
.A1(n_4101),
.A2(n_4099),
.B(n_4091),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_4095),
.A2(n_713),
.B(n_714),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_4093),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_4093),
.Y(n_4108)
);

XNOR2xp5_ASAP7_75t_L g4109 ( 
.A(n_4094),
.B(n_713),
.Y(n_4109)
);

INVxp67_ASAP7_75t_L g4110 ( 
.A(n_4090),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4098),
.Y(n_4111)
);

HB1xp67_ASAP7_75t_L g4112 ( 
.A(n_4104),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_4102),
.Y(n_4113)
);

OAI22xp5_ASAP7_75t_SL g4114 ( 
.A1(n_4103),
.A2(n_4092),
.B1(n_4096),
.B2(n_717),
.Y(n_4114)
);

CKINVDCx20_ASAP7_75t_R g4115 ( 
.A(n_4105),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_4106),
.B(n_715),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_4109),
.B(n_4107),
.Y(n_4117)
);

OAI22x1_ASAP7_75t_L g4118 ( 
.A1(n_4108),
.A2(n_715),
.B1(n_716),
.B2(n_717),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_4113),
.B(n_4110),
.Y(n_4119)
);

AOI22x1_ASAP7_75t_L g4120 ( 
.A1(n_4112),
.A2(n_4111),
.B1(n_718),
.B2(n_719),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4116),
.Y(n_4121)
);

AOI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_4117),
.A2(n_4111),
.B(n_719),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_4118),
.B(n_716),
.Y(n_4123)
);

AOI32xp33_ASAP7_75t_L g4124 ( 
.A1(n_4119),
.A2(n_4115),
.A3(n_4114),
.B1(n_722),
.B2(n_723),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_4123),
.B(n_4121),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_SL g4126 ( 
.A(n_4124),
.B(n_4122),
.Y(n_4126)
);

AOI22xp33_ASAP7_75t_L g4127 ( 
.A1(n_4126),
.A2(n_4125),
.B1(n_4120),
.B2(n_3556),
.Y(n_4127)
);

OAI221xp5_ASAP7_75t_R g4128 ( 
.A1(n_4127),
.A2(n_720),
.B1(n_721),
.B2(n_724),
.C(n_725),
.Y(n_4128)
);

AOI211xp5_ASAP7_75t_L g4129 ( 
.A1(n_4128),
.A2(n_3511),
.B(n_3502),
.C(n_3489),
.Y(n_4129)
);


endmodule