module fake_jpeg_20639_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_17;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx4_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_9),
.B1(n_18),
.B2(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_10),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_19),
.B1(n_18),
.B2(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_16),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_31),
.B(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_34)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_37),
.B1(n_30),
.B2(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_42),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_21),
.C(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_43),
.C(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_34),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_37),
.B1(n_36),
.B2(n_14),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_49),
.B1(n_27),
.B2(n_26),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_53),
.B1(n_33),
.B2(n_12),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_50),
.B(n_45),
.C(n_48),
.D(n_21),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_12),
.B(n_13),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_56),
.B1(n_45),
.B2(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_17),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_17),
.B(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_60),
.B1(n_15),
.B2(n_8),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_68),
.B(n_64),
.C(n_69),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_2),
.Y(n_72)
);


endmodule