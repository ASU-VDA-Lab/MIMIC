module real_jpeg_17439_n_18 (n_559, n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_559;
input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_0),
.A2(n_34),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_0),
.A2(n_34),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_0),
.A2(n_34),
.B1(n_442),
.B2(n_444),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_78),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_1),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_1),
.A2(n_147),
.B1(n_261),
.B2(n_264),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_1),
.A2(n_147),
.B1(n_455),
.B2(n_458),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_1),
.A2(n_147),
.B1(n_466),
.B2(n_468),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_2),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_2),
.A2(n_160),
.B1(n_335),
.B2(n_338),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_2),
.A2(n_160),
.B1(n_550),
.B2(n_552),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_4),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_114),
.B1(n_118),
.B2(n_120),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_120),
.B1(n_190),
.B2(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_5),
.A2(n_120),
.B1(n_320),
.B2(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_6),
.A2(n_66),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_6),
.A2(n_66),
.B1(n_312),
.B2(n_315),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_6),
.A2(n_66),
.B1(n_402),
.B2(n_407),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_7),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_7),
.A2(n_228),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

OAI22x1_ASAP7_75t_SL g293 ( 
.A1(n_7),
.A2(n_228),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_7),
.A2(n_228),
.B1(n_313),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_8),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_8),
.A2(n_123),
.B1(n_287),
.B2(n_291),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_8),
.A2(n_123),
.B1(n_432),
.B2(n_437),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_8),
.A2(n_119),
.B1(n_123),
.B2(n_488),
.Y(n_487)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_9),
.Y(n_99)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_9),
.Y(n_349)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_10),
.B(n_150),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_10),
.A2(n_42),
.A3(n_270),
.B1(n_394),
.B2(n_397),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_10),
.B(n_72),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_10),
.A2(n_96),
.B1(n_233),
.B2(n_487),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_10),
.A2(n_76),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_11),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_12),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_12),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_12),
.A2(n_173),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_13),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_13),
.A2(n_105),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_13),
.A2(n_105),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_13),
.A2(n_105),
.B1(n_542),
.B2(n_545),
.Y(n_541)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_14),
.Y(n_84)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_14),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_14),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_14),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_16),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_16),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_17),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_17),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_17),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_528),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_374),
.B(n_523),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_305),
.C(n_369),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_253),
.B(n_278),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_24),
.B(n_253),
.C(n_525),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_151),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_25),
.B(n_152),
.C(n_221),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_73),
.C(n_121),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_27),
.B(n_121),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_41),
.B1(n_63),
.B2(n_71),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_29),
.A2(n_72),
.B1(n_260),
.B2(n_265),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_38),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_40),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_40),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_40),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_40),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_41),
.A2(n_63),
.B1(n_71),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_41),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_41),
.A2(n_71),
.B1(n_247),
.B2(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_41),
.A2(n_71),
.B1(n_286),
.B2(n_505),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_41),
.A2(n_71),
.B1(n_328),
.B2(n_549),
.Y(n_548)
);

AO21x2_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_48),
.B(n_56),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_55),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_57),
.Y(n_227)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_57),
.Y(n_337)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_61),
.Y(n_339)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_61),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_62),
.Y(n_272)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_72),
.A2(n_260),
.B1(n_265),
.B2(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_72),
.A2(n_265),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_73),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_95),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_74),
.B(n_95),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_89),
.B2(n_90),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_SL g267 ( 
.A1(n_75),
.A2(n_76),
.B(n_124),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_76),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_76),
.B(n_419),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_SL g429 ( 
.A1(n_76),
.A2(n_418),
.B(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_76),
.B(n_300),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_76),
.B(n_177),
.Y(n_493)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_80),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_80),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_88),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_130),
.B(n_134),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_94),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_102),
.B1(n_111),
.B2(n_113),
.Y(n_95)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_96),
.A2(n_113),
.B1(n_156),
.B2(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_96),
.A2(n_168),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_96),
.A2(n_166),
.B1(n_441),
.B2(n_449),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_96),
.A2(n_465),
.B1(n_487),
.B2(n_491),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_100),
.Y(n_416)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_101),
.Y(n_295)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_101),
.Y(n_406)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22x1_ASAP7_75t_SL g292 ( 
.A1(n_103),
.A2(n_154),
.B1(n_293),
.B2(n_299),
.Y(n_292)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_108),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_109),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_116),
.Y(n_407)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_117),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_117),
.Y(n_443)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_129),
.B1(n_145),
.B2(n_150),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_122),
.A2(n_129),
.B1(n_150),
.B2(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_129),
.Y(n_239)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_134),
.A2(n_239),
.B1(n_241),
.B2(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_134),
.A2(n_239),
.B1(n_311),
.B2(n_356),
.Y(n_355)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_140),
.B2(n_143),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_141),
.Y(n_322)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_146),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_150),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_221),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_174),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_153),
.A2(n_175),
.B(n_200),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_165),
.B2(n_167),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_154),
.A2(n_234),
.B1(n_293),
.B2(n_401),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_154),
.A2(n_464),
.B1(n_471),
.B2(n_472),
.Y(n_463)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_200),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_188),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_176),
.A2(n_201),
.B1(n_269),
.B2(n_277),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_176),
.A2(n_201),
.B1(n_333),
.B2(n_340),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_176),
.A2(n_201),
.B1(n_429),
.B2(n_431),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_176),
.A2(n_201),
.B1(n_431),
.B2(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_176),
.A2(n_201),
.B1(n_384),
.B2(n_454),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_176),
.A2(n_201),
.B(n_340),
.Y(n_554)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_177),
.A2(n_214),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_177),
.A2(n_189),
.B1(n_224),
.B2(n_334),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_177),
.A2(n_224),
.B1(n_383),
.B2(n_390),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_182),
.B1(n_183),
.B2(n_186),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_185),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_185),
.Y(n_467)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_185),
.Y(n_484)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_187),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_213),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_207),
.B1(n_210),
.B2(n_212),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_206),
.Y(n_342)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_206),
.Y(n_389)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_210),
.Y(n_417)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_216),
.Y(n_343)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_237),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_222),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_232),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_225),
.Y(n_277)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_230),
.Y(n_459)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_233),
.Y(n_471)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_238),
.B(n_246),
.C(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_239),
.A2(n_240),
.B1(n_356),
.B2(n_541),
.Y(n_540)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_251),
.Y(n_553)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_252),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_255),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_258),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.C(n_268),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_268),
.Y(n_281)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_281),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_269),
.Y(n_390)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_275),
.Y(n_398)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_302),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_279),
.B(n_302),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.C(n_283),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_280),
.B(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_282),
.B(n_283),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.C(n_301),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_284),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_290),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_292),
.B(n_301),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_294),
.Y(n_488)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

A2O1A1O1Ixp25_ASAP7_75t_L g523 ( 
.A1(n_305),
.A2(n_369),
.B(n_524),
.C(n_526),
.D(n_527),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_360),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_306),
.B(n_360),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_323),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_307),
.B(n_531),
.C(n_532),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.C(n_316),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_363),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_316),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_312),
.Y(n_315)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_314),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_320),
.Y(n_506)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_320),
.Y(n_551)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_345),
.Y(n_323)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_324),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_332),
.B(n_344),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_332),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_344),
.A2(n_538),
.B1(n_555),
.B2(n_556),
.Y(n_537)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_344),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_345),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_351),
.B1(n_352),
.B2(n_359),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_346),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_347),
.A2(n_350),
.B1(n_353),
.B2(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_349),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_353),
.A2(n_359),
.B1(n_535),
.B2(n_559),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_354),
.Y(n_536)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx5_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_366),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_362),
.B1(n_364),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_364),
.Y(n_372)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_373),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_370),
.B(n_373),
.Y(n_526)
);

AOI21x1_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_408),
.B(n_522),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_376),
.B(n_378),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.C(n_391),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_379),
.A2(n_380),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_382),
.A2(n_391),
.B1(n_392),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_382),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_399),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_393),
.A2(n_399),
.B1(n_400),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_515),
.B(n_521),
.Y(n_408)
);

AOI21x1_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_497),
.B(n_514),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_461),
.B(n_496),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_439),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_412),
.B(n_439),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_427),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_413),
.A2(n_427),
.B1(n_428),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_416),
.A3(n_417),
.B1(n_418),
.B2(n_420),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_436),
.Y(n_438)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_450),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_452),
.C(n_460),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_453),
.B2(n_460),
.Y(n_450)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_475),
.B(n_495),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_473),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_473),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_470),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_489),
.B(n_494),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_486),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_485),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_493),
.Y(n_494)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_499),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_503),
.C(n_513),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_512),
.B2(n_513),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_520),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_520),
.Y(n_521)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_557),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_533),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_530),
.B(n_533),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_537),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_538),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_547),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_554),
.Y(n_547)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);


endmodule