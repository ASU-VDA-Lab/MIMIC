module fake_jpeg_13416_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_0),
.B(n_6),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_56),
.Y(n_156)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_94),
.Y(n_120)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_95),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_29),
.B(n_17),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_98),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_100),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_25),
.B(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_25),
.B(n_16),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_33),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_28),
.B(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_113),
.B(n_114),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_116),
.B(n_124),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_28),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_133),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_67),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_106),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_26),
.C(n_34),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_136),
.B(n_137),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_153),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_75),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_59),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_175),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_58),
.A2(n_33),
.B1(n_26),
.B2(n_38),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_157),
.A2(n_58),
.B1(n_68),
.B2(n_26),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_61),
.B(n_46),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_81),
.B(n_46),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_88),
.A2(n_90),
.B1(n_102),
.B2(n_93),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_20),
.B1(n_38),
.B2(n_44),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_84),
.Y(n_175)
);

INVx2_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

OR2x4_ASAP7_75t_L g290 ( 
.A(n_177),
.B(n_140),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_178),
.B(n_196),
.Y(n_263)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_179),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_64),
.B1(n_66),
.B2(n_71),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_182),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_275)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx6_ASAP7_75t_SL g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_192),
.Y(n_265)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_51),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_198),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_120),
.B(n_37),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_117),
.B(n_96),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_197),
.B(n_202),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_51),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_111),
.B(n_37),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_199),
.B(n_200),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_206),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_135),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_173),
.A2(n_82),
.B1(n_79),
.B2(n_86),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_115),
.A2(n_85),
.B1(n_83),
.B2(n_53),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_129),
.B(n_92),
.Y(n_216)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_112),
.Y(n_219)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_135),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_131),
.B(n_34),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_230),
.Y(n_250)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_154),
.A2(n_41),
.B1(n_68),
.B2(n_110),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_225),
.A2(n_228),
.B1(n_240),
.B2(n_132),
.Y(n_259)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_156),
.A2(n_41),
.B1(n_110),
.B2(n_53),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_118),
.B(n_20),
.C(n_44),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_229),
.B(n_231),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_118),
.B(n_14),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_133),
.A2(n_20),
.B1(n_52),
.B2(n_3),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_208),
.B1(n_157),
.B2(n_202),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_127),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_156),
.B(n_14),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_234),
.Y(n_268)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_235),
.Y(n_291)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_146),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_237),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_152),
.B(n_14),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_158),
.B(n_12),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_244),
.A2(n_260),
.B1(n_294),
.B2(n_197),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_180),
.A2(n_128),
.B1(n_149),
.B2(n_141),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_245),
.A2(n_287),
.B1(n_219),
.B2(n_191),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_172),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_273),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_259),
.A2(n_274),
.B1(n_243),
.B2(n_282),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_229),
.A2(n_126),
.B1(n_169),
.B2(n_119),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_198),
.B(n_126),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_206),
.A2(n_132),
.B1(n_147),
.B2(n_158),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_184),
.B(n_180),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_128),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_217),
.A2(n_149),
.B1(n_165),
.B2(n_119),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_187),
.B(n_167),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_289),
.B(n_265),
.Y(n_324)
);

INVx6_ASAP7_75t_SL g331 ( 
.A(n_290),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_181),
.A2(n_147),
.B(n_174),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_190),
.B(n_201),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_223),
.A2(n_150),
.B1(n_169),
.B2(n_162),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_197),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_297),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_210),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_298),
.A2(n_310),
.B(n_317),
.Y(n_373)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_193),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_308),
.C(n_340),
.Y(n_351)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_236),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_302),
.B(n_306),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_304),
.A2(n_315),
.B1(n_346),
.B2(n_285),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_277),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_192),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_188),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_316),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_243),
.A2(n_227),
.B1(n_224),
.B2(n_167),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_241),
.A2(n_138),
.B1(n_150),
.B2(n_162),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_311),
.A2(n_312),
.B1(n_322),
.B2(n_271),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_138),
.B1(n_140),
.B2(n_185),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_237),
.B1(n_235),
.B2(n_231),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_313),
.A2(n_294),
.B1(n_288),
.B2(n_293),
.Y(n_348)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_244),
.A2(n_203),
.B1(n_194),
.B2(n_186),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_177),
.C(n_188),
.Y(n_316)
);

AO22x1_ASAP7_75t_SL g318 ( 
.A1(n_255),
.A2(n_221),
.B1(n_205),
.B2(n_189),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_318),
.B(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_250),
.B(n_240),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_323),
.Y(n_356)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_252),
.B(n_179),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_325),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_251),
.B(n_222),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_290),
.Y(n_329)
);

INVx3_ASAP7_75t_SL g330 ( 
.A(n_242),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_330),
.A2(n_337),
.B1(n_344),
.B2(n_345),
.Y(n_366)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_250),
.B(n_212),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_333),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_262),
.Y(n_334)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_242),
.Y(n_335)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_249),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_269),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_251),
.B(n_212),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_339),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_127),
.Y(n_340)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_254),
.B(n_207),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_341),
.A2(n_270),
.B(n_257),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_253),
.B(n_171),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_343),
.Y(n_379)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

BUFx12_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_256),
.B(n_1),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_260),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_341),
.B(n_317),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_347),
.A2(n_352),
.B(n_4),
.Y(n_422)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_284),
.B(n_292),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_284),
.B(n_288),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_SL g409 ( 
.A1(n_355),
.A2(n_372),
.B(n_375),
.C(n_344),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_304),
.A2(n_283),
.B1(n_288),
.B2(n_264),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_368),
.B1(n_318),
.B2(n_322),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_308),
.A2(n_264),
.B1(n_291),
.B2(n_295),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_363),
.A2(n_364),
.B1(n_327),
.B2(n_343),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_303),
.A2(n_258),
.B1(n_286),
.B2(n_281),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_300),
.B(n_285),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_370),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_322),
.B1(n_297),
.B2(n_318),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_305),
.B(n_278),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_315),
.A2(n_266),
.B(n_270),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_280),
.B(n_296),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_374),
.A2(n_301),
.B(n_299),
.Y(n_411)
);

FAx1_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_296),
.CI(n_261),
.CON(n_375),
.SN(n_375)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_337),
.B(n_314),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_303),
.B(n_257),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_384),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_261),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_298),
.B(n_280),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_346),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_353),
.B(n_307),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_390),
.B(n_405),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_379),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_395),
.Y(n_438)
);

NOR3xp33_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_297),
.C(n_319),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_392),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_417),
.B1(n_419),
.B2(n_424),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_379),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_397),
.A2(n_388),
.B1(n_378),
.B2(n_377),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_398),
.A2(n_359),
.B1(n_375),
.B2(n_361),
.Y(n_444)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_400),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_401),
.B(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_338),
.Y(n_402)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_402),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_358),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_414),
.Y(n_457)
);

OA22x2_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_322),
.B1(n_321),
.B2(n_336),
.Y(n_404)
);

OA22x2_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_409),
.B1(n_425),
.B2(n_363),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_334),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_408),
.A2(n_423),
.B(n_427),
.Y(n_432)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_422),
.B(n_352),
.Y(n_443)
);

BUFx12_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_412),
.Y(n_448)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_413),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_335),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_381),
.B(n_330),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_415),
.B(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_386),
.B(n_344),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_356),
.B(n_1),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_362),
.B(n_2),
.Y(n_419)
);

BUFx12f_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_2),
.Y(n_421)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_387),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_389),
.B(n_4),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_SL g425 ( 
.A1(n_355),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_7),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_371),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_347),
.A2(n_9),
.B(n_10),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_396),
.A2(n_368),
.B1(n_357),
.B2(n_387),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_428),
.A2(n_444),
.B1(n_445),
.B2(n_449),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_351),
.C(n_365),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_446),
.C(n_433),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_434),
.B(n_428),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_374),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g470 ( 
.A1(n_435),
.A2(n_409),
.B(n_404),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_425),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_443),
.A2(n_427),
.B(n_423),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_396),
.A2(n_372),
.B1(n_375),
.B2(n_361),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_370),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_451),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_421),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_398),
.A2(n_372),
.B1(n_376),
.B2(n_373),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_394),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_348),
.Y(n_452)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_452),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_366),
.B1(n_373),
.B2(n_388),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_455),
.A2(n_406),
.B1(n_407),
.B2(n_404),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_426),
.A2(n_378),
.B1(n_377),
.B2(n_385),
.Y(n_456)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_408),
.A2(n_369),
.B(n_371),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_458),
.A2(n_422),
.B(n_406),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_461),
.A2(n_481),
.B(n_441),
.C(n_444),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_420),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_462),
.B(n_466),
.Y(n_489)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_438),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_451),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_467),
.Y(n_497)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_468),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_394),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_472),
.A2(n_461),
.B(n_432),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_409),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_477),
.C(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_460),
.B(n_385),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_476),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_409),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_447),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_479),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_455),
.A2(n_404),
.B1(n_418),
.B2(n_413),
.Y(n_480)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_400),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_484),
.C(n_441),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_433),
.B(n_410),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_483),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_449),
.B(n_369),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_435),
.A2(n_425),
.B(n_412),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_458),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_420),
.Y(n_488)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_491),
.B(n_490),
.Y(n_513)
);

INVx13_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

AO21x1_ASAP7_75t_L g529 ( 
.A1(n_495),
.A2(n_496),
.B(n_502),
.Y(n_529)
);

XOR2x1_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_484),
.Y(n_517)
);

NOR2x1_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_430),
.Y(n_501)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_501),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_430),
.C(n_443),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_506),
.B(n_508),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_465),
.B(n_437),
.C(n_441),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_480),
.Y(n_511)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_468),
.Y(n_512)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_512),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_490),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_437),
.Y(n_514)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_514),
.Y(n_535)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_502),
.A2(n_473),
.B(n_482),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_518),
.A2(n_523),
.B(n_496),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_498),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_522),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_501),
.A2(n_481),
.B(n_470),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_520),
.A2(n_529),
.B(n_432),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_497),
.B(n_474),
.Y(n_522)
);

FAx1_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_481),
.CI(n_472),
.CON(n_523),
.SN(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_485),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_524),
.B(n_526),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_475),
.C(n_477),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_499),
.B(n_469),
.C(n_463),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_528),
.C(n_500),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_453),
.C(n_481),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_516),
.A2(n_512),
.B1(n_493),
.B2(n_503),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_532),
.A2(n_531),
.B1(n_515),
.B2(n_530),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_507),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_534),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_514),
.A2(n_493),
.B1(n_492),
.B2(n_510),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_531),
.A2(n_511),
.B1(n_503),
.B2(n_495),
.Y(n_536)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_536),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_509),
.Y(n_538)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_538),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_539),
.A2(n_543),
.B(n_545),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_540),
.B(n_542),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_527),
.B(n_508),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_492),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_544),
.B(n_541),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_509),
.C(n_500),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_546),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_548),
.B(n_517),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_532),
.A2(n_530),
.B1(n_525),
.B2(n_520),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_551),
.A2(n_556),
.B1(n_538),
.B2(n_536),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_526),
.C(n_518),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_555),
.B(n_557),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_535),
.A2(n_523),
.B1(n_436),
.B2(n_529),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_453),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_420),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_554),
.A2(n_545),
.B1(n_547),
.B2(n_543),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_561),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_542),
.C(n_539),
.Y(n_561)
);

AOI322xp5_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_564),
.A3(n_494),
.B1(n_562),
.B2(n_550),
.C1(n_558),
.C2(n_412),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_566),
.C(n_551),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_549),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_567),
.B(n_568),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_561),
.A2(n_552),
.B(n_558),
.C(n_556),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_570),
.B(n_566),
.Y(n_572)
);

AOI322xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_569),
.A3(n_523),
.B1(n_565),
.B2(n_504),
.C1(n_442),
.C2(n_548),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_573),
.B(n_574),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_571),
.B(n_500),
.C(n_504),
.Y(n_574)
);

AOI322xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_429),
.A3(n_440),
.B1(n_439),
.B2(n_500),
.C1(n_459),
.C2(n_383),
.Y(n_576)
);

OAI321xp33_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_349),
.A3(n_383),
.B1(n_459),
.B2(n_425),
.C(n_11),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_349),
.B(n_9),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_11),
.Y(n_579)
);


endmodule