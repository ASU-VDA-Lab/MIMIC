module fake_jpeg_31437_n_431 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g148 ( 
.A(n_48),
.Y(n_148)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_16),
.A2(n_8),
.B1(n_1),
.B2(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_74),
.B1(n_41),
.B2(n_42),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_14),
.B(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_70),
.Y(n_137)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_16),
.A2(n_13),
.B1(n_1),
.B2(n_3),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_26),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_3),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_24),
.B(n_5),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_88),
.Y(n_120)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_24),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_91),
.Y(n_147)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_20),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_150),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_32),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_121),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_32),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_135),
.B1(n_74),
.B2(n_68),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_134),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_20),
.B1(n_47),
.B2(n_40),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_128),
.A2(n_143),
.B1(n_156),
.B2(n_81),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_53),
.B(n_47),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_41),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_45),
.B1(n_40),
.B2(n_33),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_92),
.A2(n_79),
.B1(n_84),
.B2(n_82),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_75),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_152),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_49),
.A2(n_65),
.B1(n_56),
.B2(n_85),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_60),
.B1(n_33),
.B2(n_45),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_159),
.Y(n_233)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_39),
.B1(n_29),
.B2(n_26),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_100),
.A2(n_51),
.B1(n_70),
.B2(n_54),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_169),
.A2(n_137),
.B1(n_125),
.B2(n_136),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_178),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_113),
.A2(n_71),
.B1(n_20),
.B2(n_151),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_175),
.A2(n_176),
.B1(n_188),
.B2(n_189),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_20),
.B1(n_46),
.B2(n_36),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_185),
.B1(n_197),
.B2(n_137),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_73),
.C(n_59),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_187),
.C(n_193),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_48),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_101),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_192),
.B(n_195),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_114),
.B(n_29),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_196),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_111),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_91),
.C(n_15),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_198),
.Y(n_204)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_135),
.A2(n_97),
.B1(n_15),
.B2(n_83),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_144),
.B1(n_151),
.B2(n_153),
.Y(n_230)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_210),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_133),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_212),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_133),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_128),
.A3(n_143),
.B1(n_156),
.B2(n_119),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_158),
.B(n_163),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_102),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_227),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_232),
.B1(n_158),
.B2(n_170),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_106),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_161),
.B1(n_189),
.B2(n_172),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_120),
.B(n_123),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_169),
.B(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_170),
.B(n_149),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_21),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_184),
.B1(n_180),
.B2(n_188),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_SL g283 ( 
.A1(n_240),
.A2(n_244),
.B(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_245),
.B1(n_260),
.B2(n_263),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_250),
.C(n_261),
.Y(n_266)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_167),
.B1(n_140),
.B2(n_154),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_158),
.B1(n_169),
.B2(n_177),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_263),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_165),
.B(n_120),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_205),
.Y(n_280)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_249),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_173),
.C(n_162),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_181),
.B1(n_168),
.B2(n_142),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_256),
.Y(n_276)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

AO22x1_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_174),
.B1(n_124),
.B2(n_118),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_224),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_199),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_195),
.C(n_160),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_227),
.C(n_217),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_217),
.B(n_225),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_277),
.B(n_248),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_206),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_217),
.B(n_235),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_246),
.B(n_211),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_278),
.B(n_279),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_209),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_285),
.B1(n_261),
.B2(n_242),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_201),
.Y(n_282)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_259),
.B(n_207),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_286),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_245),
.A2(n_232),
.B1(n_207),
.B2(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_204),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_243),
.B1(n_231),
.B2(n_251),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_241),
.B1(n_259),
.B2(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_305),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_292),
.B(n_301),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_293),
.A2(n_294),
.B1(n_299),
.B2(n_267),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_283),
.B1(n_281),
.B2(n_276),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_250),
.C(n_254),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_303),
.C(n_304),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_276),
.B1(n_280),
.B2(n_278),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_258),
.A3(n_253),
.B1(n_249),
.B2(n_203),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_258),
.B(n_226),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_233),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_224),
.C(n_203),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_266),
.B(n_226),
.C(n_239),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_218),
.B(n_229),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_264),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_311),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_202),
.B1(n_39),
.B2(n_46),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_229),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_231),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_279),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_314),
.B(n_325),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_273),
.B1(n_275),
.B2(n_274),
.Y(n_316)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_277),
.B1(n_267),
.B2(n_286),
.Y(n_319)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_279),
.C(n_277),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_328),
.C(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_291),
.A2(n_300),
.B1(n_301),
.B2(n_296),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_326),
.A2(n_311),
.B1(n_310),
.B2(n_288),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_21),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_271),
.C(n_268),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_271),
.C(n_268),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_272),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_298),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_270),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_214),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_312),
.C(n_293),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_306),
.C(n_289),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_342),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_311),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_338),
.B(n_320),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_339),
.B(n_340),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_305),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_352),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_265),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_265),
.B1(n_214),
.B2(n_36),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_347),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_223),
.Y(n_346)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_346),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_330),
.B(n_38),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_21),
.C(n_109),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_322),
.C(n_327),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_329),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_356),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_318),
.B(n_109),
.Y(n_356)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_334),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_336),
.C(n_354),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_325),
.B1(n_335),
.B2(n_320),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_363),
.A2(n_341),
.B1(n_335),
.B2(n_351),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_366),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_369),
.B(n_339),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_332),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_315),
.Y(n_372)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_385),
.C(n_361),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_357),
.B1(n_5),
.B2(n_6),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_313),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_380),
.Y(n_396)
);

AOI21x1_ASAP7_75t_SL g383 ( 
.A1(n_363),
.A2(n_340),
.B(n_338),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_383),
.A2(n_333),
.B(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_384),
.B(n_386),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_328),
.C(n_354),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_387),
.B(n_359),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_377),
.A2(n_362),
.B1(n_365),
.B2(n_358),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_390),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_392),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_393),
.B(n_397),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_382),
.B(n_370),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_395),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_362),
.B(n_313),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_377),
.A2(n_349),
.B1(n_352),
.B2(n_357),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_399),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_381),
.A2(n_44),
.B1(n_6),
.B2(n_9),
.Y(n_399)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_378),
.Y(n_401)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_385),
.C(n_374),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_403),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_391),
.B(n_375),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_396),
.B(n_384),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_409),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_379),
.Y(n_409)
);

AOI21xp33_ASAP7_75t_L g410 ( 
.A1(n_400),
.A2(n_388),
.B(n_395),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_410),
.A2(n_413),
.B(n_416),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_390),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_417),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_402),
.A2(n_397),
.B(n_6),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_412),
.B(n_10),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_407),
.A2(n_10),
.B(n_11),
.Y(n_413)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_408),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

AOI21xp33_ASAP7_75t_L g420 ( 
.A1(n_415),
.A2(n_407),
.B(n_404),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_421),
.C(n_44),
.Y(n_424)
);

OAI21xp33_ASAP7_75t_L g421 ( 
.A1(n_417),
.A2(n_401),
.B(n_10),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_411),
.C(n_414),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_423),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_425),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_426),
.A2(n_419),
.B(n_11),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_427),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_21),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_0),
.B(n_21),
.Y(n_431)
);


endmodule