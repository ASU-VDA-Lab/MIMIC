module fake_jpeg_16682_n_393 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_3),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_2),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_39),
.B(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_49),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_18),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_50),
.A2(n_16),
.B1(n_5),
.B2(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_65),
.Y(n_98)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_57),
.Y(n_109)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_7),
.C(n_12),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_16),
.C(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_26),
.B(n_36),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_13),
.B1(n_8),
.B2(n_7),
.Y(n_130)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_18),
.B1(n_37),
.B2(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_18),
.B1(n_37),
.B2(n_31),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_37),
.B1(n_36),
.B2(n_32),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_88),
.B(n_115),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_32),
.B1(n_22),
.B2(n_23),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_103),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_19),
.B(n_28),
.C(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_93),
.B(n_107),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_22),
.B1(n_28),
.B2(n_25),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_39),
.A2(n_28),
.B1(n_25),
.B2(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_34),
.B1(n_30),
.B2(n_14),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_19),
.B(n_14),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_66),
.Y(n_138)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_65),
.A2(n_14),
.B1(n_30),
.B2(n_16),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_84),
.B1(n_68),
.B2(n_72),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_10),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_118),
.A2(n_121),
.B1(n_161),
.B2(n_129),
.Y(n_208)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_59),
.B1(n_54),
.B2(n_26),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_126),
.B(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_35),
.B1(n_33),
.B2(n_17),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_127),
.A2(n_142),
.B1(n_156),
.B2(n_165),
.Y(n_194)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_128),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_83),
.B(n_5),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_131),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_147),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_86),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_149),
.B1(n_155),
.B2(n_67),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_143),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_138),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_76),
.A2(n_87),
.B1(n_75),
.B2(n_82),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_80),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_10),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_84),
.A2(n_33),
.B1(n_10),
.B2(n_4),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_48),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_17),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_151),
.B(n_157),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_101),
.B1(n_70),
.B2(n_71),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_153),
.A2(n_164),
.B1(n_132),
.B2(n_122),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_91),
.A2(n_86),
.B1(n_104),
.B2(n_108),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_5),
.B1(n_8),
.B2(n_2),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_70),
.B(n_61),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_71),
.B(n_8),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_118),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_95),
.A2(n_46),
.B1(n_57),
.B2(n_8),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_102),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_78),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_0),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_159),
.Y(n_205)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_77),
.A2(n_1),
.B1(n_3),
.B2(n_67),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_1),
.B1(n_156),
.B2(n_130),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_1),
.B(n_97),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_171),
.A2(n_173),
.B(n_154),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_148),
.B(n_147),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_175),
.B(n_198),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_191),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_97),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_192),
.C(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_110),
.B(n_102),
.C(n_116),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_179),
.B(n_184),
.Y(n_251)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_116),
.C(n_1),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_122),
.B1(n_141),
.B2(n_171),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_199),
.B(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_140),
.B(n_160),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_157),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_205),
.B(n_172),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_208),
.B1(n_180),
.B2(n_192),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_186),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_127),
.A2(n_153),
.B1(n_144),
.B2(n_125),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_216),
.B1(n_134),
.B2(n_126),
.Y(n_228)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_120),
.Y(n_230)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_119),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_142),
.B(n_144),
.C(n_159),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_153),
.A2(n_119),
.B1(n_164),
.B2(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_219),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_201),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_153),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_234),
.B1(n_253),
.B2(n_254),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_224),
.A2(n_248),
.B(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_228),
.A2(n_218),
.B1(n_249),
.B2(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_141),
.C(n_158),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_246),
.C(n_239),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_206),
.B1(n_198),
.B2(n_194),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_135),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_240),
.A2(n_241),
.B1(n_249),
.B2(n_250),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_211),
.B1(n_214),
.B2(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_173),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_256),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_187),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_188),
.A2(n_207),
.B1(n_197),
.B2(n_183),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_207),
.A2(n_193),
.B1(n_178),
.B2(n_179),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_250),
.B(n_256),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_190),
.A2(n_207),
.B1(n_176),
.B2(n_212),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_172),
.A2(n_210),
.B1(n_204),
.B2(n_174),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_229),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_182),
.B(n_174),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_181),
.A2(n_213),
.B1(n_182),
.B2(n_215),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_217),
.B1(n_247),
.B2(n_231),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_200),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_200),
.B(n_213),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g311 ( 
.A1(n_260),
.A2(n_277),
.B1(n_263),
.B2(n_269),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_261),
.B(n_266),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_263),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_265),
.A2(n_269),
.B(n_272),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_233),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_268),
.A2(n_275),
.B1(n_280),
.B2(n_292),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_217),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_270),
.B(n_271),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_231),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_228),
.B1(n_224),
.B2(n_246),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_242),
.A2(n_243),
.B1(n_219),
.B2(n_235),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_225),
.B(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_274),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g277 ( 
.A(n_254),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_220),
.B(n_244),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_278),
.A2(n_284),
.B(n_288),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_226),
.B1(n_251),
.B2(n_230),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_282),
.B(n_283),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_235),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_226),
.B(n_237),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_221),
.A2(n_243),
.B1(n_238),
.B2(n_237),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_286),
.A2(n_275),
.B1(n_260),
.B2(n_273),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_238),
.A2(n_252),
.B(n_239),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_262),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_225),
.B(n_173),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_291),
.B(n_276),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_234),
.A2(n_248),
.B1(n_223),
.B2(n_222),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_293),
.B(n_312),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_308),
.C(n_314),
.Y(n_323)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_307),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_298),
.A2(n_302),
.B(n_311),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_265),
.C(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_299),
.B(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_259),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_305),
.Y(n_331)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_264),
.C(n_284),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_292),
.B(n_259),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_281),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_285),
.B1(n_284),
.B2(n_269),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_313),
.A2(n_317),
.B1(n_283),
.B2(n_310),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_311),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_321),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_272),
.A2(n_260),
.B1(n_285),
.B2(n_267),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_262),
.B(n_273),
.C(n_291),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_282),
.C(n_270),
.Y(n_325)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_260),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_325),
.C(n_328),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_261),
.C(n_266),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_271),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_339),
.C(n_315),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_332),
.B(n_304),
.Y(n_357)
);

OA21x2_ASAP7_75t_SL g333 ( 
.A1(n_299),
.A2(n_319),
.B(n_293),
.Y(n_333)
);

XNOR2x2_ASAP7_75t_SL g348 ( 
.A(n_333),
.B(n_301),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_317),
.A2(n_302),
.B1(n_313),
.B2(n_305),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_335),
.B1(n_307),
.B2(n_312),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_306),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_300),
.Y(n_341)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_341),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_309),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_318),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_318),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_359),
.C(n_322),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_311),
.B(n_301),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_347),
.B(n_357),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_R g371 ( 
.A(n_348),
.B(n_338),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_352),
.B(n_353),
.Y(n_361)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_356),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_311),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_330),
.Y(n_368)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_358),
.B(n_350),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_321),
.C(n_296),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_298),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_362),
.Y(n_374)
);

XOR2x2_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_371),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_366),
.C(n_368),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_328),
.C(n_325),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_343),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_336),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_378),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_367),
.A2(n_331),
.B1(n_347),
.B2(n_351),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_375),
.A2(n_360),
.B1(n_363),
.B2(n_346),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_369),
.C(n_357),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_377),
.B(n_364),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);

AOI221xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_377),
.B1(n_374),
.B2(n_379),
.C(n_334),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_385),
.A2(n_360),
.B(n_345),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_384),
.A2(n_374),
.B(n_337),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_386),
.A2(n_387),
.B(n_382),
.Y(n_388)
);

A2O1A1O1Ixp25_ASAP7_75t_L g389 ( 
.A1(n_388),
.A2(n_376),
.B(n_380),
.C(n_348),
.D(n_369),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_389),
.A2(n_344),
.B1(n_376),
.B2(n_383),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_344),
.B(n_364),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_355),
.B(n_327),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_332),
.Y(n_393)
);


endmodule