module fake_jpeg_15570_n_98 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_98);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_9),
.B1(n_13),
.B2(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_4),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_9),
.B1(n_16),
.B2(n_12),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_18),
.B1(n_15),
.B2(n_10),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_25),
.B1(n_19),
.B2(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_11),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_22),
.C(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_9),
.B1(n_18),
.B2(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_33),
.B1(n_28),
.B2(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_28),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_26),
.B(n_25),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_45),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_44),
.C(n_39),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_41),
.C(n_36),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_52),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_65),
.C(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_69),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_36),
.C(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_54),
.B(n_57),
.Y(n_71)
);

AOI31xp33_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_76),
.A3(n_24),
.B(n_7),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_24),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_8),
.C(n_12),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_8),
.B(n_12),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_62),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_17),
.C(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_14),
.B(n_5),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_35),
.B1(n_27),
.B2(n_2),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_86),
.Y(n_90)
);

NAND4xp25_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_35),
.C(n_17),
.D(n_21),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_79),
.A3(n_81),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_91),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_6),
.A3(n_7),
.B1(n_21),
.B2(n_1),
.C1(n_0),
.C2(n_14),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_R g96 ( 
.A(n_93),
.B(n_0),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_6),
.B(n_0),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_1),
.C(n_95),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);


endmodule