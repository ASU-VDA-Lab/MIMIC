module real_aes_2124_n_383 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_383);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_383;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_905;
wire n_673;
wire n_518;
wire n_792;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_666;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_948;
wire n_1021;
wire n_399;
wire n_700;
wire n_958;
wire n_677;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_755;
wire n_1025;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_649;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1028;
wire n_1003;
wire n_727;
wire n_1014;
wire n_1056;
wire n_749;
wire n_385;
wire n_397;
wire n_663;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_393;
wire n_703;
wire n_652;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_0), .A2(n_235), .B1(n_753), .B2(n_845), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_1), .A2(n_69), .B1(n_488), .B2(n_625), .Y(n_980) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_2), .A2(n_117), .B1(n_602), .B2(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_3), .A2(n_128), .B1(n_695), .B2(n_822), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_4), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_5), .A2(n_254), .B1(n_458), .B2(n_566), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_6), .A2(n_78), .B1(n_485), .B2(n_860), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_7), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_8), .A2(n_342), .B1(n_816), .B2(n_817), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_9), .A2(n_67), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_10), .A2(n_376), .B1(n_469), .B2(n_472), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_11), .A2(n_210), .B1(n_759), .B2(n_761), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_12), .A2(n_198), .B1(n_599), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_13), .A2(n_260), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_14), .A2(n_301), .B1(n_592), .B2(n_594), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_15), .A2(n_317), .B1(n_455), .B2(n_653), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_16), .A2(n_86), .B1(n_862), .B2(n_863), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_17), .A2(n_138), .B1(n_488), .B2(n_625), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_18), .A2(n_189), .B1(n_459), .B2(n_566), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_19), .A2(n_195), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_20), .A2(n_259), .B1(n_519), .B2(n_520), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_21), .B(n_665), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_22), .A2(n_100), .B1(n_653), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_23), .A2(n_296), .B1(n_836), .B2(n_837), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_24), .A2(n_258), .B1(n_462), .B2(n_464), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_25), .B(n_394), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_26), .A2(n_284), .B1(n_651), .B2(n_848), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_27), .A2(n_147), .B1(n_470), .B2(n_884), .Y(n_883) );
INVx1_ASAP7_75t_SL g401 ( .A(n_28), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g1027 ( .A(n_28), .B(n_43), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_29), .A2(n_119), .B1(n_525), .B2(n_559), .Y(n_626) );
AOI22xp5_ASAP7_75t_SL g945 ( .A1(n_30), .A2(n_262), .B1(n_645), .B2(n_778), .Y(n_945) );
AOI222xp33_ASAP7_75t_L g982 ( .A1(n_31), .A2(n_311), .B1(n_347), .B2(n_574), .C1(n_983), .C2(n_984), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_32), .B(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_33), .A2(n_37), .B1(n_653), .B2(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_34), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_35), .A2(n_223), .B1(n_772), .B2(n_773), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_36), .A2(n_299), .B1(n_671), .B2(n_738), .Y(n_928) );
XNOR2x1_ASAP7_75t_SL g852 ( .A(n_38), .B(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_SL g893 ( .A1(n_38), .A2(n_853), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_38), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_39), .A2(n_265), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_40), .A2(n_109), .B1(n_473), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_41), .A2(n_104), .B1(n_825), .B2(n_826), .Y(n_824) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_42), .A2(n_389), .B(n_477), .Y(n_388) );
INVx1_ASAP7_75t_L g479 ( .A(n_42), .Y(n_479) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_43), .A2(n_353), .B1(n_400), .B2(n_404), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_44), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_45), .A2(n_294), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_46), .A2(n_110), .B1(n_599), .B2(n_698), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_47), .A2(n_194), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_48), .A2(n_96), .B1(n_530), .B2(n_531), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_49), .A2(n_280), .B1(n_657), .B2(n_890), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_50), .A2(n_116), .B1(n_758), .B2(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_51), .A2(n_283), .B1(n_879), .B2(n_880), .Y(n_878) );
INVx1_ASAP7_75t_L g402 ( .A(n_52), .Y(n_402) );
AO222x2_ASAP7_75t_SL g622 ( .A1(n_53), .A2(n_211), .B1(n_288), .B2(n_518), .C1(n_519), .C2(n_520), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_54), .A2(n_343), .B1(n_414), .B2(n_491), .Y(n_811) );
INVx1_ASAP7_75t_L g933 ( .A(n_55), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_56), .A2(n_252), .B1(n_506), .B2(n_507), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_57), .A2(n_274), .B1(n_674), .B2(n_675), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_58), .B(n_731), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_59), .A2(n_242), .B1(n_698), .B2(n_699), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_60), .A2(n_98), .B1(n_695), .B2(n_696), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_61), .A2(n_323), .B1(n_530), .B2(n_531), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_62), .A2(n_101), .B1(n_761), .B2(n_845), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_63), .A2(n_121), .B1(n_464), .B2(n_882), .Y(n_1051) );
AO222x2_ASAP7_75t_SL g517 ( .A1(n_64), .A2(n_124), .B1(n_171), .B2(n_518), .C1(n_519), .C2(n_520), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_65), .A2(n_141), .B1(n_419), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_66), .A2(n_295), .B1(n_485), .B2(n_842), .Y(n_841) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_68), .A2(n_203), .B1(n_400), .B2(n_411), .Y(n_410) );
XNOR2x1_ASAP7_75t_L g636 ( .A(n_70), .B(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_71), .A2(n_75), .B1(n_499), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_72), .A2(n_324), .B1(n_759), .B2(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_73), .A2(n_351), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_74), .A2(n_164), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI221x1_ASAP7_75t_L g652 ( .A1(n_76), .A2(n_85), .B1(n_509), .B2(n_653), .C(n_654), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_77), .A2(n_282), .B1(n_487), .B2(n_488), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g1002 ( .A1(n_79), .A2(n_335), .B1(n_485), .B2(n_842), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_80), .A2(n_129), .B1(n_593), .B2(n_594), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_81), .A2(n_168), .B1(n_421), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_82), .A2(n_331), .B1(n_499), .B2(n_534), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_83), .A2(n_202), .B1(n_671), .B2(n_738), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_84), .A2(n_266), .B1(n_445), .B2(n_566), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g1044 ( .A(n_87), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_88), .A2(n_253), .B1(n_645), .B2(n_758), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_89), .A2(n_278), .B1(n_499), .B2(n_585), .Y(n_584) );
AO22x1_ASAP7_75t_L g412 ( .A1(n_90), .A2(n_255), .B1(n_413), .B2(n_419), .Y(n_412) );
INVx1_ASAP7_75t_L g658 ( .A(n_91), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_92), .A2(n_380), .B1(n_506), .B2(n_507), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_93), .A2(n_263), .B1(n_534), .B2(n_566), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g857 ( .A1(n_94), .A2(n_300), .B1(n_421), .B2(n_690), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_95), .B(n_610), .Y(n_998) );
INVx1_ASAP7_75t_L g666 ( .A(n_97), .Y(n_666) );
INVx1_ASAP7_75t_L g643 ( .A(n_99), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_102), .A2(n_313), .B1(n_525), .B2(n_526), .Y(n_713) );
AO22x2_ASAP7_75t_L g1039 ( .A1(n_103), .A2(n_1040), .B1(n_1056), .B2(n_1057), .Y(n_1039) );
INVx1_ASAP7_75t_L g1057 ( .A(n_103), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_103), .A2(n_1062), .B1(n_1065), .B2(n_1066), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_105), .A2(n_245), .B1(n_533), .B2(n_537), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_106), .A2(n_334), .B1(n_523), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_107), .A2(n_356), .B1(n_414), .B2(n_491), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_108), .A2(n_368), .B1(n_413), .B2(n_948), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_111), .A2(n_146), .B1(n_473), .B2(n_485), .Y(n_484) );
OAI22x1_ASAP7_75t_L g956 ( .A1(n_112), .A2(n_957), .B1(n_958), .B2(n_969), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_112), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_113), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_114), .A2(n_256), .B1(n_645), .B2(n_758), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_115), .A2(n_272), .B1(n_602), .B2(n_837), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_118), .A2(n_190), .B1(n_653), .B2(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_120), .A2(n_329), .B1(n_451), .B2(n_869), .Y(n_1006) );
AO22x2_ASAP7_75t_L g407 ( .A1(n_122), .A2(n_286), .B1(n_400), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_123), .A2(n_231), .B1(n_487), .B2(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_125), .A2(n_208), .B1(n_696), .B2(n_848), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_126), .A2(n_337), .B1(n_759), .B2(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_127), .A2(n_153), .B1(n_433), .B2(n_509), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_130), .A2(n_348), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_131), .A2(n_184), .B1(n_519), .B2(n_520), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_132), .A2(n_271), .B1(n_594), .B2(n_775), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_133), .A2(n_154), .B1(n_612), .B2(n_863), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_134), .A2(n_161), .B1(n_817), .B2(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_135), .A2(n_175), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_136), .A2(n_346), .B1(n_455), .B2(n_458), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_137), .A2(n_152), .B1(n_758), .B2(n_759), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_139), .A2(n_238), .B1(n_440), .B2(n_443), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_140), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g788 ( .A(n_142), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_143), .A2(n_217), .B1(n_525), .B2(n_559), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_144), .A2(n_1056), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g1063 ( .A(n_144), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_145), .A2(n_156), .B1(n_413), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_148), .A2(n_315), .B1(n_519), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_149), .A2(n_298), .B1(n_507), .B2(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_150), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_151), .A2(n_363), .B1(n_473), .B2(n_814), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_155), .A2(n_316), .B1(n_506), .B2(n_507), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_157), .Y(n_634) );
AO22x1_ASAP7_75t_L g733 ( .A1(n_158), .A2(n_226), .B1(n_421), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_159), .A2(n_180), .B1(n_836), .B2(n_837), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_160), .B(n_572), .Y(n_797) );
INVx1_ASAP7_75t_L g1029 ( .A(n_162), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_163), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_165), .A2(n_267), .B1(n_593), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_166), .A2(n_232), .B1(n_530), .B2(n_531), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_167), .A2(n_187), .B1(n_533), .B2(n_537), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_169), .A2(n_355), .B1(n_525), .B2(n_526), .Y(n_576) );
OA22x2_ASAP7_75t_L g481 ( .A1(n_170), .A2(n_482), .B1(n_511), .B2(n_512), .Y(n_481) );
INVx1_ASAP7_75t_L g511 ( .A(n_170), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_172), .A2(n_292), .B1(n_693), .B2(n_826), .Y(n_1054) );
INVx1_ASAP7_75t_L g642 ( .A(n_173), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_174), .A2(n_361), .B1(n_485), .B2(n_860), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_176), .A2(n_209), .B1(n_674), .B2(n_675), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_177), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_178), .A2(n_247), .B1(n_500), .B2(n_825), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_179), .A2(n_220), .B1(n_641), .B2(n_822), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_181), .A2(n_287), .B1(n_755), .B2(n_888), .Y(n_975) );
XNOR2x1_ASAP7_75t_L g995 ( .A(n_182), .B(n_996), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_183), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_185), .A2(n_349), .B1(n_499), .B2(n_534), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_186), .B(n_419), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_188), .A2(n_249), .B1(n_433), .B2(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_191), .B(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_192), .A2(n_237), .B1(n_761), .B2(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_193), .A2(n_251), .B1(n_585), .B2(n_758), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_196), .A2(n_330), .B1(n_497), .B2(n_500), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_197), .A2(n_290), .B1(n_490), .B2(n_491), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_199), .A2(n_370), .B1(n_530), .B2(n_531), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_200), .A2(n_273), .B1(n_445), .B2(n_499), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_201), .A2(n_246), .B1(n_641), .B2(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g1026 ( .A(n_203), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_204), .A2(n_269), .B1(n_487), .B2(n_523), .Y(n_714) );
INVx1_ASAP7_75t_L g648 ( .A(n_205), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_206), .A2(n_264), .B1(n_753), .B2(n_755), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_207), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_212), .A2(n_372), .B1(n_749), .B2(n_751), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_213), .A2(n_306), .B1(n_531), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_214), .A2(n_373), .B1(n_751), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_215), .A2(n_365), .B1(n_451), .B2(n_776), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_216), .A2(n_248), .B1(n_506), .B2(n_507), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_218), .A2(n_377), .B1(n_599), .B2(n_828), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_219), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_221), .A2(n_374), .B1(n_519), .B2(n_520), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_222), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_224), .A2(n_243), .B1(n_421), .B2(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_225), .A2(n_382), .B1(n_593), .B2(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g1035 ( .A(n_227), .Y(n_1035) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_228), .B(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_229), .A2(n_240), .B1(n_455), .B2(n_458), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_230), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_233), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_234), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_236), .A2(n_257), .B1(n_499), .B2(n_534), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_239), .A2(n_321), .B1(n_427), .B2(n_433), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_241), .A2(n_307), .B1(n_506), .B2(n_507), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_244), .A2(n_332), .B1(n_487), .B2(n_523), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_250), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_261), .A2(n_268), .B1(n_451), .B2(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g647 ( .A(n_270), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_275), .A2(n_322), .B1(n_784), .B2(n_840), .Y(n_839) );
OA22x2_ASAP7_75t_L g970 ( .A1(n_276), .A2(n_971), .B1(n_972), .B2(n_986), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_276), .Y(n_971) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_276), .A2(n_972), .B(n_990), .Y(n_989) );
XNOR2xp5_ASAP7_75t_L g705 ( .A(n_277), .B(n_706), .Y(n_705) );
AOI22x1_ASAP7_75t_L g514 ( .A1(n_279), .A2(n_515), .B1(n_539), .B2(n_540), .Y(n_514) );
INVx1_ASAP7_75t_L g540 ( .A(n_279), .Y(n_540) );
XNOR2x1_ASAP7_75t_L g875 ( .A(n_281), .B(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_285), .B(n_937), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_286), .B(n_1025), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_289), .A2(n_312), .B1(n_534), .B2(n_566), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_291), .B(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_293), .A2(n_366), .B1(n_525), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_297), .A2(n_339), .B1(n_651), .B2(n_825), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_302), .A2(n_375), .B1(n_749), .B2(n_751), .Y(n_966) );
AND2x2_ASAP7_75t_L g730 ( .A(n_303), .B(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_304), .A2(n_319), .B1(n_451), .B2(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g400 ( .A(n_305), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_308), .Y(n_926) );
INVx1_ASAP7_75t_L g659 ( .A(n_309), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_310), .A2(n_326), .B1(n_462), .B2(n_464), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_314), .A2(n_325), .B1(n_421), .B2(n_879), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_318), .A2(n_367), .B1(n_738), .B2(n_884), .Y(n_981) );
INVx1_ASAP7_75t_L g725 ( .A(n_320), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_327), .Y(n_930) );
AND2x2_ASAP7_75t_L g392 ( .A(n_328), .B(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_333), .A2(n_381), .B1(n_470), .B2(n_603), .Y(n_687) );
INVx1_ASAP7_75t_L g668 ( .A(n_336), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_338), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_340), .A2(n_345), .B1(n_942), .B2(n_943), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_341), .A2(n_344), .B1(n_448), .B2(n_451), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_350), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_352), .B(n_555), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_354), .A2(n_362), .B1(n_674), .B2(n_939), .Y(n_938) );
OAI22x1_ASAP7_75t_L g682 ( .A1(n_357), .A2(n_683), .B1(n_684), .B2(n_703), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_357), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_358), .B(n_610), .Y(n_838) );
INVx1_ASAP7_75t_L g1021 ( .A(n_359), .Y(n_1021) );
NAND2xp5_ASAP7_75t_SL g1036 ( .A(n_359), .B(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1022 ( .A(n_360), .Y(n_1022) );
AND2x2_ASAP7_75t_R g1065 ( .A(n_360), .B(n_1021), .Y(n_1065) );
INVxp67_ASAP7_75t_L g1037 ( .A(n_364), .Y(n_1037) );
XNOR2xp5_ASAP7_75t_L g587 ( .A(n_369), .B(n_588), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_371), .Y(n_745) );
INVx1_ASAP7_75t_L g663 ( .A(n_378), .Y(n_663) );
XOR2x2_ASAP7_75t_L g805 ( .A(n_379), .B(n_806), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_1028), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_764), .B1(n_1016), .B2(n_1017), .C(n_1018), .Y(n_384) );
INVxp67_ASAP7_75t_L g1017 ( .A(n_385), .Y(n_1017) );
XNOR2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_678), .Y(n_385) );
XNOR2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_545), .Y(n_386) );
AO22x2_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_480), .B1(n_543), .B2(n_544), .Y(n_387) );
INVx1_ASAP7_75t_L g543 ( .A(n_388), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_389), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_460), .Y(n_390) );
NOR3xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_412), .C(n_425), .Y(n_391) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_SL g494 ( .A(n_395), .Y(n_494) );
INVx4_ASAP7_75t_SL g555 ( .A(n_395), .Y(n_555) );
INVx4_ASAP7_75t_SL g572 ( .A(n_395), .Y(n_572) );
BUFx2_ASAP7_75t_L g732 ( .A(n_395), .Y(n_732) );
INVx3_ASAP7_75t_L g937 ( .A(n_395), .Y(n_937) );
INVx6_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_405), .Y(n_396) );
AND2x4_ASAP7_75t_L g466 ( .A(n_397), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g474 ( .A(n_397), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g488 ( .A(n_397), .B(n_467), .Y(n_488) );
AND2x4_ASAP7_75t_L g518 ( .A(n_397), .B(n_405), .Y(n_518) );
AND2x2_ASAP7_75t_L g523 ( .A(n_397), .B(n_467), .Y(n_523) );
AND2x2_ASAP7_75t_L g526 ( .A(n_397), .B(n_475), .Y(n_526) );
AND2x2_ASAP7_75t_L g559 ( .A(n_397), .B(n_475), .Y(n_559) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_403), .Y(n_397) );
AND2x2_ASAP7_75t_L g417 ( .A(n_398), .B(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
INVx2_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
OAI22x1_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_400), .Y(n_404) );
INVx2_ASAP7_75t_L g408 ( .A(n_400), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_400), .Y(n_411) );
INVx2_ASAP7_75t_L g418 ( .A(n_403), .Y(n_418) );
AND2x2_ASAP7_75t_L g431 ( .A(n_403), .B(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
AND2x2_ASAP7_75t_L g430 ( .A(n_405), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g442 ( .A(n_405), .B(n_436), .Y(n_442) );
AND2x4_ASAP7_75t_L g457 ( .A(n_405), .B(n_417), .Y(n_457) );
AND2x6_ASAP7_75t_L g499 ( .A(n_405), .B(n_431), .Y(n_499) );
AND2x2_ASAP7_75t_L g506 ( .A(n_405), .B(n_417), .Y(n_506) );
AND2x2_ASAP7_75t_L g533 ( .A(n_405), .B(n_436), .Y(n_533) );
AND2x2_ASAP7_75t_L g564 ( .A(n_405), .B(n_417), .Y(n_564) );
AND2x4_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g416 ( .A(n_407), .B(n_409), .Y(n_416) );
AND2x2_ASAP7_75t_L g423 ( .A(n_407), .B(n_410), .Y(n_423) );
INVx1_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
INVxp67_ASAP7_75t_L g467 ( .A(n_409), .Y(n_467) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g437 ( .A(n_410), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g905 ( .A(n_413), .Y(n_905) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
INVx2_ASAP7_75t_L g608 ( .A(n_415), .Y(n_608) );
BUFx5_ASAP7_75t_L g690 ( .A(n_415), .Y(n_690) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND2x4_ASAP7_75t_L g446 ( .A(n_416), .B(n_436), .Y(n_446) );
AND2x4_ASAP7_75t_L g463 ( .A(n_416), .B(n_431), .Y(n_463) );
AND2x2_ASAP7_75t_L g487 ( .A(n_416), .B(n_431), .Y(n_487) );
AND2x4_ASAP7_75t_L g519 ( .A(n_416), .B(n_417), .Y(n_519) );
AND2x2_ASAP7_75t_L g537 ( .A(n_416), .B(n_436), .Y(n_537) );
AND2x2_ASAP7_75t_L g625 ( .A(n_416), .B(n_431), .Y(n_625) );
AND2x2_ASAP7_75t_L g471 ( .A(n_417), .B(n_437), .Y(n_471) );
AND2x4_ASAP7_75t_L g525 ( .A(n_417), .B(n_437), .Y(n_525) );
AND2x4_ASAP7_75t_L g436 ( .A(n_418), .B(n_432), .Y(n_436) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI222xp33_ASAP7_75t_L g662 ( .A1(n_420), .A2(n_663), .B1(n_664), .B2(n_666), .C1(n_667), .C2(n_668), .Y(n_662) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g948 ( .A(n_421), .Y(n_948) );
BUFx12f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g492 ( .A(n_422), .Y(n_492) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AND2x4_ASAP7_75t_L g452 ( .A(n_423), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g459 ( .A(n_423), .B(n_436), .Y(n_459) );
AND2x4_ASAP7_75t_L g507 ( .A(n_423), .B(n_436), .Y(n_507) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_423), .B(n_424), .Y(n_520) );
AND2x4_ASAP7_75t_L g531 ( .A(n_423), .B(n_453), .Y(n_531) );
AND2x2_ASAP7_75t_SL g574 ( .A(n_423), .B(n_424), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_439), .C(n_447), .D(n_454), .Y(n_425) );
INVx1_ASAP7_75t_L g915 ( .A(n_427), .Y(n_915) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g695 ( .A(n_429), .Y(n_695) );
INVx2_ASAP7_75t_SL g758 ( .A(n_429), .Y(n_758) );
INVx3_ASAP7_75t_L g888 ( .A(n_429), .Y(n_888) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g597 ( .A(n_430), .Y(n_597) );
BUFx2_ASAP7_75t_L g641 ( .A(n_430), .Y(n_641) );
AND2x2_ASAP7_75t_L g450 ( .A(n_431), .B(n_437), .Y(n_450) );
AND2x2_ASAP7_75t_SL g530 ( .A(n_431), .B(n_437), .Y(n_530) );
AND2x2_ASAP7_75t_L g800 ( .A(n_431), .B(n_437), .Y(n_800) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g510 ( .A(n_434), .Y(n_510) );
INVx2_ASAP7_75t_L g645 ( .A(n_434), .Y(n_645) );
INVx1_ASAP7_75t_SL g696 ( .A(n_434), .Y(n_696) );
INVx2_ASAP7_75t_L g755 ( .A(n_434), .Y(n_755) );
INVx2_ASAP7_75t_L g773 ( .A(n_434), .Y(n_773) );
INVx2_ASAP7_75t_L g822 ( .A(n_434), .Y(n_822) );
INVx2_ASAP7_75t_SL g873 ( .A(n_434), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_434), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_913) );
INVx8_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AND2x6_ASAP7_75t_L g534 ( .A(n_436), .B(n_437), .Y(n_534) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_438), .Y(n_476) );
INVx2_ASAP7_75t_L g754 ( .A(n_440), .Y(n_754) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_440), .Y(n_848) );
INVx4_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_SL g509 ( .A(n_441), .Y(n_509) );
INVx3_ASAP7_75t_L g566 ( .A(n_441), .Y(n_566) );
INVx2_ASAP7_75t_SL g693 ( .A(n_441), .Y(n_693) );
INVx2_ASAP7_75t_L g778 ( .A(n_441), .Y(n_778) );
INVx2_ASAP7_75t_SL g828 ( .A(n_441), .Y(n_828) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_444), .A2(n_923), .B1(n_924), .B2(n_926), .Y(n_922) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_445), .Y(n_759) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g501 ( .A(n_446), .Y(n_501) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_446), .Y(n_599) );
BUFx3_ASAP7_75t_L g651 ( .A(n_446), .Y(n_651) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g504 ( .A(n_450), .Y(n_504) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_450), .Y(n_593) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g594 ( .A(n_452), .Y(n_594) );
INVx5_ASAP7_75t_SL g660 ( .A(n_452), .Y(n_660) );
BUFx3_ASAP7_75t_L g943 ( .A(n_452), .Y(n_943) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_456), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_646) );
INVx3_ASAP7_75t_L g698 ( .A(n_456), .Y(n_698) );
INVx2_ASAP7_75t_L g761 ( .A(n_456), .Y(n_761) );
INVx1_ASAP7_75t_SL g780 ( .A(n_456), .Y(n_780) );
INVx2_ASAP7_75t_L g867 ( .A(n_456), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_456), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_918) );
INVx6_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g825 ( .A(n_457), .Y(n_825) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_SL g653 ( .A(n_459), .Y(n_653) );
INVx2_ASAP7_75t_L g700 ( .A(n_459), .Y(n_700) );
BUFx2_ASAP7_75t_SL g845 ( .A(n_459), .Y(n_845) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_468), .Y(n_460) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_463), .Y(n_612) );
BUFx2_ASAP7_75t_L g816 ( .A(n_463), .Y(n_816) );
BUFx3_ASAP7_75t_L g882 ( .A(n_463), .Y(n_882) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g613 ( .A(n_465), .Y(n_613) );
INVx2_ASAP7_75t_L g675 ( .A(n_465), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_465), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_742) );
INVx2_ASAP7_75t_L g817 ( .A(n_465), .Y(n_817) );
INVx2_ASAP7_75t_L g837 ( .A(n_465), .Y(n_837) );
INVx2_ASAP7_75t_L g863 ( .A(n_465), .Y(n_863) );
INVx6_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_471), .Y(n_485) );
INVx3_ASAP7_75t_L g739 ( .A(n_471), .Y(n_739) );
BUFx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g604 ( .A(n_474), .Y(n_604) );
INVx1_ASAP7_75t_L g672 ( .A(n_474), .Y(n_672) );
BUFx4f_ASAP7_75t_L g860 ( .A(n_474), .Y(n_860) );
BUFx3_ASAP7_75t_L g884 ( .A(n_474), .Y(n_884) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g544 ( .A(n_480), .Y(n_544) );
AOI22x1_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_513), .B1(n_541), .B2(n_542), .Y(n_480) );
INVx2_ASAP7_75t_L g542 ( .A(n_481), .Y(n_542) );
INVx1_ASAP7_75t_L g512 ( .A(n_482), .Y(n_512) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .C(n_489), .D(n_493), .Y(n_483) );
BUFx6f_ASAP7_75t_SL g602 ( .A(n_485), .Y(n_602) );
BUFx6f_ASAP7_75t_SL g840 ( .A(n_490), .Y(n_840) );
INVx1_ASAP7_75t_L g1001 ( .A(n_490), .Y(n_1001) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g785 ( .A(n_492), .Y(n_785) );
INVx2_ASAP7_75t_L g880 ( .A(n_492), .Y(n_880) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_494), .Y(n_665) );
INVx2_ASAP7_75t_L g1043 ( .A(n_494), .Y(n_1043) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .C(n_505), .D(n_508), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_500), .Y(n_950) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g585 ( .A(n_501), .Y(n_585) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g657 ( .A(n_504), .Y(n_657) );
INVx1_ASAP7_75t_L g776 ( .A(n_504), .Y(n_776) );
INVx2_ASAP7_75t_SL g541 ( .A(n_513), .Y(n_541) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AO22x2_ASAP7_75t_L g617 ( .A1(n_514), .A2(n_618), .B1(n_619), .B2(n_635), .Y(n_617) );
INVx1_ASAP7_75t_L g635 ( .A(n_514), .Y(n_635) );
INVx1_ASAP7_75t_L g539 ( .A(n_515), .Y(n_539) );
NAND2x1_ASAP7_75t_SL g515 ( .A(n_516), .B(n_527), .Y(n_515) );
NOR2xp67_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVx2_ASAP7_75t_SL g709 ( .A(n_518), .Y(n_709) );
BUFx2_ASAP7_75t_L g983 ( .A(n_518), .Y(n_983) );
INVx1_ASAP7_75t_SL g985 ( .A(n_519), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_535), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_615), .B2(n_677), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OA22x2_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_587), .B2(n_614), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
XNOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_567), .Y(n_549) );
XNOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_560), .Y(n_552) );
NAND4xp25_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .C(n_557), .D(n_558), .Y(n_553) );
INVx1_ASAP7_75t_SL g809 ( .A(n_555), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .D(n_565), .Y(n_560) );
XOR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_586), .Y(n_567) );
NAND2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_578), .Y(n_568) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
BUFx2_ASAP7_75t_L g610 ( .A(n_572), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx2_ASAP7_75t_SL g614 ( .A(n_587), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g588 ( .A(n_589), .B(n_600), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .C(n_595), .D(n_596), .Y(n_589) );
INVx1_ASAP7_75t_L g911 ( .A(n_592), .Y(n_911) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND4xp25_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .C(n_609), .D(n_611), .Y(n_600) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g741 ( .A(n_604), .Y(n_741) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g667 ( .A(n_607), .Y(n_667) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g734 ( .A(n_608), .Y(n_734) );
INVx2_ASAP7_75t_L g879 ( .A(n_608), .Y(n_879) );
BUFx2_ASAP7_75t_L g674 ( .A(n_612), .Y(n_674) );
INVx1_ASAP7_75t_L g744 ( .A(n_612), .Y(n_744) );
BUFx2_ASAP7_75t_L g836 ( .A(n_612), .Y(n_836) );
BUFx4f_ASAP7_75t_SL g862 ( .A(n_612), .Y(n_862) );
INVx2_ASAP7_75t_L g677 ( .A(n_615), .Y(n_677) );
OA22x2_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_636), .B2(n_676), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
XOR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_634), .Y(n_619) );
NAND2x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_627), .Y(n_620) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g676 ( .A(n_636), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_652), .C(n_661), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_646), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_639) );
INVx2_ASAP7_75t_L g772 ( .A(n_640), .Y(n_772) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g921 ( .A(n_653), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g750 ( .A(n_657), .Y(n_750) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_657), .Y(n_869) );
INVx2_ASAP7_75t_L g702 ( .A(n_660), .Y(n_702) );
INVx2_ASAP7_75t_L g751 ( .A(n_660), .Y(n_751) );
INVx2_ASAP7_75t_L g890 ( .A(n_660), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_660), .A2(n_910), .B1(n_911), .B2(n_912), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_669), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_664), .A2(n_904), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_903) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_722), .B1(n_723), .B2(n_763), .Y(n_680) );
INVx2_ASAP7_75t_L g763 ( .A(n_681), .Y(n_763) );
XNOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_704), .Y(n_681) );
INVx2_ASAP7_75t_L g703 ( .A(n_684), .Y(n_703) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_691), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .C(n_688), .D(n_689), .Y(n_685) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .C(n_697), .D(n_701), .Y(n_691) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g826 ( .A(n_700), .Y(n_826) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_707), .B(n_715), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_710), .B(n_711), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_762), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_725), .B(n_728), .Y(n_762) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_746), .Y(n_728) );
NOR4xp75_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .C(n_735), .D(n_742), .Y(n_729) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_735) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx4_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g814 ( .A(n_739), .Y(n_814) );
INVx3_ASAP7_75t_L g842 ( .A(n_741), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_756), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g942 ( .A(n_750), .Y(n_942) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g1016 ( .A(n_764), .Y(n_1016) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_954), .B1(n_1014), .B2(n_1015), .Y(n_764) );
INVx1_ASAP7_75t_L g1015 ( .A(n_765), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_830), .B1(n_952), .B2(n_953), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
BUFx2_ASAP7_75t_L g952 ( .A(n_767), .Y(n_952) );
OA22x2_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_789), .B1(n_790), .B2(n_829), .Y(n_767) );
INVx1_ASAP7_75t_L g829 ( .A(n_768), .Y(n_829) );
XOR2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_788), .Y(n_768) );
NOR2x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_781), .Y(n_769) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_774), .C(n_777), .D(n_779), .Y(n_770) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .C(n_786), .D(n_787), .Y(n_781) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
XNOR2x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_805), .Y(n_790) );
INVx2_ASAP7_75t_L g1010 ( .A(n_791), .Y(n_1010) );
XNOR2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_804), .Y(n_791) );
NOR2x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_798), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .C(n_796), .D(n_797), .Y(n_793) );
NAND4xp25_ASAP7_75t_L g798 ( .A(n_799), .B(n_801), .C(n_802), .D(n_803), .Y(n_798) );
NAND2x1_ASAP7_75t_L g806 ( .A(n_807), .B(n_818), .Y(n_806) );
NOR2x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .Y(n_807) );
OAI21xp5_ASAP7_75t_SL g808 ( .A1(n_809), .A2(n_810), .B(n_811), .Y(n_808) );
OAI21xp33_ASAP7_75t_L g855 ( .A1(n_809), .A2(n_856), .B(n_857), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_823), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_827), .Y(n_823) );
BUFx2_ASAP7_75t_L g925 ( .A(n_828), .Y(n_925) );
INVx1_ASAP7_75t_L g953 ( .A(n_830), .Y(n_953) );
XNOR2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_897), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_850), .B1(n_851), .B2(n_896), .Y(n_831) );
INVx5_ASAP7_75t_L g896 ( .A(n_832), .Y(n_896) );
NOR2x1_ASAP7_75t_L g833 ( .A(n_834), .B(n_843), .Y(n_833) );
NAND4xp25_ASAP7_75t_L g834 ( .A(n_835), .B(n_838), .C(n_839), .D(n_841), .Y(n_834) );
NAND4xp25_ASAP7_75t_L g843 ( .A(n_844), .B(n_846), .C(n_847), .D(n_849), .Y(n_843) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_874), .B1(n_875), .B2(n_893), .Y(n_851) );
INVx1_ASAP7_75t_SL g894 ( .A(n_853), .Y(n_894) );
AND2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_864), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_858), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_861), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_870), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVx1_ASAP7_75t_SL g874 ( .A(n_875), .Y(n_874) );
OR2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_886), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_878), .B(n_881), .C(n_883), .D(n_885), .Y(n_877) );
BUFx6f_ASAP7_75t_SL g939 ( .A(n_884), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g886 ( .A(n_887), .B(n_889), .C(n_891), .D(n_892), .Y(n_886) );
OAI22xp5_ASAP7_75t_SL g897 ( .A1(n_898), .A2(n_899), .B1(n_931), .B2(n_951), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
XNOR2x1_ASAP7_75t_L g900 ( .A(n_901), .B(n_930), .Y(n_900) );
NAND4xp75_ASAP7_75t_L g901 ( .A(n_902), .B(n_908), .C(n_917), .D(n_927), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2x1_ASAP7_75t_L g908 ( .A(n_909), .B(n_913), .Y(n_908) );
NOR2x1_ASAP7_75t_L g917 ( .A(n_918), .B(n_922), .Y(n_917) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AND2x2_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
INVx1_ASAP7_75t_L g951 ( .A(n_931), .Y(n_951) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
XNOR2xp5_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
NOR2x1_ASAP7_75t_L g934 ( .A(n_935), .B(n_944), .Y(n_934) );
NAND4xp25_ASAP7_75t_L g935 ( .A(n_936), .B(n_938), .C(n_940), .D(n_941), .Y(n_935) );
NAND4xp25_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .C(n_947), .D(n_949), .Y(n_944) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_954), .Y(n_1014) );
AO22x2_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_992), .B1(n_1012), .B2(n_1013), .Y(n_954) );
INVx2_ASAP7_75t_SL g1012 ( .A(n_955), .Y(n_1012) );
OA22x2_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_970), .B1(n_987), .B2(n_988), .Y(n_955) );
INVx1_ASAP7_75t_SL g987 ( .A(n_956), .Y(n_987) );
INVx2_ASAP7_75t_SL g969 ( .A(n_958), .Y(n_969) );
OR2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_964), .Y(n_958) );
NAND4xp25_ASAP7_75t_SL g959 ( .A(n_960), .B(n_961), .C(n_962), .D(n_963), .Y(n_959) );
NAND4xp25_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .C(n_967), .D(n_968), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_970), .A2(n_988), .B1(n_995), .B2(n_1009), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_971), .Y(n_991) );
INVx1_ASAP7_75t_L g986 ( .A(n_972), .Y(n_986) );
NOR2x1_ASAP7_75t_SL g990 ( .A(n_972), .B(n_991), .Y(n_990) );
NAND4xp75_ASAP7_75t_L g972 ( .A(n_973), .B(n_976), .C(n_979), .D(n_982), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
AND2x2_ASAP7_75t_L g976 ( .A(n_977), .B(n_978), .Y(n_976) );
AND2x2_ASAP7_75t_L g979 ( .A(n_980), .B(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx3_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx4_ASAP7_75t_L g1013 ( .A(n_992), .Y(n_1013) );
OA22x2_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_994), .B1(n_1010), .B2(n_1011), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_SL g1009 ( .A(n_995), .Y(n_1009) );
OR2x2_ASAP7_75t_L g996 ( .A(n_997), .B(n_1004), .Y(n_996) );
NAND4xp25_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .C(n_1002), .D(n_1003), .Y(n_997) );
INVx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
NAND4xp25_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .C(n_1007), .D(n_1008), .Y(n_1004) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1010), .Y(n_1011) );
INVx3_ASAP7_75t_SL g1018 ( .A(n_1019), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1023), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1020), .B(n_1024), .Y(n_1060) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1022), .Y(n_1020) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1022), .Y(n_1032) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
OAI221xp5_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1030), .B1(n_1038), .B2(n_1058), .C(n_1061), .Y(n_1028) );
INVxp67_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NOR2x1_ASAP7_75t_R g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_1032), .B(n_1034), .Y(n_1067) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
INVx3_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx2_ASAP7_75t_SL g1056 ( .A(n_1040), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_1040), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1049), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1046), .Y(n_1041) );
OAI21xp33_ASAP7_75t_SL g1042 ( .A1(n_1043), .A2(n_1044), .B(n_1045), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .Y(n_1046) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1053), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_1059), .Y(n_1058) );
CKINVDCx6p67_ASAP7_75t_R g1059 ( .A(n_1060), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g1066 ( .A(n_1067), .Y(n_1066) );
endmodule