module fake_jpeg_26009_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_51),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_64),
.B1(n_62),
.B2(n_57),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_54),
.B1(n_63),
.B2(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_44),
.B1(n_47),
.B2(n_55),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_63),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_98),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_58),
.B1(n_49),
.B2(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_100),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_97),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_58),
.B1(n_68),
.B2(n_66),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_103),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_65),
.B1(n_59),
.B2(n_56),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_67),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_46),
.C(n_45),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_114),
.B1(n_111),
.B2(n_105),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_1),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_99),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_2),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_69),
.B(n_4),
.C(n_5),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_106),
.B(n_107),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_120),
.B1(n_121),
.B2(n_6),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_13),
.C(n_14),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_123),
.Y(n_136)
);

NAND2x1_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_3),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_17),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_7),
.B(n_8),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_134),
.C(n_135),
.Y(n_138)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_18),
.C(n_21),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_141),
.C(n_133),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_144),
.A2(n_145),
.B(n_142),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_128),
.B(n_143),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_136),
.B1(n_143),
.B2(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_24),
.B(n_27),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_28),
.B(n_30),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_31),
.C(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_35),
.Y(n_154)
);


endmodule