module fake_ariane_1343_n_5263 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_5263);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_5263;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_4824;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_1032;
wire n_1592;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_5053;
wire n_1243;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_3168;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_3645;
wire n_793;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_1141;
wire n_3457;
wire n_840;
wire n_2324;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_1581;
wire n_946;
wire n_3058;
wire n_757;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_998;
wire n_3592;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_1169;
wire n_789;
wire n_3181;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_3391;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_3508;
wire n_4129;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_779;
wire n_4790;
wire n_4173;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_3738;
wire n_894;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_3113;
wire n_2751;
wire n_4183;
wire n_918;
wire n_1968;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_4333;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_994;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_856;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_1410;
wire n_939;
wire n_2297;
wire n_4203;
wire n_1325;
wire n_1223;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_3763;
wire n_933;
wire n_3499;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_2361;
wire n_1752;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_2243;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_2731;
wire n_3703;
wire n_1246;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5050;
wire n_5240;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_2133;
wire n_2497;
wire n_879;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_4138;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_4435;
wire n_3248;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_4673;
wire n_2793;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_2039;
wire n_1285;
wire n_761;
wire n_733;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1982;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_2461;
wire n_1706;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_693;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_4794;
wire n_4843;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_824;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_1627;
wire n_2903;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_876;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_790;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_973;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_5133;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_123),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_293),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_532),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_682),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_10),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_376),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_209),
.Y(n_697)
);

CKINVDCx16_ASAP7_75t_R g698 ( 
.A(n_444),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_617),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_630),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_576),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_49),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_593),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_498),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_407),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_17),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_32),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_626),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_683),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_260),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_459),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_77),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_399),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_43),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_367),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_399),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_597),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_636),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_358),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_226),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_440),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_153),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_448),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_676),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_276),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_208),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_628),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_379),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_381),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_487),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_569),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_243),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_588),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_48),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_671),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_254),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_391),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_177),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_154),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_102),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_125),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_284),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_663),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_64),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_119),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_410),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_601),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_123),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_167),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_374),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_628),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_678),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_201),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_562),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_270),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_206),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_607),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_425),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_631),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_64),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_381),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_298),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_141),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_277),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_684),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_556),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_418),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_609),
.Y(n_768)
);

BUFx10_ASAP7_75t_L g769 ( 
.A(n_434),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_178),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_450),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_233),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_54),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_667),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_208),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_521),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_195),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_321),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_35),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_240),
.Y(n_780)
);

CKINVDCx14_ASAP7_75t_R g781 ( 
.A(n_75),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_484),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_636),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_315),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_640),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_418),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_434),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_676),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_152),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_175),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_566),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_669),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_607),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_278),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_624),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_495),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_533),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_602),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_198),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_468),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_655),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_129),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_137),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_446),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_353),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_532),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_190),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_350),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_593),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_248),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_207),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_344),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_652),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_110),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_111),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_196),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_351),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_58),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_533),
.Y(n_819)
);

CKINVDCx14_ASAP7_75t_R g820 ( 
.A(n_525),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_281),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_644),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_141),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_609),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_386),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_567),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_419),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_34),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_680),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_118),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_174),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_392),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_631),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_205),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_384),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_394),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_530),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_508),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_49),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_598),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_156),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_244),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_666),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_16),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_229),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_586),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_487),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_175),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_180),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_522),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_297),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_261),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_297),
.Y(n_853)
);

BUFx2_ASAP7_75t_R g854 ( 
.A(n_352),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_672),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_131),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_342),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_660),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_658),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_115),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_227),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_535),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_568),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_387),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_95),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_77),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_506),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_474),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_119),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_167),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_28),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_59),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_336),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_667),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_200),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_133),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_482),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_519),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_143),
.Y(n_879)
);

BUFx5_ASAP7_75t_L g880 ( 
.A(n_139),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_406),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_632),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_160),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_46),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_382),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_46),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_374),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_554),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_103),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_581),
.Y(n_890)
);

CKINVDCx14_ASAP7_75t_R g891 ( 
.A(n_461),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_150),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_600),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_665),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_476),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_117),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_238),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_480),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_400),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_637),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_46),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_119),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_25),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_588),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_207),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_630),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_540),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_242),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_511),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_681),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_419),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_657),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_540),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_488),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_162),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_323),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_320),
.Y(n_917)
);

BUFx10_ASAP7_75t_L g918 ( 
.A(n_264),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_489),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_627),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_354),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_306),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_250),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_572),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_15),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_329),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_601),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_263),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_131),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_651),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_420),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_324),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_504),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_666),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_379),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_453),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_585),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_307),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_679),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_237),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_571),
.Y(n_941)
);

BUFx10_ASAP7_75t_L g942 ( 
.A(n_157),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_106),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_18),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_462),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_403),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_543),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_606),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_689),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_424),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_595),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_499),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_612),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_366),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_362),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_523),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_629),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_437),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_442),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_91),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_138),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_519),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_660),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_165),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_1),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_309),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_171),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_59),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_521),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_445),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_679),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_411),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_352),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_433),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_404),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_314),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_659),
.Y(n_977)
);

CKINVDCx14_ASAP7_75t_R g978 ( 
.A(n_402),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_383),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_87),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_689),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_484),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_501),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_231),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_327),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_329),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_445),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_91),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_618),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_591),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_461),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_463),
.Y(n_992)
);

BUFx8_ASAP7_75t_SL g993 ( 
.A(n_499),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_181),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_506),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_555),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_130),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_439),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_310),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_559),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_110),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_199),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_514),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_145),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_71),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_556),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_327),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_261),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_26),
.Y(n_1009)
);

BUFx5_ASAP7_75t_L g1010 ( 
.A(n_197),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_554),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_291),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_342),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_318),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_31),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_51),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_210),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_312),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_511),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_677),
.Y(n_1020)
);

CKINVDCx12_ASAP7_75t_R g1021 ( 
.A(n_74),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_665),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_508),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_377),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_626),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_464),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_820),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_891),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_902),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_902),
.Y(n_1030)
);

CKINVDCx16_ASAP7_75t_R g1031 ( 
.A(n_781),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_978),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_880),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_758),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_965),
.B(n_0),
.Y(n_1035)
);

CKINVDCx16_ASAP7_75t_R g1036 ( 
.A(n_698),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_993),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1001),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_762),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_758),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_1005),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_880),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_845),
.Y(n_1043)
);

INVxp33_ASAP7_75t_L g1044 ( 
.A(n_700),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_845),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_910),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_778),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_880),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_838),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_910),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_882),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_935),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_761),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_935),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_940),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_940),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_764),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_766),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_767),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_949),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_880),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_949),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_719),
.B(n_0),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_880),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_695),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_768),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1009),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_854),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_707),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_740),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_748),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_760),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_771),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_701),
.B(n_0),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_773),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_774),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_814),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_1015),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_782),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_784),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_786),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_839),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_694),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_871),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_889),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_787),
.Y(n_1086)
);

CKINVDCx16_ASAP7_75t_R g1087 ( 
.A(n_769),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_943),
.Y(n_1088)
);

BUFx2_ASAP7_75t_SL g1089 ( 
.A(n_880),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_788),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_968),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_1021),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_988),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_703),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_869),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_869),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_789),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_791),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_872),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_872),
.Y(n_1100)
);

INVxp33_ASAP7_75t_L g1101 ( 
.A(n_859),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_792),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_717),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_880),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_884),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_884),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_880),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1010),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1010),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1010),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_718),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1010),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_793),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_694),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1010),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1010),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1010),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1010),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_794),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_704),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_721),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_730),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_722),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_723),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_694),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_795),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_797),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_799),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_801),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_803),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_777),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_868),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_724),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_804),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_805),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_870),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_694),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_725),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_731),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_769),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_806),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_732),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_694),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_807),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_808),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_737),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_738),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_810),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_739),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1000),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_811),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_746),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_749),
.Y(n_1153)
);

BUFx2_ASAP7_75t_SL g1154 ( 
.A(n_705),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_705),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_750),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_705),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_812),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_751),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_754),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_755),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_691),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_757),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_813),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_759),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_763),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_816),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_765),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_772),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_817),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_819),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_705),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_705),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_720),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_822),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_775),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_776),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_783),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_785),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_823),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_720),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_720),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_720),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_769),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_802),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_809),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_843),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_836),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_796),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_824),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_837),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_835),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_897),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_720),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_825),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_826),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_855),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_701),
.B(n_1),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_827),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_864),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_829),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_873),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_874),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_831),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_727),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_875),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_727),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_883),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_879),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_727),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_832),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_888),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_894),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_833),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_895),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_912),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_904),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_906),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_840),
.Y(n_1219)
);

NOR2xp67_ASAP7_75t_L g1220 ( 
.A(n_780),
.B(n_1),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_841),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_911),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_727),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_913),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_929),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_950),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_933),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_937),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_727),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_946),
.Y(n_1230)
);

CKINVDCx16_ASAP7_75t_R g1231 ( 
.A(n_843),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_947),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_952),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_843),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_955),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_957),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_842),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_967),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_961),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_971),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_790),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_780),
.B(n_2),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_979),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_996),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1003),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_790),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_790),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_790),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_975),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1004),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1006),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1007),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_983),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_846),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1026),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_790),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_800),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_691),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_702),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_800),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_848),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_850),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_821),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_821),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_851),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_834),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_852),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_834),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_853),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_990),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_856),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_857),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_861),
.Y(n_1273)
);

INVxp33_ASAP7_75t_L g1274 ( 
.A(n_861),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1018),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_878),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_798),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_878),
.Y(n_1278)
);

NOR2xp67_ASAP7_75t_L g1279 ( 
.A(n_863),
.B(n_2),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_887),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_887),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_858),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_798),
.Y(n_1283)
);

BUFx8_ASAP7_75t_SL g1284 ( 
.A(n_706),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_892),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_892),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_931),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_798),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_931),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_798),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_863),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_989),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_706),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_862),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_876),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_798),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_989),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_877),
.Y(n_1298)
);

CKINVDCx16_ASAP7_75t_R g1299 ( 
.A(n_917),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_712),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_964),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_964),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_964),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_964),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_964),
.Y(n_1305)
);

NOR2xp67_ASAP7_75t_L g1306 ( 
.A(n_711),
.B(n_2),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_973),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_973),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_692),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_973),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_973),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_973),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_992),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_992),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_992),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_992),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_992),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_881),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_712),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_779),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_885),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_917),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_890),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_714),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_917),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_815),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_818),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_828),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_714),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_918),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_893),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_898),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_830),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_844),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_860),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_918),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_899),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_752),
.B(n_3),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_900),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_886),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_905),
.Y(n_1341)
);

BUFx10_ASAP7_75t_L g1342 ( 
.A(n_734),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_896),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_918),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_735),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_901),
.Y(n_1346)
);

BUFx8_ASAP7_75t_SL g1347 ( 
.A(n_734),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_907),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_903),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_741),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_908),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_914),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_934),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_934),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_915),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_916),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_925),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_944),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_934),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_741),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_744),
.Y(n_1361)
);

NOR2xp67_ASAP7_75t_L g1362 ( 
.A(n_847),
.B(n_3),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_744),
.B(n_3),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_942),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_919),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_942),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_745),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_920),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_745),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_865),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_865),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_866),
.B(n_4),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_921),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_866),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_960),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_960),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_980),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_942),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_980),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_922),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_923),
.Y(n_1381)
);

NOR2xp67_ASAP7_75t_L g1382 ( 
.A(n_1016),
.B(n_4),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1016),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_924),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_977),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_693),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_926),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_927),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_693),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_770),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1120),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1121),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1123),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1284),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1309),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1124),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1065),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1347),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1037),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1320),
.B(n_928),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1133),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1037),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1138),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1111),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1139),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1142),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_R g1407 ( 
.A(n_1134),
.B(n_930),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1065),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1078),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1146),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1147),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1149),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1078),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1152),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1153),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1156),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1159),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_1108),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1226),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1160),
.Y(n_1420)
);

CKINVDCx16_ASAP7_75t_R g1421 ( 
.A(n_1031),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1253),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1161),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1326),
.B(n_932),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1163),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1135),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1165),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1166),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1094),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1168),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1141),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1169),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1144),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1094),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1145),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1148),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1053),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1345),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1176),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1177),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1178),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1179),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1027),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1185),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1027),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1330),
.B(n_1293),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1186),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1188),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1191),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1390),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1028),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1028),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1103),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1038),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1053),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1103),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_SL g1457 ( 
.A(n_1342),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1057),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1330),
.B(n_936),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1057),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1197),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1330),
.B(n_938),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1058),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1200),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1388),
.B(n_945),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1202),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1203),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1041),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1206),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1058),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1059),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1059),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1066),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1172),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1162),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1208),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1212),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1122),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1327),
.B(n_948),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1172),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1066),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1073),
.B(n_951),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1213),
.Y(n_1483)
);

BUFx2_ASAP7_75t_SL g1484 ( 
.A(n_1342),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1122),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1324),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1073),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1076),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1131),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1108),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1076),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1079),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1388),
.B(n_953),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1079),
.Y(n_1494)
);

CKINVDCx14_ASAP7_75t_R g1495 ( 
.A(n_1032),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1143),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1080),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1328),
.B(n_954),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1080),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1081),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1215),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1081),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1086),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1274),
.B(n_696),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1086),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1131),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1370),
.Y(n_1507)
);

INVxp33_ASAP7_75t_SL g1508 ( 
.A(n_1032),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1217),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1143),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1300),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1218),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1090),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1189),
.Y(n_1514)
);

INVxp33_ASAP7_75t_SL g1515 ( 
.A(n_1039),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1090),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1189),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1222),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1224),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1192),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1097),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1225),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1227),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1192),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1209),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1228),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1230),
.Y(n_1527)
);

CKINVDCx14_ASAP7_75t_R g1528 ( 
.A(n_1342),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1232),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1258),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1209),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1233),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1097),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1216),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1235),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1216),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_1087),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1098),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1098),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1322),
.B(n_956),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1236),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1083),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1172),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1172),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1239),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1102),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1240),
.Y(n_1547)
);

INVxp33_ASAP7_75t_SL g1548 ( 
.A(n_1039),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1047),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1102),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1243),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1113),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1379),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1244),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1210),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1157),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1245),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1083),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1250),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1113),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1119),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1251),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1252),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1255),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1238),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1132),
.B(n_849),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1069),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1119),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_L g1569 ( 
.A(n_1126),
.B(n_958),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1044),
.B(n_696),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1070),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1126),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1071),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1127),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1127),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1238),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1249),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1249),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1128),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1128),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1072),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1129),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1075),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1077),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1082),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1210),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1129),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1130),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1270),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1084),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1270),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1275),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1130),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1151),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1085),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1210),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1088),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1275),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1091),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1151),
.Y(n_1600)
);

INVxp33_ASAP7_75t_SL g1601 ( 
.A(n_1047),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1158),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1093),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1158),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1164),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1029),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1030),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1333),
.B(n_1334),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1107),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1210),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1109),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1335),
.B(n_1340),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1110),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1223),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1112),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1101),
.B(n_697),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1300),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1319),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1164),
.Y(n_1619)
);

CKINVDCx16_ASAP7_75t_R g1620 ( 
.A(n_1140),
.Y(n_1620)
);

BUFx2_ASAP7_75t_SL g1621 ( 
.A(n_1319),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1167),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1167),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1170),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1170),
.Y(n_1625)
);

NOR2xp67_ASAP7_75t_L g1626 ( 
.A(n_1171),
.B(n_697),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1049),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1116),
.Y(n_1628)
);

CKINVDCx16_ASAP7_75t_R g1629 ( 
.A(n_1231),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1049),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1117),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1329),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1118),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1171),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1154),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1329),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1034),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1223),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1175),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1040),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1043),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_1350),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1175),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1045),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1180),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1050),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1157),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1180),
.Y(n_1648)
);

INVxp33_ASAP7_75t_L g1649 ( 
.A(n_1092),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1052),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1190),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1054),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1350),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1055),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1056),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1060),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1183),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1190),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1051),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1223),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1195),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1136),
.B(n_909),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1195),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1062),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_1361),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1361),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1375),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1183),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1248),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1248),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1196),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1196),
.Y(n_1672)
);

CKINVDCx20_ASAP7_75t_R g1673 ( 
.A(n_1375),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1343),
.B(n_699),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_1036),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1083),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1199),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1346),
.B(n_699),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1290),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1349),
.B(n_708),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1357),
.B(n_708),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1290),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1199),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1234),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1291),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1344),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1292),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1297),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1322),
.B(n_1023),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1358),
.B(n_709),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1201),
.Y(n_1691)
);

CKINVDCx20_ASAP7_75t_R g1692 ( 
.A(n_1299),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1201),
.Y(n_1693)
);

INVxp33_ASAP7_75t_L g1694 ( 
.A(n_1322),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1204),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1336),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1446),
.B(n_1322),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1558),
.B(n_1325),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1674),
.A2(n_1063),
.B1(n_1385),
.B2(n_1187),
.Y(n_1699)
);

BUFx12f_ASAP7_75t_L g1700 ( 
.A(n_1394),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1685),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1504),
.B(n_1383),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1586),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1609),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1586),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1586),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1586),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1558),
.B(n_1325),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1570),
.B(n_1383),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1542),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1586),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1611),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1391),
.B(n_1325),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1617),
.A2(n_1068),
.B1(n_1051),
.B2(n_1035),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1450),
.B(n_1344),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1668),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1558),
.B(n_1325),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1613),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1676),
.B(n_1378),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1474),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1669),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1378),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1670),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1615),
.Y(n_1724)
);

INVx5_ASAP7_75t_L g1725 ( 
.A(n_1676),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1395),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1679),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1628),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1631),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1633),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1635),
.B(n_1378),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1687),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1474),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1480),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1480),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1608),
.B(n_1089),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1678),
.A2(n_1184),
.B1(n_1187),
.B2(n_1204),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1688),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1543),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1438),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1612),
.B(n_1353),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1606),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1543),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1542),
.B(n_1353),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1544),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1694),
.B(n_1360),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1544),
.A2(n_1042),
.B(n_1033),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1555),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1555),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1596),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1596),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1607),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1392),
.B(n_1393),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1610),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1675),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1459),
.B(n_1354),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1637),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1640),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1662),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1610),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1398),
.Y(n_1762)
);

AND2x2_ASAP7_75t_SL g1763 ( 
.A(n_1421),
.B(n_1198),
.Y(n_1763)
);

CKINVDCx6p67_ASAP7_75t_R g1764 ( 
.A(n_1457),
.Y(n_1764)
);

BUFx8_ASAP7_75t_L g1765 ( 
.A(n_1457),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1484),
.A2(n_1363),
.B1(n_1242),
.B2(n_1259),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1614),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1614),
.Y(n_1768)
);

AND2x2_ASAP7_75t_SL g1769 ( 
.A(n_1537),
.B(n_1354),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1457),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1426),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1638),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1462),
.B(n_1367),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1680),
.A2(n_1184),
.B1(n_1214),
.B2(n_1211),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1617),
.A2(n_1211),
.B1(n_1219),
.B2(n_1214),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1638),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1465),
.B(n_1369),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1660),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1641),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1660),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1496),
.B(n_1359),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1644),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1646),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1567),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1650),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1571),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1510),
.B(n_1359),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1616),
.B(n_1364),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1652),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1675),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1396),
.B(n_1364),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1654),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1655),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1656),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1664),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1573),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1581),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1583),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1468),
.Y(n_1799)
);

OAI22x1_ASAP7_75t_L g1800 ( 
.A1(n_1511),
.A2(n_1150),
.B1(n_1193),
.B2(n_1067),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1584),
.Y(n_1801)
);

OAI22x1_ASAP7_75t_R g1802 ( 
.A1(n_1618),
.A2(n_710),
.B1(n_713),
.B2(n_709),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1556),
.B(n_1647),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1401),
.B(n_1366),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1657),
.B(n_1366),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1403),
.B(n_1371),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1585),
.Y(n_1807)
);

OA21x2_ASAP7_75t_L g1808 ( 
.A1(n_1493),
.A2(n_1042),
.B(n_1033),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1590),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1540),
.B(n_1374),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1595),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1405),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1406),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1410),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1597),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1411),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1682),
.B(n_1418),
.Y(n_1817)
);

OA21x2_ASAP7_75t_L g1818 ( 
.A1(n_1689),
.A2(n_1061),
.B(n_1048),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_SL g1819 ( 
.A(n_1515),
.B(n_1219),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1599),
.B(n_1376),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1412),
.B(n_1377),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1681),
.A2(n_1237),
.B1(n_1254),
.B2(n_1221),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1490),
.B(n_1386),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1603),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1414),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1566),
.B(n_1221),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1415),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1416),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1417),
.A2(n_1061),
.B(n_1048),
.Y(n_1829)
);

OA21x2_ASAP7_75t_L g1830 ( 
.A1(n_1420),
.A2(n_1104),
.B(n_1064),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1423),
.B(n_1074),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1425),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1427),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1397),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1404),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1454),
.B(n_1237),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1428),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1400),
.B(n_1389),
.Y(n_1838)
);

AND2x6_ASAP7_75t_L g1839 ( 
.A(n_1430),
.B(n_1064),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1432),
.B(n_1220),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1424),
.B(n_1254),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1684),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1690),
.A2(n_1262),
.B1(n_1265),
.B2(n_1261),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1439),
.B(n_1279),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1440),
.Y(n_1845)
);

XNOR2x1_ASAP7_75t_L g1846 ( 
.A(n_1419),
.B(n_1261),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1479),
.B(n_1498),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1441),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1442),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1475),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1444),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1447),
.Y(n_1852)
);

OA21x2_ASAP7_75t_L g1853 ( 
.A1(n_1448),
.A2(n_1115),
.B(n_1104),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1449),
.A2(n_1115),
.B(n_1302),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1461),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1486),
.Y(n_1856)
);

OAI22x1_ASAP7_75t_R g1857 ( 
.A1(n_1618),
.A2(n_713),
.B1(n_715),
.B2(n_710),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1464),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1686),
.B(n_1262),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1466),
.A2(n_1305),
.B(n_1303),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1467),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1469),
.B(n_1265),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1476),
.B(n_1372),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1477),
.B(n_1267),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1483),
.B(n_1046),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1501),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1509),
.B(n_1267),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1512),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1433),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1435),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1518),
.B(n_1519),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1482),
.B(n_1569),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1522),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1523),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1526),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1527),
.B(n_1269),
.Y(n_1876)
);

INVx5_ASAP7_75t_L g1877 ( 
.A(n_1620),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1529),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1436),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1532),
.B(n_1535),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1541),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1545),
.B(n_1269),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1426),
.Y(n_1883)
);

INVx5_ASAP7_75t_L g1884 ( 
.A(n_1629),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1547),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1632),
.A2(n_1272),
.B1(n_1282),
.B2(n_1271),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1551),
.B(n_1046),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1422),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1507),
.B(n_1271),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1554),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1557),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1431),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1559),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1562),
.Y(n_1894)
);

INVx5_ASAP7_75t_L g1895 ( 
.A(n_1528),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1563),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1632),
.A2(n_1642),
.B1(n_1653),
.B2(n_1636),
.Y(n_1897)
);

INVx5_ASAP7_75t_L g1898 ( 
.A(n_1564),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1431),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1399),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1530),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1553),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1626),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1437),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1455),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1458),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1508),
.B(n_1272),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1508),
.B(n_1282),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1460),
.B(n_1294),
.Y(n_1909)
);

INVxp67_ASAP7_75t_L g1910 ( 
.A(n_1621),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1463),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1470),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1471),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1472),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1473),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1443),
.A2(n_1310),
.B(n_1307),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1481),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1549),
.B(n_1382),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1533),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1487),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1533),
.A2(n_1295),
.B1(n_1298),
.B2(n_1294),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1488),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1491),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1492),
.Y(n_1924)
);

INVx5_ASAP7_75t_L g1925 ( 
.A(n_1495),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1494),
.Y(n_1926)
);

OA21x2_ASAP7_75t_L g1927 ( 
.A1(n_1443),
.A2(n_1312),
.B(n_1311),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1604),
.A2(n_716),
.B1(n_726),
.B2(n_715),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1627),
.B(n_1306),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1497),
.Y(n_1930)
);

CKINVDCx8_ASAP7_75t_R g1931 ( 
.A(n_1402),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1630),
.B(n_1338),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1499),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1500),
.B(n_1295),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1502),
.B(n_1365),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1649),
.B(n_1095),
.Y(n_1936)
);

OA21x2_ASAP7_75t_L g1937 ( 
.A1(n_1445),
.A2(n_1315),
.B(n_1313),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1503),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1505),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1659),
.B(n_1362),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1513),
.Y(n_1941)
);

OA21x2_ASAP7_75t_L g1942 ( 
.A1(n_1445),
.A2(n_1317),
.B(n_1316),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1516),
.B(n_1298),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1397),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1604),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1521),
.B(n_1318),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1538),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1451),
.A2(n_1137),
.B(n_1125),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1539),
.B(n_1318),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1546),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1550),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1605),
.A2(n_1695),
.B1(n_1622),
.B2(n_1623),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1605),
.A2(n_726),
.B1(n_728),
.B2(n_716),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1552),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1560),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1561),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1568),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1572),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1574),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1575),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1579),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1580),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1582),
.Y(n_1963)
);

OA21x2_ASAP7_75t_L g1964 ( 
.A1(n_1451),
.A2(n_1137),
.B(n_1125),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1587),
.B(n_1321),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1588),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1636),
.A2(n_1323),
.B1(n_1331),
.B2(n_1321),
.Y(n_1967)
);

OA21x2_ASAP7_75t_L g1968 ( 
.A1(n_1452),
.A2(n_1173),
.B(n_1155),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1642),
.A2(n_1331),
.B1(n_1332),
.B2(n_1323),
.Y(n_1969)
);

OA21x2_ASAP7_75t_L g1970 ( 
.A1(n_1452),
.A2(n_1173),
.B(n_1155),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1593),
.B(n_1332),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1684),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1594),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1600),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1602),
.B(n_1337),
.Y(n_1975)
);

NAND2xp33_ASAP7_75t_L g1976 ( 
.A(n_1619),
.B(n_1337),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1515),
.A2(n_1246),
.B(n_1114),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1619),
.B(n_1339),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1634),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1645),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1648),
.Y(n_1981)
);

AND2x2_ASAP7_75t_SL g1982 ( 
.A(n_1548),
.B(n_1174),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1622),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1651),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1658),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1762),
.Y(n_1986)
);

OAI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1847),
.A2(n_1695),
.B1(n_1624),
.B2(n_1625),
.Y(n_1987)
);

OAI22xp33_ASAP7_75t_SL g1988 ( 
.A1(n_1766),
.A2(n_1624),
.B1(n_1625),
.B2(n_1623),
.Y(n_1988)
);

AO22x2_ASAP7_75t_L g1989 ( 
.A1(n_1846),
.A2(n_1665),
.B1(n_1666),
.B2(n_1653),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1841),
.A2(n_1643),
.B1(n_1639),
.B2(n_1661),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1715),
.B(n_1639),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1854),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1854),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1760),
.B(n_1643),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1841),
.A2(n_1671),
.B1(n_1672),
.B2(n_1663),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1741),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1726),
.B(n_1677),
.Y(n_1997)
);

OAI22xp33_ASAP7_75t_R g1998 ( 
.A1(n_1907),
.A2(n_941),
.B1(n_985),
.B2(n_939),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1854),
.Y(n_1999)
);

OAI22xp33_ASAP7_75t_SL g2000 ( 
.A1(n_1826),
.A2(n_1691),
.B1(n_1693),
.B2(n_1683),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1889),
.B(n_1339),
.Y(n_2001)
);

AO22x2_ASAP7_75t_L g2002 ( 
.A1(n_1846),
.A2(n_1802),
.B1(n_1857),
.B2(n_1897),
.Y(n_2002)
);

AO22x2_ASAP7_75t_L g2003 ( 
.A1(n_1928),
.A2(n_1666),
.B1(n_1667),
.B2(n_1665),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1762),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1704),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1784),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1704),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1799),
.B(n_1341),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1784),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1909),
.B(n_1548),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1982),
.A2(n_1601),
.B1(n_1348),
.B2(n_1351),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1819),
.A2(n_1348),
.B1(n_1351),
.B2(n_1341),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1712),
.Y(n_2013)
);

AO22x2_ASAP7_75t_L g2014 ( 
.A1(n_1953),
.A2(n_1673),
.B1(n_1667),
.B2(n_1409),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1784),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1978),
.B(n_1352),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_SL g2017 ( 
.A1(n_1834),
.A2(n_1673),
.B1(n_1409),
.B2(n_1413),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_SL g2018 ( 
.A1(n_1699),
.A2(n_1355),
.B1(n_1356),
.B2(n_1352),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1784),
.Y(n_2019)
);

NAND2xp33_ASAP7_75t_SL g2020 ( 
.A(n_1869),
.B(n_1355),
.Y(n_2020)
);

OR2x6_ASAP7_75t_L g2021 ( 
.A(n_1700),
.B(n_1429),
.Y(n_2021)
);

OAI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1952),
.A2(n_1838),
.B1(n_1843),
.B2(n_1822),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1982),
.A2(n_1601),
.B1(n_1365),
.B2(n_1368),
.Y(n_2023)
);

OAI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1738),
.A2(n_1368),
.B1(n_1373),
.B2(n_1356),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1777),
.A2(n_1380),
.B1(n_1381),
.B2(n_1373),
.Y(n_2025)
);

OAI22xp33_ASAP7_75t_SL g2026 ( 
.A1(n_1862),
.A2(n_1381),
.B1(n_1384),
.B2(n_1380),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1712),
.Y(n_2027)
);

OA22x2_ASAP7_75t_L g2028 ( 
.A1(n_1800),
.A2(n_1387),
.B1(n_1384),
.B2(n_1696),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1786),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1786),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1728),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1835),
.B(n_1387),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1786),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1888),
.B(n_1936),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1786),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1925),
.B(n_728),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1796),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1718),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1836),
.B(n_1850),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1718),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1796),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1936),
.B(n_1692),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1901),
.B(n_1692),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1737),
.B(n_729),
.Y(n_2044)
);

OAI22xp33_ASAP7_75t_R g2045 ( 
.A1(n_1907),
.A2(n_733),
.B1(n_736),
.B2(n_729),
.Y(n_2045)
);

OAI22xp33_ASAP7_75t_R g2046 ( 
.A1(n_1908),
.A2(n_736),
.B1(n_742),
.B2(n_733),
.Y(n_2046)
);

OR2x6_ASAP7_75t_L g2047 ( 
.A(n_1700),
.B(n_1429),
.Y(n_2047)
);

AO22x2_ASAP7_75t_L g2048 ( 
.A1(n_1918),
.A2(n_1413),
.B1(n_1408),
.B2(n_1434),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1777),
.A2(n_1696),
.B1(n_743),
.B2(n_747),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_1773),
.A2(n_743),
.B1(n_747),
.B2(n_742),
.Y(n_2050)
);

OAI22xp33_ASAP7_75t_SL g2051 ( 
.A1(n_1864),
.A2(n_867),
.B1(n_959),
.B2(n_753),
.Y(n_2051)
);

AO22x2_ASAP7_75t_L g2052 ( 
.A1(n_1918),
.A2(n_1408),
.B1(n_1453),
.B2(n_1434),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1773),
.A2(n_756),
.B1(n_867),
.B2(n_753),
.Y(n_2053)
);

OAI22xp5_ASAP7_75t_SL g2054 ( 
.A1(n_1834),
.A2(n_1456),
.B1(n_1478),
.B2(n_1453),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1901),
.B(n_1456),
.Y(n_2055)
);

OAI22xp33_ASAP7_75t_SL g2056 ( 
.A1(n_1867),
.A2(n_962),
.B1(n_963),
.B2(n_756),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1810),
.A2(n_962),
.B1(n_963),
.B2(n_959),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_1944),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1810),
.B(n_966),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1902),
.B(n_1478),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1796),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_1877),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1944),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1702),
.A2(n_969),
.B1(n_970),
.B2(n_966),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1796),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1702),
.A2(n_970),
.B1(n_972),
.B2(n_969),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1724),
.Y(n_2067)
);

OR2x6_ASAP7_75t_L g2068 ( 
.A(n_1870),
.B(n_1485),
.Y(n_2068)
);

OAI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1742),
.A2(n_1983),
.B1(n_1921),
.B2(n_1899),
.Y(n_2069)
);

OAI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1809),
.A2(n_974),
.B1(n_976),
.B2(n_972),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1724),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1729),
.Y(n_2072)
);

AO22x2_ASAP7_75t_L g2073 ( 
.A1(n_1918),
.A2(n_1489),
.B1(n_1506),
.B2(n_1485),
.Y(n_2073)
);

OAI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1983),
.A2(n_976),
.B1(n_981),
.B2(n_974),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1902),
.B(n_1489),
.Y(n_2075)
);

OAI22xp33_ASAP7_75t_SL g2076 ( 
.A1(n_1876),
.A2(n_984),
.B1(n_986),
.B2(n_981),
.Y(n_2076)
);

BUFx6f_ASAP7_75t_L g2077 ( 
.A(n_1728),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1934),
.B(n_1949),
.Y(n_2078)
);

AO22x2_ASAP7_75t_L g2079 ( 
.A1(n_1929),
.A2(n_1514),
.B1(n_1517),
.B2(n_1506),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1934),
.B(n_1514),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1716),
.Y(n_2081)
);

OAI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1899),
.A2(n_984),
.B1(n_986),
.B2(n_982),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1949),
.B(n_1517),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1908),
.B(n_1945),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1729),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1788),
.A2(n_987),
.B1(n_991),
.B2(n_982),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1730),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1856),
.B(n_1520),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1788),
.A2(n_991),
.B1(n_994),
.B2(n_987),
.Y(n_2089)
);

AO22x2_ASAP7_75t_L g2090 ( 
.A1(n_1929),
.A2(n_1932),
.B1(n_1940),
.B2(n_1935),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1809),
.A2(n_995),
.B1(n_997),
.B2(n_994),
.Y(n_2091)
);

OR2x6_ASAP7_75t_L g2092 ( 
.A(n_1870),
.B(n_1520),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1797),
.Y(n_2093)
);

INVxp67_ASAP7_75t_SL g2094 ( 
.A(n_1710),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1709),
.A2(n_997),
.B1(n_998),
.B2(n_995),
.Y(n_2095)
);

XOR2xp5_ASAP7_75t_L g2096 ( 
.A(n_1771),
.B(n_1524),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1709),
.A2(n_999),
.B1(n_1002),
.B2(n_998),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_1697),
.A2(n_1002),
.B1(n_1008),
.B2(n_999),
.Y(n_2098)
);

AO22x2_ASAP7_75t_L g2099 ( 
.A1(n_1929),
.A2(n_1525),
.B1(n_1531),
.B2(n_1524),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1797),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_SL g2101 ( 
.A1(n_1882),
.A2(n_1012),
.B1(n_1013),
.B2(n_1008),
.Y(n_2101)
);

AO22x2_ASAP7_75t_L g2102 ( 
.A1(n_1932),
.A2(n_1531),
.B1(n_1534),
.B2(n_1525),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1919),
.B(n_1534),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1943),
.B(n_1536),
.Y(n_2104)
);

OAI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_1899),
.A2(n_1012),
.B1(n_1013),
.B2(n_1011),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1730),
.Y(n_2106)
);

AO22x2_ASAP7_75t_L g2107 ( 
.A1(n_1932),
.A2(n_1565),
.B1(n_1576),
.B2(n_1536),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1946),
.B(n_1565),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1797),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1879),
.B(n_1576),
.Y(n_2110)
);

OAI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_1899),
.A2(n_1014),
.B1(n_1017),
.B2(n_1011),
.Y(n_2111)
);

INVx2_ASAP7_75t_SL g2112 ( 
.A(n_1877),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1925),
.B(n_1895),
.Y(n_2113)
);

XNOR2xp5_ASAP7_75t_L g2114 ( 
.A(n_1771),
.B(n_1577),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1879),
.B(n_1577),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1797),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1801),
.Y(n_2117)
);

AO22x2_ASAP7_75t_L g2118 ( 
.A1(n_1940),
.A2(n_1589),
.B1(n_1591),
.B2(n_1578),
.Y(n_2118)
);

OAI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_1774),
.A2(n_1017),
.B1(n_1019),
.B2(n_1014),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1697),
.A2(n_1020),
.B1(n_1022),
.B2(n_1019),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1697),
.A2(n_1022),
.B1(n_1023),
.B2(n_1020),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1733),
.A2(n_1025),
.B1(n_1024),
.B2(n_1257),
.Y(n_2122)
);

OAI22xp33_ASAP7_75t_SL g2123 ( 
.A1(n_1935),
.A2(n_1024),
.B1(n_1025),
.B2(n_1286),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1801),
.Y(n_2124)
);

OAI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_1809),
.A2(n_1246),
.B1(n_1114),
.B2(n_1181),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1830),
.Y(n_2126)
);

INVx8_ASAP7_75t_L g2127 ( 
.A(n_1925),
.Y(n_2127)
);

XNOR2xp5_ASAP7_75t_L g2128 ( 
.A(n_1892),
.B(n_1578),
.Y(n_2128)
);

OAI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1883),
.A2(n_1263),
.B1(n_1264),
.B2(n_1260),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1801),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_1716),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_1733),
.A2(n_1268),
.B1(n_1273),
.B2(n_1266),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1830),
.Y(n_2133)
);

NOR2x1p5_ASAP7_75t_L g2134 ( 
.A(n_1764),
.B(n_1276),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1965),
.B(n_1591),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1801),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1925),
.B(n_1241),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1782),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1716),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_1756),
.Y(n_2140)
);

AO22x2_ASAP7_75t_L g2141 ( 
.A1(n_1940),
.A2(n_1589),
.B1(n_1598),
.B2(n_1592),
.Y(n_2141)
);

OAI22xp33_ASAP7_75t_SL g2142 ( 
.A1(n_1912),
.A2(n_1280),
.B1(n_1281),
.B2(n_1278),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1883),
.B(n_1592),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1931),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1815),
.A2(n_1246),
.B1(n_1114),
.B2(n_1181),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_1713),
.A2(n_1287),
.B1(n_1289),
.B2(n_1285),
.Y(n_2146)
);

OAI22xp33_ASAP7_75t_SL g2147 ( 
.A1(n_1912),
.A2(n_1099),
.B1(n_1100),
.B2(n_1096),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_1790),
.B(n_1598),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1713),
.A2(n_1106),
.B1(n_1105),
.B2(n_1174),
.Y(n_2149)
);

AOI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_1713),
.A2(n_1194),
.B1(n_1205),
.B2(n_1182),
.Y(n_2150)
);

AO22x2_ASAP7_75t_L g2151 ( 
.A1(n_1924),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1754),
.A2(n_1194),
.B1(n_1205),
.B2(n_1182),
.Y(n_2152)
);

AO22x2_ASAP7_75t_L g2153 ( 
.A1(n_1924),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_1754),
.A2(n_1256),
.B1(n_1277),
.B2(n_1207),
.Y(n_2154)
);

OAI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1883),
.A2(n_1256),
.B1(n_1277),
.B2(n_1207),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1811),
.Y(n_2156)
);

OA22x2_ASAP7_75t_L g2157 ( 
.A1(n_1800),
.A2(n_1288),
.B1(n_1296),
.B2(n_1283),
.Y(n_2157)
);

AO22x2_ASAP7_75t_L g2158 ( 
.A1(n_1941),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_1925),
.B(n_7),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1754),
.A2(n_1283),
.B1(n_1296),
.B2(n_1288),
.Y(n_2160)
);

AO22x2_ASAP7_75t_L g2161 ( 
.A1(n_1941),
.A2(n_1959),
.B1(n_1973),
.B2(n_1960),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1880),
.A2(n_1308),
.B1(n_1314),
.B2(n_1241),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_1880),
.A2(n_1308),
.B1(n_1314),
.B2(n_1241),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_SL g2164 ( 
.A1(n_1959),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2164)
);

INVx1_ASAP7_75t_SL g2165 ( 
.A(n_1842),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1763),
.B(n_1314),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1880),
.A2(n_1229),
.B1(n_1247),
.B2(n_1223),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1763),
.B(n_8),
.Y(n_2168)
);

OA22x2_ASAP7_75t_L g2169 ( 
.A1(n_1775),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_1747),
.A2(n_1247),
.B1(n_1301),
.B2(n_1229),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_1747),
.A2(n_1247),
.B1(n_1301),
.B2(n_1229),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1769),
.B(n_1869),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1782),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_1769),
.B(n_9),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1783),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1783),
.Y(n_2176)
);

OAI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_1960),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2177)
);

OAI22xp33_ASAP7_75t_L g2178 ( 
.A1(n_1892),
.A2(n_1247),
.B1(n_1301),
.B2(n_1229),
.Y(n_2178)
);

OAI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_1869),
.A2(n_1304),
.B1(n_1301),
.B2(n_13),
.Y(n_2179)
);

OR2x6_ASAP7_75t_L g2180 ( 
.A(n_1972),
.B(n_1304),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1798),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1811),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1906),
.B(n_11),
.Y(n_2183)
);

OAI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_1973),
.A2(n_1985),
.B1(n_1955),
.B2(n_1958),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1811),
.Y(n_2185)
);

AO22x2_ASAP7_75t_L g2186 ( 
.A1(n_1985),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1811),
.Y(n_2187)
);

AO22x2_ASAP7_75t_L g2188 ( 
.A1(n_1863),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_2188)
);

OAI22xp33_ASAP7_75t_L g2189 ( 
.A1(n_1911),
.A2(n_1304),
.B1(n_16),
.B2(n_14),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1906),
.B(n_14),
.Y(n_2190)
);

OAI22xp33_ASAP7_75t_SL g2191 ( 
.A1(n_1904),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2191)
);

OAI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_1911),
.A2(n_1304),
.B1(n_19),
.B2(n_17),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1830),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1853),
.Y(n_2194)
);

OA22x2_ASAP7_75t_L g2195 ( 
.A1(n_1886),
.A2(n_1967),
.B1(n_1969),
.B2(n_1714),
.Y(n_2195)
);

OAI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_1911),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2196)
);

AO22x2_ASAP7_75t_L g2197 ( 
.A1(n_1863),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1906),
.B(n_1914),
.Y(n_2198)
);

OAI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_1911),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2199)
);

AND2x2_ASAP7_75t_SL g2200 ( 
.A(n_1976),
.B(n_21),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_1831),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2201)
);

OAI22xp33_ASAP7_75t_SL g2202 ( 
.A1(n_1905),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_2202)
);

OAI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1955),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1824),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1914),
.B(n_1933),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1914),
.B(n_24),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1853),
.Y(n_2207)
);

OA22x2_ASAP7_75t_L g2208 ( 
.A1(n_1900),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1853),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1933),
.B(n_26),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_SL g2211 ( 
.A1(n_1900),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1829),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_1895),
.B(n_27),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_1877),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1955),
.B(n_129),
.Y(n_2215)
);

AO22x2_ASAP7_75t_L g2216 ( 
.A1(n_1863),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_1971),
.B(n_29),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1829),
.Y(n_2218)
);

AO22x2_ASAP7_75t_L g2219 ( 
.A1(n_1831),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2219)
);

OA22x2_ASAP7_75t_L g2220 ( 
.A1(n_1913),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_1933),
.B(n_33),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_SL g2222 ( 
.A1(n_1931),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2222)
);

INVx4_ASAP7_75t_L g2223 ( 
.A(n_1895),
.Y(n_2223)
);

OR2x6_ASAP7_75t_L g2224 ( 
.A(n_1955),
.B(n_33),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1831),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1947),
.B(n_36),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_1840),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1860),
.Y(n_2228)
);

OAI22xp33_ASAP7_75t_SL g2229 ( 
.A1(n_1915),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1860),
.Y(n_2230)
);

OAI22xp33_ASAP7_75t_R g2231 ( 
.A1(n_1917),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1824),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_1947),
.B(n_39),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1824),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1716),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_1840),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2236)
);

OAI22xp33_ASAP7_75t_SL g2237 ( 
.A1(n_1920),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2237)
);

OAI22xp33_ASAP7_75t_L g2238 ( 
.A1(n_1958),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2238)
);

OAI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_1958),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2239)
);

AO22x2_ASAP7_75t_L g2240 ( 
.A1(n_1840),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_1844),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1824),
.Y(n_2242)
);

OAI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_1958),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1947),
.B(n_47),
.Y(n_2244)
);

AND2x2_ASAP7_75t_SL g2245 ( 
.A(n_1976),
.B(n_48),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_SL g2246 ( 
.A1(n_1922),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2246)
);

INVx8_ASAP7_75t_L g2247 ( 
.A(n_1877),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_1844),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2248)
);

OAI22xp33_ASAP7_75t_SL g2249 ( 
.A1(n_1923),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_2249)
);

AO22x2_ASAP7_75t_L g2250 ( 
.A1(n_1844),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1757),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_2251)
);

OR2x6_ASAP7_75t_L g2252 ( 
.A(n_1966),
.B(n_55),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1798),
.Y(n_2253)
);

AO22x2_ASAP7_75t_L g2254 ( 
.A1(n_1806),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_2254)
);

OAI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_1966),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_1815),
.A2(n_132),
.B1(n_133),
.B2(n_130),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_1954),
.B(n_56),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1954),
.B(n_57),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1807),
.Y(n_2259)
);

OAI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_1966),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2260)
);

AO22x2_ASAP7_75t_L g2261 ( 
.A1(n_1806),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_1806),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1807),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1821),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1825),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1825),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_1821),
.A2(n_1837),
.B1(n_1849),
.B2(n_1815),
.Y(n_2267)
);

OR2x6_ASAP7_75t_L g2268 ( 
.A(n_1966),
.B(n_63),
.Y(n_2268)
);

AO22x2_ASAP7_75t_L g2269 ( 
.A1(n_1821),
.A2(n_66),
.B1(n_63),
.B2(n_65),
.Y(n_2269)
);

OR2x6_ASAP7_75t_L g2270 ( 
.A(n_1984),
.B(n_65),
.Y(n_2270)
);

AO22x2_ASAP7_75t_L g2271 ( 
.A1(n_1791),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_1765),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1954),
.B(n_66),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1981),
.B(n_1984),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_1837),
.A2(n_1849),
.B1(n_1833),
.B2(n_1825),
.Y(n_2275)
);

OAI22xp33_ASAP7_75t_SL g2276 ( 
.A1(n_1926),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_1981),
.B(n_67),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_1837),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_1877),
.Y(n_2279)
);

AO22x2_ASAP7_75t_L g2280 ( 
.A1(n_1791),
.A2(n_1804),
.B1(n_1938),
.B2(n_1930),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1825),
.Y(n_2281)
);

OR2x6_ASAP7_75t_L g2282 ( 
.A(n_1984),
.B(n_1910),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_1728),
.Y(n_2283)
);

BUFx10_ASAP7_75t_L g2284 ( 
.A(n_1984),
.Y(n_2284)
);

INVx1_ASAP7_75t_SL g2285 ( 
.A(n_1884),
.Y(n_2285)
);

INVx2_ASAP7_75t_SL g2286 ( 
.A(n_1884),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_SL g2287 ( 
.A1(n_1939),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2287)
);

AND2x2_ASAP7_75t_SL g2288 ( 
.A(n_1770),
.B(n_70),
.Y(n_2288)
);

OAI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_1975),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2289)
);

OAI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1950),
.A2(n_1951),
.B1(n_1957),
.B2(n_1956),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1860),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_1849),
.A2(n_1708),
.B1(n_1717),
.B2(n_1698),
.Y(n_2292)
);

OAI22xp33_ASAP7_75t_SL g2293 ( 
.A1(n_1961),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_2293)
);

AO22x2_ASAP7_75t_L g2294 ( 
.A1(n_1791),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2294)
);

OAI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_1962),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1981),
.B(n_75),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_1884),
.B(n_76),
.Y(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_1963),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_2298)
);

OAI22xp33_ASAP7_75t_SL g2299 ( 
.A1(n_1974),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2299)
);

AO22x2_ASAP7_75t_L g2300 ( 
.A1(n_1804),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_SL g2301 ( 
.A1(n_1979),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_SL g2302 ( 
.A1(n_1980),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_2302)
);

INVxp67_ASAP7_75t_L g2303 ( 
.A(n_1859),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_1895),
.B(n_81),
.Y(n_2304)
);

INVx2_ASAP7_75t_SL g2305 ( 
.A(n_1884),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1884),
.B(n_82),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1993),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_1991),
.B(n_1865),
.Y(n_2308)
);

XNOR2xp5_ASAP7_75t_L g2309 ( 
.A(n_2096),
.B(n_1872),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2005),
.Y(n_2310)
);

NAND3xp33_ASAP7_75t_L g2311 ( 
.A(n_1990),
.B(n_1745),
.C(n_1823),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2126),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2005),
.Y(n_2313)
);

INVx2_ASAP7_75t_SL g2314 ( 
.A(n_2284),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2069),
.B(n_1725),
.Y(n_2315)
);

INVx4_ASAP7_75t_L g2316 ( 
.A(n_2247),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2078),
.B(n_1820),
.Y(n_2317)
);

INVx5_ASAP7_75t_L g2318 ( 
.A(n_2247),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2059),
.B(n_1820),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_2063),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2007),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2303),
.B(n_1781),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2010),
.B(n_1787),
.Y(n_2323)
);

NAND2xp33_ASAP7_75t_L g2324 ( 
.A(n_2127),
.B(n_1725),
.Y(n_2324)
);

INVxp33_ASAP7_75t_L g2325 ( 
.A(n_2008),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2126),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2007),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_1998),
.A2(n_1828),
.B1(n_1845),
.B2(n_1827),
.Y(n_2328)
);

INVx2_ASAP7_75t_SL g2329 ( 
.A(n_2284),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2022),
.B(n_1903),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2133),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2013),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2223),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2267),
.B(n_1725),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2275),
.B(n_1725),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2133),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2084),
.B(n_1805),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_1987),
.B(n_2034),
.Y(n_2338)
);

NAND3xp33_ASAP7_75t_L g2339 ( 
.A(n_2025),
.B(n_1858),
.C(n_1833),
.Y(n_2339)
);

INVx4_ASAP7_75t_L g2340 ( 
.A(n_2127),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_2223),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2184),
.B(n_1725),
.Y(n_2342)
);

NAND2xp33_ASAP7_75t_L g2343 ( 
.A(n_2198),
.B(n_1719),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2193),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2200),
.B(n_1728),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2245),
.B(n_1833),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2013),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2027),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2172),
.A2(n_1804),
.B1(n_1858),
.B2(n_1833),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2027),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2031),
.B(n_1858),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2205),
.B(n_1865),
.Y(n_2352)
);

OR2x6_ASAP7_75t_L g2353 ( 
.A(n_2068),
.B(n_1770),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2193),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2044),
.B(n_1887),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2194),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2031),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2031),
.B(n_1858),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2085),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2085),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2087),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_2077),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2087),
.Y(n_2363)
);

OR2x6_ASAP7_75t_L g2364 ( 
.A(n_2068),
.B(n_1770),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1994),
.B(n_1887),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2106),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2106),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2194),
.Y(n_2368)
);

BUFx3_ASAP7_75t_L g2369 ( 
.A(n_2113),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2207),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2077),
.B(n_1868),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2038),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2001),
.B(n_1731),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2207),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2040),
.Y(n_2375)
);

INVxp67_ASAP7_75t_L g2376 ( 
.A(n_2042),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2067),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_2113),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2209),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_2140),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_1995),
.B(n_2016),
.Y(n_2381)
);

AND2x4_ASAP7_75t_SL g2382 ( 
.A(n_2282),
.B(n_1764),
.Y(n_2382)
);

INVx4_ASAP7_75t_L g2383 ( 
.A(n_1986),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2077),
.B(n_1868),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_L g2385 ( 
.A1(n_1998),
.A2(n_1828),
.B1(n_1845),
.B2(n_1827),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2166),
.B(n_1868),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2271),
.A2(n_1852),
.B1(n_1855),
.B2(n_1848),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2004),
.Y(n_2388)
);

CKINVDCx20_ASAP7_75t_R g2389 ( 
.A(n_2017),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2209),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_2272),
.Y(n_2391)
);

OR2x6_ASAP7_75t_L g2392 ( 
.A(n_2092),
.B(n_2021),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2071),
.Y(n_2393)
);

INVxp67_ASAP7_75t_L g2394 ( 
.A(n_2055),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_1992),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2072),
.Y(n_2396)
);

BUFx3_ASAP7_75t_L g2397 ( 
.A(n_2144),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1992),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2011),
.B(n_2023),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_1999),
.Y(n_2400)
);

OAI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2262),
.A2(n_1874),
.B1(n_1881),
.B2(n_1868),
.Y(n_2401)
);

AOI22xp33_ASAP7_75t_L g2402 ( 
.A1(n_2271),
.A2(n_1852),
.B1(n_1855),
.B2(n_1848),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_2274),
.B(n_1895),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2138),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_2114),
.Y(n_2405)
);

AND3x2_ASAP7_75t_L g2406 ( 
.A(n_2080),
.B(n_1765),
.C(n_1861),
.Y(n_2406)
);

BUFx8_ASAP7_75t_SL g2407 ( 
.A(n_2021),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_1999),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_1997),
.B(n_1759),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2173),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2175),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_2283),
.Y(n_2412)
);

AOI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_2294),
.A2(n_1893),
.B1(n_1896),
.B2(n_1891),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2060),
.B(n_1759),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2176),
.Y(n_2415)
);

BUFx10_ASAP7_75t_L g2416 ( 
.A(n_2104),
.Y(n_2416)
);

AOI22xp33_ASAP7_75t_L g2417 ( 
.A1(n_2294),
.A2(n_1893),
.B1(n_1896),
.B2(n_1891),
.Y(n_2417)
);

BUFx6f_ASAP7_75t_L g2418 ( 
.A(n_2283),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2181),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2094),
.B(n_1874),
.Y(n_2420)
);

AO22x2_ASAP7_75t_L g2421 ( 
.A1(n_2168),
.A2(n_1866),
.B1(n_1861),
.B2(n_1813),
.Y(n_2421)
);

INVxp67_ASAP7_75t_L g2422 ( 
.A(n_2075),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2253),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2259),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2110),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2263),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2283),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2228),
.Y(n_2428)
);

INVx4_ASAP7_75t_L g2429 ( 
.A(n_2282),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2132),
.Y(n_2430)
);

CKINVDCx20_ASAP7_75t_R g2431 ( 
.A(n_2128),
.Y(n_2431)
);

BUFx10_ASAP7_75t_L g2432 ( 
.A(n_2108),
.Y(n_2432)
);

NOR2x1p5_ASAP7_75t_L g2433 ( 
.A(n_2039),
.B(n_2148),
.Y(n_2433)
);

NAND2xp33_ASAP7_75t_L g2434 ( 
.A(n_2020),
.B(n_1722),
.Y(n_2434)
);

OR2x6_ASAP7_75t_L g2435 ( 
.A(n_2092),
.B(n_1874),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_2081),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2228),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2230),
.Y(n_2438)
);

BUFx3_ASAP7_75t_L g2439 ( 
.A(n_2115),
.Y(n_2439)
);

CKINVDCx16_ASAP7_75t_R g2440 ( 
.A(n_2054),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2150),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_2047),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2290),
.B(n_1874),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2152),
.Y(n_2444)
);

OAI22x1_ASAP7_75t_L g2445 ( 
.A1(n_2049),
.A2(n_1866),
.B1(n_1927),
.B2(n_1916),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2183),
.B(n_1890),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2190),
.B(n_1890),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2206),
.B(n_1890),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_1988),
.B(n_1881),
.Y(n_2449)
);

AOI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2045),
.A2(n_1890),
.B1(n_1894),
.B2(n_1881),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2210),
.B(n_1894),
.Y(n_2451)
);

OAI21xp33_ASAP7_75t_SL g2452 ( 
.A1(n_2288),
.A2(n_1977),
.B(n_1871),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2081),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2154),
.Y(n_2454)
);

INVx4_ASAP7_75t_L g2455 ( 
.A(n_2159),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2135),
.B(n_1881),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2160),
.Y(n_2457)
);

XNOR2xp5_ASAP7_75t_L g2458 ( 
.A(n_1989),
.B(n_1916),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2131),
.B(n_1894),
.Y(n_2459)
);

INVx2_ASAP7_75t_SL g2460 ( 
.A(n_2165),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2043),
.B(n_1710),
.Y(n_2461)
);

AOI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_2045),
.A2(n_1894),
.B1(n_1927),
.B2(n_1916),
.Y(n_2462)
);

BUFx3_ASAP7_75t_L g2463 ( 
.A(n_2047),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_2018),
.B(n_1817),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_2058),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2280),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2280),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2221),
.B(n_2226),
.Y(n_2468)
);

BUFx3_ASAP7_75t_L g2469 ( 
.A(n_2131),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2230),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2291),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2233),
.B(n_1851),
.Y(n_2472)
);

BUFx6f_ASAP7_75t_L g2473 ( 
.A(n_2139),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2149),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2244),
.B(n_1873),
.Y(n_2475)
);

BUFx10_ASAP7_75t_L g2476 ( 
.A(n_2159),
.Y(n_2476)
);

INVxp33_ASAP7_75t_L g2477 ( 
.A(n_2088),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2291),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_2139),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2257),
.B(n_1875),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2161),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_2235),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2143),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2258),
.B(n_2273),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2161),
.Y(n_2485)
);

OR2x6_ASAP7_75t_L g2486 ( 
.A(n_2224),
.B(n_1812),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2212),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2146),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2006),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2009),
.Y(n_2490)
);

HB1xp67_ASAP7_75t_L g2491 ( 
.A(n_1996),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2212),
.Y(n_2492)
);

INVx2_ASAP7_75t_SL g2493 ( 
.A(n_2180),
.Y(n_2493)
);

INVx4_ASAP7_75t_L g2494 ( 
.A(n_2213),
.Y(n_2494)
);

INVx1_ASAP7_75t_SL g2495 ( 
.A(n_2103),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2015),
.Y(n_2496)
);

INVx3_ASAP7_75t_L g2497 ( 
.A(n_2235),
.Y(n_2497)
);

CKINVDCx16_ASAP7_75t_R g2498 ( 
.A(n_2083),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2218),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2019),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2218),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2029),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2030),
.Y(n_2503)
);

BUFx3_ASAP7_75t_L g2504 ( 
.A(n_2062),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2033),
.Y(n_2505)
);

AND3x2_ASAP7_75t_L g2506 ( 
.A(n_2032),
.B(n_1765),
.C(n_1814),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2035),
.Y(n_2507)
);

BUFx2_ASAP7_75t_L g2508 ( 
.A(n_2180),
.Y(n_2508)
);

AND2x4_ASAP7_75t_L g2509 ( 
.A(n_2134),
.B(n_1816),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2037),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2277),
.B(n_1832),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2041),
.Y(n_2512)
);

AOI22xp33_ASAP7_75t_L g2513 ( 
.A1(n_2300),
.A2(n_1927),
.B1(n_1942),
.B2(n_1937),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2296),
.B(n_1878),
.Y(n_2514)
);

AND2x6_ASAP7_75t_L g2515 ( 
.A(n_2213),
.B(n_1885),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2061),
.Y(n_2516)
);

NAND3xp33_ASAP7_75t_L g2517 ( 
.A(n_2050),
.B(n_1898),
.C(n_1753),
.Y(n_2517)
);

OR2x6_ASAP7_75t_L g2518 ( 
.A(n_2224),
.B(n_1701),
.Y(n_2518)
);

AOI21x1_ASAP7_75t_L g2519 ( 
.A1(n_2292),
.A2(n_1977),
.B(n_1818),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2057),
.B(n_1732),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2065),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2304),
.B(n_1898),
.Y(n_2522)
);

BUFx3_ASAP7_75t_L g2523 ( 
.A(n_2112),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2093),
.Y(n_2524)
);

INVx4_ASAP7_75t_L g2525 ( 
.A(n_2304),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2300),
.A2(n_1942),
.B1(n_1937),
.B2(n_1948),
.Y(n_2526)
);

BUFx4f_ASAP7_75t_L g2527 ( 
.A(n_2252),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2100),
.Y(n_2528)
);

CKINVDCx16_ASAP7_75t_R g2529 ( 
.A(n_2252),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_L g2530 ( 
.A1(n_2254),
.A2(n_2269),
.B1(n_2261),
.B2(n_2240),
.Y(n_2530)
);

BUFx8_ASAP7_75t_SL g2531 ( 
.A(n_2268),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2109),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2116),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_SL g2534 ( 
.A(n_2268),
.B(n_1839),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2117),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2174),
.B(n_1739),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2124),
.Y(n_2537)
);

INVx5_ASAP7_75t_L g2538 ( 
.A(n_2214),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2130),
.B(n_1898),
.Y(n_2539)
);

INVx2_ASAP7_75t_SL g2540 ( 
.A(n_2090),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_2136),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2156),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2182),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2000),
.Y(n_2544)
);

OR2x2_ASAP7_75t_L g2545 ( 
.A(n_2053),
.B(n_1743),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2217),
.B(n_1758),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2185),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2187),
.Y(n_2548)
);

INVxp67_ASAP7_75t_SL g2549 ( 
.A(n_2204),
.Y(n_2549)
);

AOI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2254),
.A2(n_1942),
.B1(n_1937),
.B2(n_1948),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2119),
.B(n_1803),
.Y(n_2551)
);

BUFx6f_ASAP7_75t_L g2552 ( 
.A(n_2232),
.Y(n_2552)
);

INVx2_ASAP7_75t_SL g2553 ( 
.A(n_2090),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2285),
.B(n_1779),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2129),
.B(n_1785),
.Y(n_2555)
);

INVx4_ASAP7_75t_L g2556 ( 
.A(n_2270),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2234),
.Y(n_2557)
);

INVx3_ASAP7_75t_L g2558 ( 
.A(n_2242),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2265),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2266),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2046),
.A2(n_1792),
.B1(n_1793),
.B2(n_1789),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2122),
.B(n_1794),
.Y(n_2562)
);

XNOR2xp5_ASAP7_75t_L g2563 ( 
.A(n_1989),
.B(n_1795),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2024),
.B(n_1721),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2281),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2297),
.B(n_1898),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2306),
.B(n_1898),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2279),
.B(n_1948),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_L g2569 ( 
.A(n_2305),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_2098),
.B(n_1721),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2125),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2286),
.B(n_1964),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2123),
.B(n_1721),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2145),
.Y(n_2574)
);

INVxp67_ASAP7_75t_L g2575 ( 
.A(n_2079),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2151),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2157),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2002),
.B(n_1964),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2151),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2261),
.A2(n_1964),
.B1(n_1970),
.B2(n_1968),
.Y(n_2580)
);

INVxp33_ASAP7_75t_L g2581 ( 
.A(n_2079),
.Y(n_2581)
);

INVx1_ASAP7_75t_SL g2582 ( 
.A(n_2270),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2153),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2142),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2153),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2086),
.B(n_1968),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2147),
.Y(n_2587)
);

INVx2_ASAP7_75t_SL g2588 ( 
.A(n_2048),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2167),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2278),
.Y(n_2590)
);

INVx4_ASAP7_75t_SL g2591 ( 
.A(n_2222),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2158),
.Y(n_2592)
);

NOR2x1p5_ASAP7_75t_L g2593 ( 
.A(n_2002),
.B(n_1776),
.Y(n_2593)
);

INVxp67_ASAP7_75t_SL g2594 ( 
.A(n_2082),
.Y(n_2594)
);

AND2x4_ASAP7_75t_L g2595 ( 
.A(n_2036),
.B(n_1839),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2269),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2105),
.B(n_1968),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2251),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2158),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2186),
.Y(n_2600)
);

NOR2xp33_ASAP7_75t_L g2601 ( 
.A(n_2120),
.B(n_1721),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2186),
.Y(n_2602)
);

OAI21xp33_ASAP7_75t_SL g2603 ( 
.A1(n_2264),
.A2(n_2225),
.B(n_2201),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2219),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2012),
.B(n_1723),
.Y(n_2605)
);

AND2x6_ASAP7_75t_L g2606 ( 
.A(n_2227),
.B(n_1734),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_2026),
.Y(n_2607)
);

NAND2xp33_ASAP7_75t_R g2608 ( 
.A(n_2046),
.B(n_1970),
.Y(n_2608)
);

AND2x4_ASAP7_75t_L g2609 ( 
.A(n_2215),
.B(n_1839),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2048),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2111),
.B(n_1723),
.Y(n_2611)
);

BUFx10_ASAP7_75t_L g2612 ( 
.A(n_2195),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2220),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2219),
.A2(n_1970),
.B1(n_1839),
.B2(n_1723),
.Y(n_2614)
);

BUFx2_ASAP7_75t_L g2615 ( 
.A(n_2099),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2240),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2236),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2137),
.B(n_2121),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_SL g2619 ( 
.A(n_2155),
.B(n_1723),
.Y(n_2619)
);

INVx3_ASAP7_75t_L g2620 ( 
.A(n_2250),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2241),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2089),
.B(n_1727),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2248),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2250),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2064),
.B(n_1727),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2188),
.Y(n_2626)
);

INVxp67_ASAP7_75t_SL g2627 ( 
.A(n_2189),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2188),
.Y(n_2628)
);

CKINVDCx20_ASAP7_75t_R g2629 ( 
.A(n_2211),
.Y(n_2629)
);

AND2x6_ASAP7_75t_L g2630 ( 
.A(n_2162),
.B(n_1734),
.Y(n_2630)
);

AOI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2231),
.A2(n_1839),
.B1(n_1727),
.B2(n_1818),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2099),
.Y(n_2632)
);

NOR2xp33_ASAP7_75t_L g2633 ( 
.A(n_2066),
.B(n_1727),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2051),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2192),
.B(n_1772),
.Y(n_2635)
);

BUFx10_ASAP7_75t_L g2636 ( 
.A(n_2074),
.Y(n_2636)
);

BUFx3_ASAP7_75t_L g2637 ( 
.A(n_2052),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2095),
.B(n_1720),
.Y(n_2638)
);

NOR2xp33_ASAP7_75t_L g2639 ( 
.A(n_2097),
.B(n_2056),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2052),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2014),
.B(n_1720),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2070),
.B(n_1808),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_2076),
.B(n_1808),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_2196),
.B(n_1772),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2199),
.B(n_1772),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2101),
.B(n_1808),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2197),
.Y(n_2647)
);

INVx3_ASAP7_75t_L g2648 ( 
.A(n_2197),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2216),
.Y(n_2649)
);

BUFx6f_ASAP7_75t_L g2650 ( 
.A(n_2216),
.Y(n_2650)
);

AND2x6_ASAP7_75t_L g2651 ( 
.A(n_2163),
.B(n_1735),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2170),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2169),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2256),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2208),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2171),
.Y(n_2656)
);

BUFx4f_ASAP7_75t_L g2657 ( 
.A(n_2231),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2091),
.B(n_1818),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2246),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2203),
.Y(n_2660)
);

CKINVDCx6p67_ASAP7_75t_R g2661 ( 
.A(n_2102),
.Y(n_2661)
);

BUFx2_ASAP7_75t_L g2662 ( 
.A(n_2465),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2317),
.B(n_2028),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2372),
.Y(n_2664)
);

OAI221xp5_ASAP7_75t_L g2665 ( 
.A1(n_2399),
.A2(n_2381),
.B1(n_2657),
.B2(n_2603),
.C(n_2338),
.Y(n_2665)
);

AND2x6_ASAP7_75t_L g2666 ( 
.A(n_2650),
.B(n_1720),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2375),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2612),
.B(n_2365),
.Y(n_2668)
);

INVx1_ASAP7_75t_SL g2669 ( 
.A(n_2380),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2432),
.B(n_2179),
.Y(n_2670)
);

AND2x6_ASAP7_75t_L g2671 ( 
.A(n_2650),
.B(n_1751),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2377),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2419),
.Y(n_2673)
);

INVx4_ASAP7_75t_SL g2674 ( 
.A(n_2515),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2330),
.B(n_1751),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2393),
.Y(n_2676)
);

INVxp67_ASAP7_75t_SL g2677 ( 
.A(n_2395),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2396),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2419),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2432),
.B(n_2238),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2310),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2313),
.Y(n_2682)
);

OR2x6_ASAP7_75t_L g2683 ( 
.A(n_2486),
.B(n_2102),
.Y(n_2683)
);

AO22x2_ASAP7_75t_L g2684 ( 
.A1(n_2604),
.A2(n_2014),
.B1(n_2003),
.B2(n_2107),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2404),
.Y(n_2685)
);

INVxp33_ASAP7_75t_L g2686 ( 
.A(n_2491),
.Y(n_2686)
);

INVx2_ASAP7_75t_SL g2687 ( 
.A(n_2397),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2612),
.B(n_2003),
.Y(n_2688)
);

NAND3xp33_ASAP7_75t_L g2689 ( 
.A(n_2399),
.B(n_2243),
.C(n_2239),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2410),
.Y(n_2690)
);

CKINVDCx20_ASAP7_75t_R g2691 ( 
.A(n_2465),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2381),
.B(n_2287),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2411),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2415),
.Y(n_2694)
);

INVxp67_ASAP7_75t_L g2695 ( 
.A(n_2460),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2330),
.B(n_1751),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2321),
.Y(n_2697)
);

INVx1_ASAP7_75t_SL g2698 ( 
.A(n_2409),
.Y(n_2698)
);

A2O1A1Ixp33_ASAP7_75t_L g2699 ( 
.A1(n_2551),
.A2(n_1776),
.B(n_1736),
.C(n_1740),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2612),
.B(n_2107),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2423),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2424),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2327),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2426),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2325),
.B(n_2301),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2332),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2369),
.B(n_1776),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_2325),
.B(n_2302),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2347),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2323),
.B(n_2295),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2348),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_2397),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2350),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2359),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2498),
.B(n_2298),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2360),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2495),
.B(n_2118),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2338),
.B(n_2191),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2416),
.B(n_2255),
.Y(n_2719)
);

INVxp67_ASAP7_75t_L g2720 ( 
.A(n_2443),
.Y(n_2720)
);

INVx1_ASAP7_75t_SL g2721 ( 
.A(n_2320),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2369),
.B(n_1735),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2361),
.Y(n_2723)
);

INVxp67_ASAP7_75t_L g2724 ( 
.A(n_2443),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2363),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2366),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2319),
.B(n_1736),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2308),
.B(n_2118),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2455),
.B(n_1740),
.Y(n_2729)
);

OAI221xp5_ASAP7_75t_L g2730 ( 
.A1(n_2657),
.A2(n_2202),
.B1(n_2249),
.B2(n_2237),
.C(n_2229),
.Y(n_2730)
);

AND2x6_ASAP7_75t_L g2731 ( 
.A(n_2650),
.B(n_1772),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2414),
.B(n_2141),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2416),
.B(n_2260),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2367),
.Y(n_2734)
);

INVxp67_ASAP7_75t_SL g2735 ( 
.A(n_2395),
.Y(n_2735)
);

INVxp67_ASAP7_75t_L g2736 ( 
.A(n_2461),
.Y(n_2736)
);

INVx8_ASAP7_75t_L g2737 ( 
.A(n_2318),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2577),
.Y(n_2738)
);

BUFx4_ASAP7_75t_L g2739 ( 
.A(n_2407),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2659),
.B(n_2141),
.Y(n_2740)
);

NAND2x1p5_ASAP7_75t_L g2741 ( 
.A(n_2318),
.B(n_1748),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2318),
.Y(n_2742)
);

INVx3_ASAP7_75t_L g2743 ( 
.A(n_2318),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2466),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2340),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2337),
.B(n_1744),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2416),
.B(n_2164),
.Y(n_2747)
);

BUFx2_ASAP7_75t_L g2748 ( 
.A(n_2435),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2467),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2481),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2357),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2386),
.B(n_1744),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2394),
.Y(n_2753)
);

INVx8_ASAP7_75t_L g2754 ( 
.A(n_2515),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2312),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2312),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2326),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2326),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2331),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2386),
.B(n_1746),
.Y(n_2760)
);

NAND2x1p5_ASAP7_75t_L g2761 ( 
.A(n_2378),
.B(n_1748),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2331),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2659),
.B(n_2073),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2477),
.B(n_2276),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2336),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2382),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2388),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2455),
.B(n_1746),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2551),
.B(n_1749),
.Y(n_2769)
);

AO22x2_ASAP7_75t_L g2770 ( 
.A1(n_2604),
.A2(n_2610),
.B1(n_2637),
.B2(n_2588),
.Y(n_2770)
);

AND2x6_ASAP7_75t_L g2771 ( 
.A(n_2650),
.B(n_1778),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2485),
.Y(n_2772)
);

OAI22xp5_ASAP7_75t_SL g2773 ( 
.A1(n_2629),
.A2(n_2073),
.B1(n_2299),
.B2(n_2293),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2576),
.Y(n_2774)
);

NAND3x1_ASAP7_75t_L g2775 ( 
.A(n_2620),
.B(n_2177),
.C(n_2289),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2456),
.B(n_1749),
.Y(n_2776)
);

INVx8_ASAP7_75t_L g2777 ( 
.A(n_2515),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2477),
.B(n_1778),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2422),
.B(n_2376),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2576),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2579),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2336),
.Y(n_2782)
);

INVx2_ASAP7_75t_SL g2783 ( 
.A(n_2382),
.Y(n_2783)
);

INVx4_ASAP7_75t_L g2784 ( 
.A(n_2316),
.Y(n_2784)
);

INVx2_ASAP7_75t_SL g2785 ( 
.A(n_2527),
.Y(n_2785)
);

BUFx6f_ASAP7_75t_L g2786 ( 
.A(n_2357),
.Y(n_2786)
);

BUFx4f_ASAP7_75t_L g2787 ( 
.A(n_2392),
.Y(n_2787)
);

INVxp67_ASAP7_75t_L g2788 ( 
.A(n_2456),
.Y(n_2788)
);

INVx3_ASAP7_75t_L g2789 ( 
.A(n_2340),
.Y(n_2789)
);

INVxp67_ASAP7_75t_L g2790 ( 
.A(n_2633),
.Y(n_2790)
);

AND2x4_ASAP7_75t_L g2791 ( 
.A(n_2494),
.B(n_1750),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2636),
.B(n_2178),
.Y(n_2792)
);

BUFx2_ASAP7_75t_L g2793 ( 
.A(n_2435),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2433),
.B(n_1750),
.Y(n_2794)
);

BUFx6f_ASAP7_75t_L g2795 ( 
.A(n_2357),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2579),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2344),
.Y(n_2797)
);

INVx5_ASAP7_75t_L g2798 ( 
.A(n_2515),
.Y(n_2798)
);

INVx4_ASAP7_75t_L g2799 ( 
.A(n_2316),
.Y(n_2799)
);

INVx4_ASAP7_75t_L g2800 ( 
.A(n_2378),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2494),
.B(n_1752),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2435),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2583),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2344),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2373),
.B(n_1752),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2653),
.B(n_1755),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2536),
.B(n_1755),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2357),
.Y(n_2808)
);

BUFx3_ASAP7_75t_L g2809 ( 
.A(n_2407),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2362),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2373),
.B(n_1761),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2439),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2354),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2598),
.B(n_1761),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2583),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2585),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2585),
.Y(n_2817)
);

HB1xp67_ASAP7_75t_L g2818 ( 
.A(n_2439),
.Y(n_2818)
);

NAND2xp33_ASAP7_75t_L g2819 ( 
.A(n_2515),
.B(n_1703),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2354),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2599),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2356),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2599),
.Y(n_2823)
);

INVxp33_ASAP7_75t_SL g2824 ( 
.A(n_2391),
.Y(n_2824)
);

HB1xp67_ASAP7_75t_L g2825 ( 
.A(n_2425),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2362),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2600),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2356),
.Y(n_2828)
);

INVx5_ASAP7_75t_L g2829 ( 
.A(n_2362),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2636),
.B(n_1778),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2600),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2590),
.B(n_2322),
.Y(n_2832)
);

INVxp67_ASAP7_75t_L g2833 ( 
.A(n_2633),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2592),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2352),
.B(n_1767),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2592),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2489),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2355),
.B(n_2594),
.Y(n_2838)
);

OR2x2_ASAP7_75t_SL g2839 ( 
.A(n_2440),
.B(n_2529),
.Y(n_2839)
);

BUFx3_ASAP7_75t_L g2840 ( 
.A(n_2463),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_2405),
.B(n_1778),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2490),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2464),
.B(n_1780),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2362),
.Y(n_2844)
);

BUFx6f_ASAP7_75t_L g2845 ( 
.A(n_2412),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2496),
.Y(n_2846)
);

AND2x6_ASAP7_75t_L g2847 ( 
.A(n_2620),
.B(n_1780),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2368),
.Y(n_2848)
);

INVx6_ASAP7_75t_L g2849 ( 
.A(n_2476),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_2463),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2368),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2500),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2412),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_2545),
.B(n_2520),
.Y(n_2854)
);

INVx3_ASAP7_75t_L g2855 ( 
.A(n_2412),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2502),
.Y(n_2856)
);

NAND2x1p5_ASAP7_75t_L g2857 ( 
.A(n_2525),
.B(n_1748),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2510),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2653),
.B(n_1767),
.Y(n_2859)
);

OAI221xp5_ASAP7_75t_L g2860 ( 
.A1(n_2530),
.A2(n_1768),
.B1(n_1780),
.B2(n_1706),
.C(n_1707),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2512),
.Y(n_2861)
);

AO22x2_ASAP7_75t_L g2862 ( 
.A1(n_2610),
.A2(n_1768),
.B1(n_84),
.B2(n_82),
.Y(n_2862)
);

INVx4_ASAP7_75t_L g2863 ( 
.A(n_2525),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2516),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2521),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2524),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2398),
.B(n_1780),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2370),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_SL g2869 ( 
.A(n_2534),
.B(n_2527),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2486),
.Y(n_2870)
);

BUFx3_ASAP7_75t_L g2871 ( 
.A(n_2431),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2528),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2429),
.B(n_1703),
.Y(n_2873)
);

AND2x4_ASAP7_75t_L g2874 ( 
.A(n_2429),
.B(n_1703),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2533),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2564),
.B(n_1703),
.Y(n_2876)
);

BUFx6f_ASAP7_75t_L g2877 ( 
.A(n_2412),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2537),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2543),
.Y(n_2879)
);

BUFx6f_ASAP7_75t_L g2880 ( 
.A(n_2418),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2548),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2503),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2591),
.B(n_83),
.Y(n_2883)
);

AND2x4_ASAP7_75t_L g2884 ( 
.A(n_2403),
.B(n_1705),
.Y(n_2884)
);

OR2x2_ASAP7_75t_L g2885 ( 
.A(n_2483),
.B(n_83),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2370),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2464),
.B(n_2345),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2398),
.B(n_1705),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2400),
.B(n_1705),
.Y(n_2889)
);

AND2x4_ASAP7_75t_L g2890 ( 
.A(n_2403),
.B(n_1705),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2374),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2564),
.B(n_1706),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2374),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2503),
.Y(n_2894)
);

BUFx2_ASAP7_75t_L g2895 ( 
.A(n_2486),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2505),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2418),
.Y(n_2897)
);

AND2x4_ASAP7_75t_L g2898 ( 
.A(n_2403),
.B(n_1706),
.Y(n_2898)
);

AND2x4_ASAP7_75t_L g2899 ( 
.A(n_2314),
.B(n_1706),
.Y(n_2899)
);

BUFx3_ASAP7_75t_L g2900 ( 
.A(n_2431),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2345),
.B(n_1707),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2591),
.B(n_84),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2379),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2379),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2346),
.B(n_1707),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2390),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2346),
.B(n_1707),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2505),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2390),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2469),
.B(n_1711),
.Y(n_2910)
);

INVx3_ASAP7_75t_L g2911 ( 
.A(n_2418),
.Y(n_2911)
);

INVx2_ASAP7_75t_SL g2912 ( 
.A(n_2506),
.Y(n_2912)
);

NAND3x1_ASAP7_75t_L g2913 ( 
.A(n_2648),
.B(n_86),
.C(n_85),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2530),
.A2(n_1711),
.B1(n_86),
.B2(n_84),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2400),
.B(n_1711),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2383),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2408),
.B(n_1711),
.Y(n_2917)
);

NAND2x1p5_ASAP7_75t_L g2918 ( 
.A(n_2469),
.B(n_85),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_2617),
.B(n_132),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2408),
.B(n_85),
.Y(n_2920)
);

AOI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2629),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2507),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_L g2923 ( 
.A(n_2418),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2507),
.Y(n_2924)
);

INVx5_ASAP7_75t_L g2925 ( 
.A(n_2476),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2535),
.Y(n_2926)
);

NAND2x1p5_ASAP7_75t_L g2927 ( 
.A(n_2479),
.B(n_2482),
.Y(n_2927)
);

AND2x6_ASAP7_75t_L g2928 ( 
.A(n_2648),
.B(n_87),
.Y(n_2928)
);

CKINVDCx5p33_ASAP7_75t_R g2929 ( 
.A(n_2383),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2531),
.Y(n_2930)
);

BUFx2_ASAP7_75t_L g2931 ( 
.A(n_2518),
.Y(n_2931)
);

INVx4_ASAP7_75t_L g2932 ( 
.A(n_2476),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2535),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2557),
.Y(n_2934)
);

AO22x2_ASAP7_75t_L g2935 ( 
.A1(n_2637),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_2935)
);

INVx5_ASAP7_75t_L g2936 ( 
.A(n_2606),
.Y(n_2936)
);

NAND3x1_ASAP7_75t_L g2937 ( 
.A(n_2639),
.B(n_90),
.C(n_89),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2557),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2508),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2559),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2559),
.Y(n_2941)
);

INVx3_ASAP7_75t_L g2942 ( 
.A(n_2453),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2453),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2621),
.B(n_88),
.Y(n_2944)
);

AND2x4_ASAP7_75t_L g2945 ( 
.A(n_2329),
.B(n_89),
.Y(n_2945)
);

NAND3xp33_ASAP7_75t_L g2946 ( 
.A(n_2311),
.B(n_135),
.C(n_134),
.Y(n_2946)
);

BUFx2_ASAP7_75t_L g2947 ( 
.A(n_2518),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2623),
.B(n_2307),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2428),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2428),
.Y(n_2950)
);

NAND3xp33_ASAP7_75t_L g2951 ( 
.A(n_2639),
.B(n_135),
.C(n_134),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2531),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2560),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2591),
.B(n_90),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2664),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2720),
.B(n_2654),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2667),
.Y(n_2957)
);

NAND3xp33_ASAP7_75t_SL g2958 ( 
.A(n_2692),
.B(n_2607),
.C(n_2544),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2672),
.Y(n_2959)
);

A2O1A1Ixp33_ASAP7_75t_L g2960 ( 
.A1(n_2665),
.A2(n_2570),
.B(n_2601),
.C(n_2339),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2720),
.B(n_2578),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2676),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2724),
.B(n_2437),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2673),
.Y(n_2964)
);

O2A1O1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2665),
.A2(n_2546),
.B(n_2449),
.C(n_2605),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2724),
.B(n_2437),
.Y(n_2966)
);

INVxp33_ASAP7_75t_L g2967 ( 
.A(n_2662),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2832),
.B(n_2438),
.Y(n_2968)
);

INVx3_ASAP7_75t_L g2969 ( 
.A(n_2798),
.Y(n_2969)
);

NOR3xp33_ASAP7_75t_L g2970 ( 
.A(n_2692),
.B(n_2449),
.C(n_2605),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2679),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2681),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2668),
.B(n_2854),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2832),
.B(n_2838),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_SL g2975 ( 
.A(n_2869),
.B(n_2556),
.Y(n_2975)
);

AOI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2819),
.A2(n_2343),
.B(n_2315),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2838),
.B(n_2450),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2705),
.B(n_2593),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_SL g2979 ( 
.A(n_2788),
.B(n_2556),
.Y(n_2979)
);

AND2x4_ASAP7_75t_L g2980 ( 
.A(n_2674),
.B(n_2540),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2790),
.B(n_2438),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2705),
.B(n_2655),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2824),
.B(n_2518),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_2721),
.B(n_2309),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2684),
.A2(n_2458),
.B1(n_2661),
.B2(n_2563),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2678),
.Y(n_2986)
);

BUFx3_ASAP7_75t_L g2987 ( 
.A(n_2712),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2685),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2788),
.B(n_2618),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2682),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2697),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2703),
.Y(n_2992)
);

BUFx6f_ASAP7_75t_SL g2993 ( 
.A(n_2809),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2723),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2798),
.B(n_2618),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2721),
.B(n_2582),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2710),
.B(n_2328),
.Y(n_2997)
);

NOR2x1p5_ASAP7_75t_L g2998 ( 
.A(n_2871),
.B(n_2442),
.Y(n_2998)
);

BUFx6f_ASAP7_75t_L g2999 ( 
.A(n_2737),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2708),
.B(n_2389),
.Y(n_3000)
);

AND2x4_ASAP7_75t_SL g3001 ( 
.A(n_2691),
.B(n_2392),
.Y(n_3001)
);

HB1xp67_ASAP7_75t_L g3002 ( 
.A(n_2698),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2698),
.B(n_2328),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2669),
.B(n_2385),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2725),
.Y(n_3005)
);

HB1xp67_ASAP7_75t_L g3006 ( 
.A(n_2753),
.Y(n_3006)
);

AND2x2_ASAP7_75t_SL g3007 ( 
.A(n_2787),
.B(n_2616),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2755),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2690),
.Y(n_3009)
);

O2A1O1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2718),
.A2(n_2555),
.B(n_2315),
.C(n_2475),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2756),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2693),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2686),
.B(n_2389),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2715),
.B(n_2634),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_SL g3015 ( 
.A1(n_2684),
.A2(n_2615),
.B1(n_2632),
.B2(n_2640),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2694),
.Y(n_3016)
);

INVx8_ASAP7_75t_L g3017 ( 
.A(n_2737),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2790),
.B(n_2833),
.Y(n_3018)
);

AOI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2684),
.A2(n_2581),
.B1(n_2649),
.B2(n_2616),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2669),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2701),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2757),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2798),
.B(n_2618),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2736),
.B(n_2385),
.Y(n_3024)
);

NAND2xp33_ASAP7_75t_L g3025 ( 
.A(n_2731),
.B(n_2453),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_2900),
.B(n_2655),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2753),
.B(n_2392),
.Y(n_3027)
);

NOR2x1p5_ASAP7_75t_L g3028 ( 
.A(n_2767),
.B(n_2649),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_SL g3029 ( 
.A1(n_2773),
.A2(n_2624),
.B1(n_2628),
.B2(n_2626),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2758),
.Y(n_3030)
);

NOR2xp67_ASAP7_75t_L g3031 ( 
.A(n_2785),
.B(n_2493),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_2930),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2728),
.B(n_2647),
.Y(n_3033)
);

INVxp67_ASAP7_75t_SL g3034 ( 
.A(n_2677),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2759),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2737),
.Y(n_3036)
);

OR2x2_ASAP7_75t_L g3037 ( 
.A(n_2736),
.B(n_2717),
.Y(n_3037)
);

AO221x1_ASAP7_75t_L g3038 ( 
.A1(n_2935),
.A2(n_2401),
.B1(n_2596),
.B2(n_2660),
.C(n_2421),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2732),
.B(n_2613),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2702),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2704),
.Y(n_3041)
);

NOR2xp33_ASAP7_75t_L g3042 ( 
.A(n_2887),
.B(n_2509),
.Y(n_3042)
);

AOI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_2689),
.A2(n_2608),
.B1(n_2627),
.B2(n_2601),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2762),
.Y(n_3044)
);

O2A1O1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_2680),
.A2(n_2472),
.B(n_2511),
.C(n_2480),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_SL g3046 ( 
.A(n_2798),
.B(n_2631),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2883),
.B(n_2613),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2818),
.B(n_2509),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2833),
.B(n_2470),
.Y(n_3049)
);

A2O1A1Ixp33_ASAP7_75t_L g3050 ( 
.A1(n_2689),
.A2(n_2570),
.B(n_2658),
.C(n_2462),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2948),
.B(n_2470),
.Y(n_3051)
);

OAI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2914),
.A2(n_2402),
.B1(n_2413),
.B2(n_2387),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2779),
.B(n_2561),
.Y(n_3053)
);

AOI22xp33_ASAP7_75t_L g3054 ( 
.A1(n_2773),
.A2(n_2581),
.B1(n_2575),
.B2(n_2641),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2765),
.Y(n_3055)
);

INVx3_ASAP7_75t_L g3056 ( 
.A(n_2754),
.Y(n_3056)
);

INVx3_ASAP7_75t_L g3057 ( 
.A(n_2754),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2706),
.Y(n_3058)
);

INVx4_ASAP7_75t_L g3059 ( 
.A(n_2829),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2869),
.B(n_2948),
.Y(n_3060)
);

AND2x4_ASAP7_75t_L g3061 ( 
.A(n_2674),
.B(n_2553),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2919),
.B(n_2695),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2677),
.B(n_2471),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2782),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2695),
.B(n_2387),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2797),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_2818),
.B(n_2841),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2804),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2735),
.B(n_2471),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2747),
.B(n_2509),
.Y(n_3070)
);

OAI22xp5_ASAP7_75t_L g3071 ( 
.A1(n_2914),
.A2(n_2402),
.B1(n_2417),
.B2(n_2413),
.Y(n_3071)
);

NOR2xp67_ASAP7_75t_L g3072 ( 
.A(n_2687),
.B(n_2538),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2939),
.B(n_2353),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2944),
.B(n_2417),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2813),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2709),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2820),
.Y(n_3077)
);

INVx8_ASAP7_75t_L g3078 ( 
.A(n_2754),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2735),
.B(n_2478),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2822),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2711),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2746),
.B(n_2478),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2746),
.B(n_2307),
.Y(n_3083)
);

BUFx3_ASAP7_75t_L g3084 ( 
.A(n_2840),
.Y(n_3084)
);

A2O1A1Ixp33_ASAP7_75t_L g3085 ( 
.A1(n_2951),
.A2(n_2658),
.B(n_2452),
.C(n_2646),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_2952),
.Y(n_3086)
);

NOR2xp67_ASAP7_75t_L g3087 ( 
.A(n_2766),
.B(n_2538),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2713),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2714),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_2740),
.A2(n_2602),
.B1(n_2401),
.B2(n_2587),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2944),
.B(n_2488),
.Y(n_3091)
);

NAND2x1_ASAP7_75t_L g3092 ( 
.A(n_2844),
.B(n_2333),
.Y(n_3092)
);

NAND2x1_ASAP7_75t_L g3093 ( 
.A(n_2844),
.B(n_2333),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2716),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_SL g3095 ( 
.A(n_2925),
.B(n_2349),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_SL g3096 ( 
.A(n_2925),
.B(n_2800),
.Y(n_3096)
);

NOR2xp67_ASAP7_75t_SL g3097 ( 
.A(n_2929),
.B(n_2538),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2825),
.B(n_2584),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2939),
.B(n_2353),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_2764),
.B(n_2353),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2675),
.B(n_2421),
.Y(n_3101)
);

INVx3_ASAP7_75t_L g3102 ( 
.A(n_2777),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2675),
.B(n_2421),
.Y(n_3103)
);

NOR3x1_ASAP7_75t_L g3104 ( 
.A(n_2730),
.B(n_2514),
.C(n_2573),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2696),
.B(n_2468),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2696),
.B(n_2484),
.Y(n_3106)
);

AND2x6_ASAP7_75t_SL g3107 ( 
.A(n_2739),
.B(n_2364),
.Y(n_3107)
);

AND2x6_ASAP7_75t_SL g3108 ( 
.A(n_2683),
.B(n_2364),
.Y(n_3108)
);

INVx3_ASAP7_75t_L g3109 ( 
.A(n_2777),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2828),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2726),
.Y(n_3111)
);

O2A1O1Ixp5_ASAP7_75t_L g3112 ( 
.A1(n_2719),
.A2(n_2611),
.B(n_2342),
.C(n_2334),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2925),
.B(n_2569),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2805),
.B(n_2606),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2902),
.B(n_2954),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2805),
.B(n_2811),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_2763),
.B(n_2364),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2811),
.B(n_2606),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2843),
.B(n_2769),
.Y(n_3119)
);

AOI22xp5_ASAP7_75t_L g3120 ( 
.A1(n_2764),
.A2(n_2608),
.B1(n_2638),
.B2(n_2554),
.Y(n_3120)
);

INVx2_ASAP7_75t_SL g3121 ( 
.A(n_2787),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_2683),
.A2(n_2614),
.B1(n_2445),
.B2(n_2606),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2843),
.B(n_2769),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2727),
.B(n_2606),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2848),
.Y(n_3125)
);

BUFx12f_ASAP7_75t_L g3126 ( 
.A(n_2839),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2727),
.B(n_2560),
.Y(n_3127)
);

BUFx6f_ASAP7_75t_L g3128 ( 
.A(n_2742),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2733),
.A2(n_2609),
.B1(n_2562),
.B2(n_2611),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2734),
.Y(n_3130)
);

BUFx3_ASAP7_75t_L g3131 ( 
.A(n_2850),
.Y(n_3131)
);

AOI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_2928),
.A2(n_2609),
.B1(n_2625),
.B2(n_2622),
.Y(n_3132)
);

BUFx6f_ASAP7_75t_L g3133 ( 
.A(n_2742),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2851),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2812),
.B(n_2406),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2925),
.B(n_2569),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2742),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2868),
.Y(n_3138)
);

O2A1O1Ixp33_ASAP7_75t_L g3139 ( 
.A1(n_2730),
.A2(n_2343),
.B(n_2434),
.C(n_2573),
.Y(n_3139)
);

OAI22xp5_ASAP7_75t_SL g3140 ( 
.A1(n_2683),
.A2(n_2921),
.B1(n_2951),
.B2(n_2946),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2738),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2886),
.Y(n_3142)
);

CKINVDCx5p33_ASAP7_75t_R g3143 ( 
.A(n_2916),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2670),
.B(n_2436),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2774),
.B(n_2436),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2780),
.B(n_2497),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2825),
.B(n_2497),
.Y(n_3147)
);

INVx2_ASAP7_75t_SL g3148 ( 
.A(n_2783),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2794),
.B(n_2474),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2781),
.B(n_2796),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2803),
.B(n_2586),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_SL g3152 ( 
.A(n_2800),
.B(n_2569),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2815),
.B(n_2446),
.Y(n_3153)
);

A2O1A1Ixp33_ASAP7_75t_SL g3154 ( 
.A1(n_2901),
.A2(n_2434),
.B(n_2646),
.C(n_2643),
.Y(n_3154)
);

AOI22xp5_ASAP7_75t_L g3155 ( 
.A1(n_2928),
.A2(n_2609),
.B1(n_2522),
.B2(n_2595),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_SL g3156 ( 
.A(n_2936),
.B(n_2569),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2870),
.B(n_2614),
.Y(n_3157)
);

INVxp67_ASAP7_75t_L g3158 ( 
.A(n_2663),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2816),
.B(n_2831),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2817),
.B(n_2430),
.Y(n_3160)
);

NAND3xp33_ASAP7_75t_L g3161 ( 
.A(n_2946),
.B(n_2643),
.C(n_2517),
.Y(n_3161)
);

OAI22xp5_ASAP7_75t_L g3162 ( 
.A1(n_2860),
.A2(n_2448),
.B1(n_2451),
.B2(n_2447),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2888),
.A2(n_2324),
.B(n_2342),
.Y(n_3163)
);

BUFx6f_ASAP7_75t_L g3164 ( 
.A(n_2829),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2936),
.B(n_2453),
.Y(n_3165)
);

INVxp67_ASAP7_75t_L g3166 ( 
.A(n_2885),
.Y(n_3166)
);

INVx1_ASAP7_75t_SL g3167 ( 
.A(n_2895),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2821),
.B(n_2542),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2837),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2823),
.B(n_2542),
.Y(n_3170)
);

OR2x6_ASAP7_75t_L g3171 ( 
.A(n_2777),
.B(n_2522),
.Y(n_3171)
);

NOR2xp33_ASAP7_75t_L g3172 ( 
.A(n_2931),
.B(n_2504),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_2936),
.B(n_2473),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_2888),
.A2(n_2324),
.B(n_2487),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2827),
.B(n_2547),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2891),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2889),
.A2(n_2492),
.B(n_2487),
.Y(n_3177)
);

AOI22xp5_ASAP7_75t_L g3178 ( 
.A1(n_2928),
.A2(n_2937),
.B1(n_2775),
.B2(n_2792),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_3000),
.B(n_2945),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2974),
.B(n_2750),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2972),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2955),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_2980),
.B(n_2936),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_2987),
.Y(n_3184)
);

OAI21xp33_ASAP7_75t_SL g3185 ( 
.A1(n_2977),
.A2(n_2860),
.B(n_2920),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2957),
.Y(n_3186)
);

INVx4_ASAP7_75t_L g3187 ( 
.A(n_3017),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2974),
.B(n_2772),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3119),
.B(n_2744),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2959),
.Y(n_3190)
);

AO22x1_ASAP7_75t_L g3191 ( 
.A1(n_3014),
.A2(n_2928),
.B1(n_2912),
.B2(n_2688),
.Y(n_3191)
);

BUFx2_ASAP7_75t_L g3192 ( 
.A(n_2973),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_3164),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_2980),
.B(n_2674),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2962),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_3119),
.B(n_2749),
.Y(n_3196)
);

BUFx2_ASAP7_75t_L g3197 ( 
.A(n_3027),
.Y(n_3197)
);

NAND2x1p5_ASAP7_75t_L g3198 ( 
.A(n_2969),
.B(n_2829),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_3006),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2990),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2986),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2988),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3009),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3012),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3016),
.Y(n_3205)
);

HB1xp67_ASAP7_75t_L g3206 ( 
.A(n_3002),
.Y(n_3206)
);

AOI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_2997),
.A2(n_3140),
.B1(n_2970),
.B2(n_2935),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3123),
.B(n_2893),
.Y(n_3208)
);

BUFx6f_ASAP7_75t_L g3209 ( 
.A(n_3164),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3021),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_3010),
.B(n_2830),
.Y(n_3211)
);

BUFx3_ASAP7_75t_L g3212 ( 
.A(n_3084),
.Y(n_3212)
);

AOI22xp33_ASAP7_75t_L g3213 ( 
.A1(n_3038),
.A2(n_2862),
.B1(n_2935),
.B2(n_2700),
.Y(n_3213)
);

HB1xp67_ASAP7_75t_L g3214 ( 
.A(n_3067),
.Y(n_3214)
);

BUFx6f_ASAP7_75t_L g3215 ( 
.A(n_3164),
.Y(n_3215)
);

CKINVDCx8_ASAP7_75t_R g3216 ( 
.A(n_3107),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3040),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_2982),
.B(n_2945),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2991),
.Y(n_3219)
);

AOI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_3043),
.A2(n_2862),
.B1(n_2913),
.B2(n_2671),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2956),
.B(n_2947),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2992),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_2978),
.B(n_2862),
.Y(n_3223)
);

INVx5_ASAP7_75t_L g3224 ( 
.A(n_3078),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_3018),
.Y(n_3225)
);

NOR2xp33_ASAP7_75t_L g3226 ( 
.A(n_2984),
.B(n_2784),
.Y(n_3226)
);

BUFx2_ASAP7_75t_L g3227 ( 
.A(n_3143),
.Y(n_3227)
);

INVx2_ASAP7_75t_SL g3228 ( 
.A(n_3131),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3123),
.B(n_2903),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_3032),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2968),
.B(n_2904),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3041),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_2967),
.B(n_3018),
.Y(n_3233)
);

HB1xp67_ASAP7_75t_L g3234 ( 
.A(n_3048),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_L g3235 ( 
.A1(n_2958),
.A2(n_2770),
.B1(n_2513),
.B2(n_2671),
.Y(n_3235)
);

INVx4_ASAP7_75t_L g3236 ( 
.A(n_3017),
.Y(n_3236)
);

CKINVDCx5p33_ASAP7_75t_R g3237 ( 
.A(n_3086),
.Y(n_3237)
);

INVx4_ASAP7_75t_L g3238 ( 
.A(n_3017),
.Y(n_3238)
);

INVx5_ASAP7_75t_L g3239 ( 
.A(n_3078),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_3042),
.A2(n_2671),
.B1(n_2666),
.B2(n_2834),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3053),
.B(n_2784),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_3059),
.Y(n_3242)
);

INVx2_ASAP7_75t_SL g3243 ( 
.A(n_3001),
.Y(n_3243)
);

AND2x2_ASAP7_75t_SL g3244 ( 
.A(n_3007),
.B(n_2975),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3169),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3058),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2994),
.Y(n_3247)
);

CKINVDCx5p33_ASAP7_75t_R g3248 ( 
.A(n_2993),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_3059),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3005),
.Y(n_3250)
);

CKINVDCx16_ASAP7_75t_R g3251 ( 
.A(n_2993),
.Y(n_3251)
);

INVx5_ASAP7_75t_L g3252 ( 
.A(n_3078),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_3020),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3076),
.Y(n_3254)
);

BUFx12f_ASAP7_75t_L g3255 ( 
.A(n_3126),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2968),
.B(n_2906),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3081),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3088),
.Y(n_3258)
);

INVx1_ASAP7_75t_SL g3259 ( 
.A(n_3167),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3089),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2956),
.B(n_2909),
.Y(n_3261)
);

INVx2_ASAP7_75t_SL g3262 ( 
.A(n_2998),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3105),
.B(n_2949),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3094),
.Y(n_3264)
);

OR2x2_ASAP7_75t_SL g3265 ( 
.A(n_3062),
.B(n_2849),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_3115),
.B(n_2806),
.Y(n_3266)
);

HB1xp67_ASAP7_75t_L g3267 ( 
.A(n_3098),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3105),
.B(n_2950),
.Y(n_3268)
);

AOI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_2989),
.A2(n_2671),
.B1(n_2666),
.B2(n_2836),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_SL g3270 ( 
.A(n_3060),
.B(n_2829),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3091),
.B(n_2748),
.Y(n_3271)
);

OAI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_3120),
.A2(n_2918),
.B1(n_2920),
.B2(n_2835),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3178),
.A2(n_2666),
.B1(n_2847),
.B2(n_2778),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3149),
.B(n_2793),
.Y(n_3274)
);

INVx4_ASAP7_75t_L g3275 ( 
.A(n_2999),
.Y(n_3275)
);

INVx4_ASAP7_75t_L g3276 ( 
.A(n_2999),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_3117),
.Y(n_3277)
);

INVx6_ASAP7_75t_L g3278 ( 
.A(n_3028),
.Y(n_3278)
);

BUFx6f_ASAP7_75t_L g3279 ( 
.A(n_2999),
.Y(n_3279)
);

BUFx4f_ASAP7_75t_L g3280 ( 
.A(n_3036),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3106),
.B(n_2731),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_2964),
.Y(n_3282)
);

BUFx12f_ASAP7_75t_L g3283 ( 
.A(n_3148),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3106),
.B(n_2731),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3111),
.Y(n_3285)
);

CKINVDCx5p33_ASAP7_75t_R g3286 ( 
.A(n_2996),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3116),
.B(n_2731),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2971),
.Y(n_3288)
);

AND2x4_ASAP7_75t_L g3289 ( 
.A(n_3061),
.B(n_2802),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3116),
.B(n_2771),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3051),
.B(n_2771),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_3036),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3130),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3051),
.B(n_2771),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3141),
.Y(n_3295)
);

BUFx12f_ASAP7_75t_L g3296 ( 
.A(n_3121),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3008),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_2983),
.B(n_3013),
.Y(n_3298)
);

INVx2_ASAP7_75t_SL g3299 ( 
.A(n_3128),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2963),
.B(n_2771),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3047),
.B(n_2859),
.Y(n_3301)
);

INVx5_ASAP7_75t_L g3302 ( 
.A(n_3171),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3011),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3022),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3030),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3035),
.Y(n_3306)
);

INVx3_ASAP7_75t_L g3307 ( 
.A(n_3036),
.Y(n_3307)
);

BUFx2_ASAP7_75t_L g3308 ( 
.A(n_3128),
.Y(n_3308)
);

INVx2_ASAP7_75t_SL g3309 ( 
.A(n_3128),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2963),
.B(n_2666),
.Y(n_3310)
);

BUFx3_ASAP7_75t_L g3311 ( 
.A(n_3135),
.Y(n_3311)
);

BUFx6f_ASAP7_75t_L g3312 ( 
.A(n_3133),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3044),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2966),
.B(n_2814),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3055),
.Y(n_3315)
);

BUFx8_ASAP7_75t_L g3316 ( 
.A(n_3133),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_3052),
.A2(n_2770),
.B1(n_2513),
.B2(n_2842),
.Y(n_3317)
);

BUFx3_ASAP7_75t_L g3318 ( 
.A(n_3026),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3064),
.Y(n_3319)
);

INVx4_ASAP7_75t_L g3320 ( 
.A(n_3133),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3066),
.Y(n_3321)
);

BUFx12f_ASAP7_75t_L g3322 ( 
.A(n_3137),
.Y(n_3322)
);

BUFx4f_ASAP7_75t_L g3323 ( 
.A(n_3137),
.Y(n_3323)
);

AND2x4_ASAP7_75t_L g3324 ( 
.A(n_3061),
.B(n_2890),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3068),
.Y(n_3325)
);

BUFx4f_ASAP7_75t_L g3326 ( 
.A(n_3137),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_2966),
.B(n_2814),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3075),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_3073),
.B(n_2799),
.Y(n_3329)
);

BUFx6f_ASAP7_75t_L g3330 ( 
.A(n_3056),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3077),
.Y(n_3331)
);

BUFx3_ASAP7_75t_L g3332 ( 
.A(n_3172),
.Y(n_3332)
);

AND3x2_ASAP7_75t_SL g3333 ( 
.A(n_3108),
.B(n_2770),
.C(n_2918),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3080),
.Y(n_3334)
);

HB1xp67_ASAP7_75t_L g3335 ( 
.A(n_3147),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3110),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3125),
.Y(n_3337)
);

AND2x4_ASAP7_75t_L g3338 ( 
.A(n_3171),
.B(n_2884),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_2981),
.B(n_2847),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2981),
.B(n_2847),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3049),
.B(n_2847),
.Y(n_3341)
);

BUFx2_ASAP7_75t_L g3342 ( 
.A(n_3099),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3134),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3138),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3049),
.B(n_2882),
.Y(n_3345)
);

AND2x4_ASAP7_75t_L g3346 ( 
.A(n_3171),
.B(n_2884),
.Y(n_3346)
);

BUFx2_ASAP7_75t_L g3347 ( 
.A(n_3166),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3142),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2961),
.B(n_3082),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3176),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3159),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3159),
.Y(n_3352)
);

AND2x4_ASAP7_75t_L g3353 ( 
.A(n_3056),
.B(n_2898),
.Y(n_3353)
);

CKINVDCx5p33_ASAP7_75t_R g3354 ( 
.A(n_2979),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3150),
.Y(n_3355)
);

BUFx3_ASAP7_75t_L g3356 ( 
.A(n_3037),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_2976),
.A2(n_2334),
.B(n_2335),
.Y(n_3357)
);

INVx1_ASAP7_75t_SL g3358 ( 
.A(n_3065),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3160),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_3070),
.B(n_2799),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2961),
.B(n_2894),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3168),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3004),
.B(n_2846),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3039),
.B(n_2707),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3024),
.B(n_2852),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3168),
.Y(n_3366)
);

BUFx3_ASAP7_75t_L g3367 ( 
.A(n_3057),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_3100),
.B(n_2863),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_3170),
.Y(n_3369)
);

OR2x2_ASAP7_75t_L g3370 ( 
.A(n_3033),
.B(n_2856),
.Y(n_3370)
);

BUFx6f_ASAP7_75t_L g3371 ( 
.A(n_3057),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3170),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3175),
.Y(n_3373)
);

NOR2xp33_ASAP7_75t_L g3374 ( 
.A(n_3144),
.B(n_2863),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_3102),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3175),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3145),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3158),
.B(n_2745),
.Y(n_3378)
);

BUFx3_ASAP7_75t_L g3379 ( 
.A(n_3102),
.Y(n_3379)
);

BUFx4f_ASAP7_75t_SL g3380 ( 
.A(n_2995),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3003),
.B(n_2858),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3145),
.Y(n_3382)
);

INVx1_ASAP7_75t_SL g3383 ( 
.A(n_3023),
.Y(n_3383)
);

AND2x4_ASAP7_75t_L g3384 ( 
.A(n_3109),
.B(n_2898),
.Y(n_3384)
);

BUFx6f_ASAP7_75t_L g3385 ( 
.A(n_3109),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_3146),
.Y(n_3386)
);

BUFx3_ASAP7_75t_L g3387 ( 
.A(n_2969),
.Y(n_3387)
);

INVx3_ASAP7_75t_L g3388 ( 
.A(n_3092),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_3214),
.B(n_2745),
.Y(n_3389)
);

A2O1A1Ixp33_ASAP7_75t_L g3390 ( 
.A1(n_3185),
.A2(n_2965),
.B(n_3139),
.C(n_3085),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3225),
.B(n_3074),
.Y(n_3391)
);

INVx4_ASAP7_75t_L g3392 ( 
.A(n_3322),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3267),
.B(n_3114),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3185),
.A2(n_3162),
.B(n_3034),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3286),
.B(n_3226),
.Y(n_3395)
);

BUFx4f_ASAP7_75t_L g3396 ( 
.A(n_3255),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3182),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3282),
.Y(n_3398)
);

OAI21x1_ASAP7_75t_L g3399 ( 
.A1(n_3357),
.A2(n_3163),
.B(n_3112),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3288),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3211),
.A2(n_3162),
.B(n_3025),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3314),
.A2(n_2960),
.B(n_3050),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3186),
.Y(n_3403)
);

BUFx4f_ASAP7_75t_L g3404 ( 
.A(n_3279),
.Y(n_3404)
);

BUFx4f_ASAP7_75t_L g3405 ( 
.A(n_3279),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3297),
.Y(n_3406)
);

OAI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_3272),
.A2(n_3045),
.B(n_3161),
.Y(n_3407)
);

OAI21x1_ASAP7_75t_L g3408 ( 
.A1(n_3272),
.A2(n_3174),
.B(n_3177),
.Y(n_3408)
);

CKINVDCx20_ASAP7_75t_R g3409 ( 
.A(n_3251),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3190),
.Y(n_3410)
);

OAI21xp33_ASAP7_75t_SL g3411 ( 
.A1(n_3220),
.A2(n_3046),
.B(n_3122),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3314),
.A2(n_3069),
.B(n_3063),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3335),
.B(n_3234),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3207),
.A2(n_3220),
.B1(n_3241),
.B2(n_3374),
.Y(n_3414)
);

INVx3_ASAP7_75t_L g3415 ( 
.A(n_3193),
.Y(n_3415)
);

OA22x2_ASAP7_75t_L g3416 ( 
.A1(n_3207),
.A2(n_3223),
.B1(n_3240),
.B2(n_3273),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3305),
.Y(n_3417)
);

XNOR2xp5_ASAP7_75t_L g3418 ( 
.A(n_3230),
.B(n_3031),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3192),
.B(n_3114),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3327),
.A2(n_3069),
.B(n_3063),
.Y(n_3420)
);

OAI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3378),
.A2(n_3129),
.B(n_3154),
.Y(n_3421)
);

BUFx6f_ASAP7_75t_L g3422 ( 
.A(n_3280),
.Y(n_3422)
);

OAI21x1_ASAP7_75t_L g3423 ( 
.A1(n_3388),
.A2(n_2519),
.B(n_3124),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3271),
.B(n_3118),
.Y(n_3424)
);

CKINVDCx20_ASAP7_75t_R g3425 ( 
.A(n_3237),
.Y(n_3425)
);

INVxp67_ASAP7_75t_L g3426 ( 
.A(n_3253),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3359),
.B(n_3118),
.Y(n_3427)
);

O2A1O1Ixp33_ASAP7_75t_L g3428 ( 
.A1(n_3206),
.A2(n_3152),
.B(n_3096),
.C(n_3146),
.Y(n_3428)
);

A2O1A1Ixp33_ASAP7_75t_L g3429 ( 
.A1(n_3179),
.A2(n_3029),
.B(n_3071),
.C(n_3052),
.Y(n_3429)
);

OAI21x1_ASAP7_75t_L g3430 ( 
.A1(n_3388),
.A2(n_3124),
.B(n_2892),
.Y(n_3430)
);

A2O1A1Ixp33_ASAP7_75t_L g3431 ( 
.A1(n_3273),
.A2(n_3071),
.B(n_2985),
.C(n_3132),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3199),
.B(n_3104),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3195),
.Y(n_3433)
);

NAND2x1p5_ASAP7_75t_L g3434 ( 
.A(n_3224),
.B(n_3097),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_SL g3435 ( 
.A(n_3216),
.B(n_2932),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_3327),
.A2(n_3079),
.B(n_3156),
.Y(n_3436)
);

OAI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3354),
.A2(n_3155),
.B1(n_3090),
.B2(n_3054),
.Y(n_3437)
);

INVxp67_ASAP7_75t_L g3438 ( 
.A(n_3233),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_SL g3439 ( 
.A(n_3244),
.B(n_2932),
.Y(n_3439)
);

INVx4_ASAP7_75t_L g3440 ( 
.A(n_3224),
.Y(n_3440)
);

OAI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_3235),
.A2(n_2927),
.B1(n_3103),
.B2(n_3101),
.Y(n_3441)
);

OAI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3360),
.A2(n_3284),
.B(n_3281),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3218),
.B(n_3342),
.Y(n_3443)
);

BUFx6f_ASAP7_75t_L g3444 ( 
.A(n_3280),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_3287),
.A2(n_3079),
.B(n_2876),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3332),
.B(n_2789),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3221),
.B(n_3082),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3213),
.A2(n_2927),
.B1(n_3101),
.B2(n_3103),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3287),
.A2(n_3173),
.B(n_3165),
.Y(n_3449)
);

O2A1O1Ixp33_ASAP7_75t_L g3450 ( 
.A1(n_3259),
.A2(n_3095),
.B(n_3136),
.C(n_3113),
.Y(n_3450)
);

CKINVDCx20_ASAP7_75t_R g3451 ( 
.A(n_3248),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3370),
.B(n_3153),
.Y(n_3452)
);

INVx4_ASAP7_75t_L g3453 ( 
.A(n_3224),
.Y(n_3453)
);

NAND2x1_ASAP7_75t_L g3454 ( 
.A(n_3242),
.B(n_2855),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_3290),
.A2(n_3284),
.B(n_3281),
.Y(n_3455)
);

NOR2xp67_ASAP7_75t_SL g3456 ( 
.A(n_3239),
.B(n_2743),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_L g3457 ( 
.A(n_3298),
.B(n_2789),
.Y(n_3457)
);

INVxp67_ASAP7_75t_SL g3458 ( 
.A(n_3290),
.Y(n_3458)
);

BUFx6f_ASAP7_75t_L g3459 ( 
.A(n_3212),
.Y(n_3459)
);

CKINVDCx6p67_ASAP7_75t_R g3460 ( 
.A(n_3296),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3259),
.B(n_3358),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3339),
.A2(n_2335),
.B(n_2642),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_3380),
.B(n_3368),
.Y(n_3463)
);

AOI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_3266),
.A2(n_3157),
.B1(n_2778),
.B2(n_3019),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3313),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3364),
.B(n_3015),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3339),
.A2(n_2499),
.B(n_2492),
.Y(n_3467)
);

CKINVDCx10_ASAP7_75t_R g3468 ( 
.A(n_3262),
.Y(n_3468)
);

BUFx3_ASAP7_75t_L g3469 ( 
.A(n_3184),
.Y(n_3469)
);

OAI22xp5_ASAP7_75t_L g3470 ( 
.A1(n_3265),
.A2(n_2849),
.B1(n_2595),
.B2(n_2482),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3358),
.B(n_3153),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3340),
.A2(n_2501),
.B(n_2499),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3274),
.B(n_3127),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3227),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_3318),
.B(n_3072),
.Y(n_3475)
);

OAI21xp33_ASAP7_75t_L g3476 ( 
.A1(n_3317),
.A2(n_3349),
.B(n_3341),
.Y(n_3476)
);

INVx1_ASAP7_75t_SL g3477 ( 
.A(n_3311),
.Y(n_3477)
);

AOI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3340),
.A2(n_2501),
.B(n_2776),
.Y(n_3478)
);

BUFx6f_ASAP7_75t_L g3479 ( 
.A(n_3323),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3355),
.B(n_3127),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3351),
.B(n_3083),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3352),
.B(n_3083),
.Y(n_3482)
);

OAI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3341),
.A2(n_2907),
.B(n_2905),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3180),
.B(n_2861),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3240),
.A2(n_2849),
.B1(n_2595),
.B2(n_2479),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3315),
.Y(n_3486)
);

BUFx12f_ASAP7_75t_L g3487 ( 
.A(n_3316),
.Y(n_3487)
);

BUFx2_ASAP7_75t_SL g3488 ( 
.A(n_3228),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3329),
.B(n_136),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3300),
.A2(n_2776),
.B(n_2889),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_3193),
.B(n_3087),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3201),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3300),
.A2(n_2917),
.B(n_2915),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3180),
.B(n_2864),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3188),
.B(n_2865),
.Y(n_3495)
);

BUFx2_ASAP7_75t_L g3496 ( 
.A(n_3316),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3277),
.B(n_3197),
.Y(n_3497)
);

AOI21xp33_ASAP7_75t_L g3498 ( 
.A1(n_3363),
.A2(n_3151),
.B(n_2760),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3310),
.A2(n_2917),
.B(n_2915),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3188),
.B(n_2866),
.Y(n_3500)
);

CKINVDCx5p33_ASAP7_75t_R g3501 ( 
.A(n_3283),
.Y(n_3501)
);

O2A1O1Ixp33_ASAP7_75t_L g3502 ( 
.A1(n_3347),
.A2(n_2644),
.B(n_2645),
.C(n_2459),
.Y(n_3502)
);

INVx5_ASAP7_75t_L g3503 ( 
.A(n_3193),
.Y(n_3503)
);

AOI22xp5_ASAP7_75t_L g3504 ( 
.A1(n_3301),
.A2(n_2645),
.B1(n_2644),
.B2(n_2635),
.Y(n_3504)
);

AND2x4_ASAP7_75t_L g3505 ( 
.A(n_3356),
.B(n_3151),
.Y(n_3505)
);

OAI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3269),
.A2(n_2567),
.B1(n_2566),
.B2(n_2523),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3202),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3310),
.A2(n_3294),
.B(n_3291),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3349),
.B(n_2872),
.Y(n_3509)
);

INVxp67_ASAP7_75t_L g3510 ( 
.A(n_3308),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3203),
.Y(n_3511)
);

O2A1O1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3189),
.A2(n_2459),
.B(n_2835),
.C(n_2707),
.Y(n_3512)
);

OAI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_3291),
.A2(n_2699),
.B(n_2358),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3321),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3294),
.A2(n_2635),
.B(n_2752),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_SL g3516 ( 
.A(n_3187),
.B(n_2873),
.Y(n_3516)
);

AOI22x1_ASAP7_75t_L g3517 ( 
.A1(n_3187),
.A2(n_2743),
.B1(n_2943),
.B2(n_2942),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3204),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3189),
.B(n_2875),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3243),
.B(n_3307),
.Y(n_3520)
);

AO21x1_ASAP7_75t_L g3521 ( 
.A1(n_3196),
.A2(n_2358),
.B(n_2351),
.Y(n_3521)
);

AOI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_3269),
.A2(n_2873),
.B1(n_2874),
.B2(n_2619),
.Y(n_3522)
);

O2A1O1Ixp33_ASAP7_75t_L g3523 ( 
.A1(n_3196),
.A2(n_2351),
.B(n_2384),
.C(n_2371),
.Y(n_3523)
);

AOI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_3270),
.A2(n_2760),
.B(n_2752),
.Y(n_3524)
);

A2O1A1Ixp33_ASAP7_75t_SL g3525 ( 
.A1(n_3242),
.A2(n_2943),
.B(n_2942),
.C(n_2897),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_SL g3526 ( 
.A(n_3209),
.B(n_2751),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3365),
.B(n_2878),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3345),
.A2(n_3093),
.B(n_2384),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3345),
.A2(n_2371),
.B(n_2619),
.Y(n_3529)
);

OAI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3236),
.A2(n_2504),
.B1(n_2523),
.B2(n_2473),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3236),
.A2(n_2473),
.B1(n_2910),
.B2(n_2538),
.Y(n_3531)
);

OAI21x1_ASAP7_75t_L g3532 ( 
.A1(n_3208),
.A2(n_2867),
.B(n_2741),
.Y(n_3532)
);

AOI21x1_ASAP7_75t_L g3533 ( 
.A1(n_3191),
.A2(n_3229),
.B(n_3208),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_SL g3534 ( 
.A(n_3238),
.B(n_2874),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_SL g3535 ( 
.A(n_3209),
.B(n_2751),
.Y(n_3535)
);

OAI21xp33_ASAP7_75t_SL g3536 ( 
.A1(n_3377),
.A2(n_2550),
.B(n_2526),
.Y(n_3536)
);

INVx3_ASAP7_75t_L g3537 ( 
.A(n_3209),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_3261),
.A2(n_2867),
.B(n_2597),
.Y(n_3538)
);

A2O1A1Ixp33_ASAP7_75t_L g3539 ( 
.A1(n_3361),
.A2(n_2550),
.B(n_2768),
.C(n_2729),
.Y(n_3539)
);

OAI22xp33_ASAP7_75t_L g3540 ( 
.A1(n_3278),
.A2(n_2807),
.B1(n_2420),
.B2(n_2473),
.Y(n_3540)
);

AOI21x1_ASAP7_75t_L g3541 ( 
.A1(n_3229),
.A2(n_2881),
.B(n_2879),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3386),
.B(n_2896),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3215),
.B(n_2923),
.Y(n_3543)
);

AOI221xp5_ASAP7_75t_L g3544 ( 
.A1(n_3205),
.A2(n_2526),
.B1(n_2574),
.B2(n_2571),
.C(n_2729),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3263),
.B(n_2908),
.Y(n_3545)
);

NOR3xp33_ASAP7_75t_L g3546 ( 
.A(n_3275),
.B(n_2897),
.C(n_2855),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3307),
.B(n_136),
.Y(n_3547)
);

A2O1A1Ixp33_ASAP7_75t_L g3548 ( 
.A1(n_3361),
.A2(n_2768),
.B(n_2801),
.C(n_2791),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_SL g3549 ( 
.A(n_3238),
.B(n_2899),
.Y(n_3549)
);

NAND2xp33_ASAP7_75t_L g3550 ( 
.A(n_3330),
.B(n_3385),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3210),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3217),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3263),
.B(n_2922),
.Y(n_3553)
);

O2A1O1Ixp5_ASAP7_75t_L g3554 ( 
.A1(n_3323),
.A2(n_2911),
.B(n_2539),
.C(n_2427),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3261),
.A2(n_2910),
.B(n_2539),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3268),
.A2(n_2857),
.B(n_2572),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3215),
.B(n_2751),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3268),
.B(n_2924),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3278),
.A2(n_2926),
.B1(n_2934),
.B2(n_2933),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3232),
.Y(n_3560)
);

OAI21x1_ASAP7_75t_L g3561 ( 
.A1(n_3249),
.A2(n_2741),
.B(n_2857),
.Y(n_3561)
);

NAND2x1p5_ASAP7_75t_L g3562 ( 
.A(n_3239),
.B(n_3252),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3362),
.B(n_2938),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_3367),
.B(n_3379),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_SL g3565 ( 
.A(n_3215),
.B(n_2853),
.Y(n_3565)
);

NOR2xp67_ASAP7_75t_L g3566 ( 
.A(n_3239),
.B(n_2911),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3372),
.B(n_2940),
.Y(n_3567)
);

A2O1A1Ixp33_ASAP7_75t_SL g3568 ( 
.A1(n_3249),
.A2(n_2427),
.B(n_2341),
.C(n_2547),
.Y(n_3568)
);

OAI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3198),
.A2(n_2568),
.B(n_2761),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_3387),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3245),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3373),
.B(n_2941),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3252),
.A2(n_2899),
.B1(n_2791),
.B2(n_2801),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3382),
.A2(n_2890),
.B(n_2795),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_3312),
.B(n_2786),
.Y(n_3575)
);

OAI21x1_ASAP7_75t_L g3576 ( 
.A1(n_3198),
.A2(n_2761),
.B(n_2580),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3376),
.B(n_2953),
.Y(n_3577)
);

OR2x2_ASAP7_75t_L g3578 ( 
.A(n_3277),
.B(n_2786),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3246),
.B(n_2786),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_SL g3580 ( 
.A(n_3312),
.B(n_3330),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3326),
.A2(n_2808),
.B(n_2795),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3326),
.A2(n_2808),
.B(n_2795),
.Y(n_3582)
);

CKINVDCx5p33_ASAP7_75t_R g3583 ( 
.A(n_3279),
.Y(n_3583)
);

O2A1O1Ixp5_ASAP7_75t_SL g3584 ( 
.A1(n_3254),
.A2(n_2565),
.B(n_2558),
.C(n_2589),
.Y(n_3584)
);

AO22x1_ASAP7_75t_L g3585 ( 
.A1(n_3194),
.A2(n_2722),
.B1(n_2651),
.B2(n_2630),
.Y(n_3585)
);

OR2x6_ASAP7_75t_L g3586 ( 
.A(n_3183),
.B(n_3194),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3366),
.B(n_2808),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3325),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3369),
.B(n_2810),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3231),
.A2(n_2826),
.B(n_2810),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3257),
.Y(n_3591)
);

A2O1A1Ixp33_ASAP7_75t_L g3592 ( 
.A1(n_3381),
.A2(n_2722),
.B(n_2565),
.C(n_2558),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3258),
.B(n_2810),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3231),
.A2(n_2845),
.B(n_2826),
.Y(n_3594)
);

BUFx6f_ASAP7_75t_L g3595 ( 
.A(n_3292),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3312),
.Y(n_3596)
);

OAI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3383),
.A2(n_2651),
.B(n_2630),
.Y(n_3597)
);

O2A1O1Ixp33_ASAP7_75t_L g3598 ( 
.A1(n_3260),
.A2(n_3264),
.B(n_3293),
.C(n_3285),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3256),
.A2(n_2845),
.B(n_2826),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3256),
.A2(n_2853),
.B(n_2845),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3295),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3394),
.A2(n_3302),
.B(n_3383),
.Y(n_3602)
);

OAI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3390),
.A2(n_3407),
.B(n_3401),
.Y(n_3603)
);

OAI21x1_ASAP7_75t_L g3604 ( 
.A1(n_3584),
.A2(n_3344),
.B(n_3343),
.Y(n_3604)
);

INVx3_ASAP7_75t_L g3605 ( 
.A(n_3469),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3413),
.B(n_3299),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3461),
.B(n_3447),
.Y(n_3607)
);

OAI21x1_ASAP7_75t_L g3608 ( 
.A1(n_3399),
.A2(n_3350),
.B(n_3348),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3424),
.B(n_3309),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3473),
.B(n_3320),
.Y(n_3610)
);

OAI21x1_ASAP7_75t_L g3611 ( 
.A1(n_3408),
.A2(n_3304),
.B(n_3303),
.Y(n_3611)
);

AO21x1_ASAP7_75t_L g3612 ( 
.A1(n_3414),
.A2(n_3320),
.B(n_3289),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_L g3613 ( 
.A(n_3395),
.B(n_3275),
.Y(n_3613)
);

CKINVDCx5p33_ASAP7_75t_R g3614 ( 
.A(n_3451),
.Y(n_3614)
);

INVx3_ASAP7_75t_L g3615 ( 
.A(n_3570),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3423),
.A2(n_3319),
.B(n_3306),
.Y(n_3616)
);

BUFx2_ASAP7_75t_L g3617 ( 
.A(n_3570),
.Y(n_3617)
);

OAI21x1_ASAP7_75t_L g3618 ( 
.A1(n_3541),
.A2(n_3462),
.B(n_3529),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_3402),
.A2(n_3597),
.B(n_3585),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3443),
.B(n_3289),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3452),
.B(n_3181),
.Y(n_3621)
);

INVx3_ASAP7_75t_L g3622 ( 
.A(n_3459),
.Y(n_3622)
);

CKINVDCx8_ASAP7_75t_R g3623 ( 
.A(n_3468),
.Y(n_3623)
);

OAI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3489),
.A2(n_3384),
.B(n_3353),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3497),
.B(n_3338),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_SL g3626 ( 
.A1(n_3432),
.A2(n_3276),
.B(n_3333),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_SL g3627 ( 
.A(n_3457),
.B(n_3292),
.Y(n_3627)
);

OA22x2_ASAP7_75t_L g3628 ( 
.A1(n_3464),
.A2(n_3183),
.B1(n_3324),
.B2(n_3338),
.Y(n_3628)
);

AOI221x1_ASAP7_75t_L g3629 ( 
.A1(n_3547),
.A2(n_3334),
.B1(n_3331),
.B2(n_3328),
.C(n_3222),
.Y(n_3629)
);

AO31x2_ASAP7_75t_L g3630 ( 
.A1(n_3521),
.A2(n_3337),
.A3(n_3336),
.B(n_3219),
.Y(n_3630)
);

NOR2xp67_ASAP7_75t_L g3631 ( 
.A(n_3455),
.B(n_3302),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3412),
.A2(n_3302),
.B(n_3252),
.Y(n_3632)
);

OAI21x1_ASAP7_75t_SL g3633 ( 
.A1(n_3421),
.A2(n_3428),
.B(n_3598),
.Y(n_3633)
);

AO21x1_ASAP7_75t_L g3634 ( 
.A1(n_3484),
.A2(n_3276),
.B(n_3346),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3420),
.A2(n_3346),
.B(n_3353),
.Y(n_3635)
);

AOI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3533),
.A2(n_3475),
.B(n_3454),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3490),
.A2(n_3384),
.B(n_3371),
.Y(n_3637)
);

OAI22xp5_ASAP7_75t_L g3638 ( 
.A1(n_3429),
.A2(n_3330),
.B1(n_3375),
.B2(n_3371),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3438),
.B(n_3200),
.Y(n_3639)
);

NAND2x1p5_ASAP7_75t_L g3640 ( 
.A(n_3404),
.B(n_3292),
.Y(n_3640)
);

INVx3_ASAP7_75t_L g3641 ( 
.A(n_3459),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_SL g3642 ( 
.A(n_3439),
.B(n_3371),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3478),
.A2(n_3385),
.B(n_3375),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3397),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3398),
.Y(n_3645)
);

OAI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3524),
.A2(n_2580),
.B(n_3247),
.Y(n_3646)
);

INVx3_ASAP7_75t_L g3647 ( 
.A(n_3459),
.Y(n_3647)
);

AO21x1_ASAP7_75t_L g3648 ( 
.A1(n_3494),
.A2(n_3324),
.B(n_3250),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3403),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3538),
.A2(n_3576),
.B(n_3532),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3393),
.B(n_3375),
.Y(n_3651)
);

BUFx3_ASAP7_75t_L g3652 ( 
.A(n_3474),
.Y(n_3652)
);

AOI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3512),
.A2(n_3385),
.B(n_2877),
.Y(n_3653)
);

BUFx6f_ASAP7_75t_L g3654 ( 
.A(n_3422),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_L g3655 ( 
.A1(n_3515),
.A2(n_2656),
.B(n_2652),
.Y(n_3655)
);

INVx6_ASAP7_75t_SL g3656 ( 
.A(n_3586),
.Y(n_3656)
);

OAI21x1_ASAP7_75t_L g3657 ( 
.A1(n_3528),
.A2(n_2656),
.B(n_2652),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3505),
.B(n_91),
.Y(n_3658)
);

AND2x4_ASAP7_75t_L g3659 ( 
.A(n_3458),
.B(n_2853),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3411),
.A2(n_2651),
.B(n_2630),
.Y(n_3660)
);

OAI22xp5_ASAP7_75t_L g3661 ( 
.A1(n_3431),
.A2(n_2880),
.B1(n_2923),
.B2(n_2877),
.Y(n_3661)
);

BUFx2_ASAP7_75t_L g3662 ( 
.A(n_3510),
.Y(n_3662)
);

OAI21x1_ASAP7_75t_L g3663 ( 
.A1(n_3561),
.A2(n_2454),
.B(n_2444),
.Y(n_3663)
);

BUFx6f_ASAP7_75t_L g3664 ( 
.A(n_3422),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3505),
.B(n_92),
.Y(n_3665)
);

OAI21x1_ASAP7_75t_L g3666 ( 
.A1(n_3493),
.A2(n_2457),
.B(n_2441),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3499),
.A2(n_2880),
.B(n_2877),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3513),
.A2(n_2341),
.B(n_2549),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3495),
.B(n_92),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3568),
.A2(n_2923),
.B(n_2880),
.Y(n_3670)
);

INVx3_ASAP7_75t_SL g3671 ( 
.A(n_3501),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3436),
.A2(n_2541),
.B(n_2532),
.Y(n_3672)
);

AND2x2_ASAP7_75t_SL g3673 ( 
.A(n_3396),
.B(n_2532),
.Y(n_3673)
);

OAI21x1_ASAP7_75t_L g3674 ( 
.A1(n_3555),
.A2(n_2651),
.B(n_2630),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3525),
.A2(n_2541),
.B(n_2532),
.Y(n_3675)
);

AOI31xp67_ASAP7_75t_L g3676 ( 
.A1(n_3416),
.A2(n_2651),
.A3(n_2630),
.B(n_94),
.Y(n_3676)
);

OAI21x1_ASAP7_75t_L g3677 ( 
.A1(n_3556),
.A2(n_2541),
.B(n_2532),
.Y(n_3677)
);

OAI22x1_ASAP7_75t_L g3678 ( 
.A1(n_3477),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3678)
);

OA22x2_ASAP7_75t_L g3679 ( 
.A1(n_3464),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3679)
);

OAI21xp5_ASAP7_75t_L g3680 ( 
.A1(n_3411),
.A2(n_3554),
.B(n_3450),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3523),
.A2(n_2552),
.B(n_2541),
.Y(n_3681)
);

INVxp67_ASAP7_75t_L g3682 ( 
.A(n_3488),
.Y(n_3682)
);

OAI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3502),
.A2(n_93),
.B(n_95),
.Y(n_3683)
);

INVx5_ASAP7_75t_L g3684 ( 
.A(n_3440),
.Y(n_3684)
);

NAND3xp33_ASAP7_75t_L g3685 ( 
.A(n_3544),
.B(n_2552),
.C(n_96),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3467),
.A2(n_2552),
.B(n_96),
.Y(n_3686)
);

A2O1A1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3476),
.A2(n_2552),
.B(n_98),
.C(n_96),
.Y(n_3687)
);

HB1xp67_ASAP7_75t_L g3688 ( 
.A(n_3419),
.Y(n_3688)
);

OAI21x1_ASAP7_75t_L g3689 ( 
.A1(n_3472),
.A2(n_97),
.B(n_98),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3410),
.Y(n_3690)
);

AOI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_3449),
.A2(n_97),
.B(n_98),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3433),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3500),
.B(n_3519),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3445),
.A2(n_97),
.B(n_99),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3400),
.Y(n_3695)
);

OAI21x1_ASAP7_75t_L g3696 ( 
.A1(n_3430),
.A2(n_99),
.B(n_100),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3391),
.B(n_99),
.Y(n_3697)
);

O2A1O1Ixp5_ASAP7_75t_L g3698 ( 
.A1(n_3442),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_3698)
);

OAI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3504),
.A2(n_100),
.B(n_101),
.Y(n_3699)
);

OAI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3504),
.A2(n_101),
.B(n_102),
.Y(n_3700)
);

OAI21x1_ASAP7_75t_L g3701 ( 
.A1(n_3569),
.A2(n_103),
.B(n_104),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3590),
.A2(n_3599),
.B(n_3594),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3471),
.B(n_103),
.Y(n_3703)
);

OAI21x1_ASAP7_75t_L g3704 ( 
.A1(n_3600),
.A2(n_104),
.B(n_105),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3427),
.B(n_104),
.Y(n_3705)
);

OAI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3536),
.A2(n_105),
.B(n_106),
.Y(n_3706)
);

OAI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3574),
.A2(n_105),
.B(n_106),
.Y(n_3707)
);

A2O1A1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3476),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_3708)
);

NOR2xp67_ASAP7_75t_L g3709 ( 
.A(n_3440),
.B(n_137),
.Y(n_3709)
);

OAI21x1_ASAP7_75t_L g3710 ( 
.A1(n_3483),
.A2(n_107),
.B(n_108),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3509),
.B(n_107),
.Y(n_3711)
);

CKINVDCx5p33_ASAP7_75t_R g3712 ( 
.A(n_3425),
.Y(n_3712)
);

OAI21x1_ASAP7_75t_L g3713 ( 
.A1(n_3506),
.A2(n_3562),
.B(n_3517),
.Y(n_3713)
);

BUFx6f_ASAP7_75t_L g3714 ( 
.A(n_3422),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3492),
.B(n_108),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3507),
.B(n_109),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3511),
.B(n_109),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3518),
.B(n_110),
.Y(n_3718)
);

OAI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3389),
.A2(n_111),
.B(n_112),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3551),
.B(n_111),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3550),
.A2(n_3463),
.B(n_3526),
.Y(n_3721)
);

OAI21xp33_ASAP7_75t_L g3722 ( 
.A1(n_3437),
.A2(n_112),
.B(n_113),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3535),
.A2(n_112),
.B(n_113),
.Y(n_3723)
);

BUFx12f_ASAP7_75t_L g3724 ( 
.A(n_3487),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3543),
.A2(n_113),
.B(n_114),
.Y(n_3725)
);

AO31x2_ASAP7_75t_L g3726 ( 
.A1(n_3441),
.A2(n_116),
.A3(n_114),
.B(n_115),
.Y(n_3726)
);

OR2x2_ASAP7_75t_L g3727 ( 
.A(n_3552),
.B(n_114),
.Y(n_3727)
);

NAND3xp33_ASAP7_75t_L g3728 ( 
.A(n_3593),
.B(n_3508),
.C(n_3579),
.Y(n_3728)
);

A2O1A1Ixp33_ASAP7_75t_L g3729 ( 
.A1(n_3536),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3560),
.B(n_116),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3571),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3426),
.A2(n_120),
.B1(n_121),
.B2(n_118),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3591),
.B(n_117),
.Y(n_3733)
);

O2A1O1Ixp5_ASAP7_75t_L g3734 ( 
.A1(n_3580),
.A2(n_121),
.B(n_118),
.C(n_120),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3601),
.Y(n_3735)
);

NAND2x1p5_ASAP7_75t_L g3736 ( 
.A(n_3404),
.B(n_138),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3596),
.B(n_120),
.Y(n_3737)
);

INVx2_ASAP7_75t_SL g3738 ( 
.A(n_3583),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_3557),
.A2(n_121),
.B(n_122),
.Y(n_3739)
);

BUFx2_ASAP7_75t_L g3740 ( 
.A(n_3496),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3485),
.A2(n_122),
.B(n_123),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3565),
.A2(n_122),
.B(n_124),
.Y(n_3742)
);

AO31x2_ASAP7_75t_L g3743 ( 
.A1(n_3448),
.A2(n_3539),
.A3(n_3567),
.B(n_3563),
.Y(n_3743)
);

AO21x1_ASAP7_75t_L g3744 ( 
.A1(n_3527),
.A2(n_124),
.B(n_125),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3406),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3549),
.A2(n_3548),
.B(n_3575),
.Y(n_3746)
);

OAI21x1_ASAP7_75t_L g3747 ( 
.A1(n_3434),
.A2(n_124),
.B(n_125),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3417),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_3466),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3480),
.B(n_126),
.Y(n_3750)
);

AOI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_3516),
.A2(n_126),
.B(n_127),
.Y(n_3751)
);

BUFx6f_ASAP7_75t_L g3752 ( 
.A(n_3444),
.Y(n_3752)
);

AOI221x1_ASAP7_75t_L g3753 ( 
.A1(n_3446),
.A2(n_3546),
.B1(n_3520),
.B2(n_3498),
.C(n_3564),
.Y(n_3753)
);

BUFx5_ASAP7_75t_L g3754 ( 
.A(n_3453),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3465),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3481),
.B(n_127),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3486),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3514),
.Y(n_3758)
);

NAND3xp33_ASAP7_75t_L g3759 ( 
.A(n_3587),
.B(n_128),
.C(n_139),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3588),
.Y(n_3760)
);

AOI221x1_ASAP7_75t_L g3761 ( 
.A1(n_3415),
.A2(n_128),
.B1(n_142),
.B2(n_140),
.C(n_143),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_3534),
.A2(n_140),
.B(n_142),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3470),
.A2(n_144),
.B(n_145),
.Y(n_3763)
);

OA21x2_ASAP7_75t_L g3764 ( 
.A1(n_3482),
.A2(n_144),
.B(n_146),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3531),
.A2(n_146),
.B(n_147),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3540),
.A2(n_3405),
.B(n_3491),
.Y(n_3766)
);

NAND3xp33_ASAP7_75t_L g3767 ( 
.A(n_3589),
.B(n_149),
.C(n_148),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3522),
.A2(n_687),
.B1(n_688),
.B2(n_686),
.Y(n_3768)
);

OAI22xp5_ASAP7_75t_L g3769 ( 
.A1(n_3522),
.A2(n_687),
.B1(n_688),
.B2(n_686),
.Y(n_3769)
);

BUFx2_ASAP7_75t_L g3770 ( 
.A(n_3415),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3537),
.B(n_147),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3405),
.A2(n_148),
.B(n_149),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3581),
.A2(n_3582),
.B(n_3573),
.Y(n_3773)
);

AOI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3530),
.A2(n_150),
.B(n_151),
.Y(n_3774)
);

OAI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3409),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_3775)
);

AOI21x1_ASAP7_75t_SL g3776 ( 
.A1(n_3468),
.A2(n_154),
.B(n_155),
.Y(n_3776)
);

OAI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_3460),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3777)
);

INVx1_ASAP7_75t_SL g3778 ( 
.A(n_3578),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3537),
.A2(n_3577),
.B(n_3572),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3559),
.A2(n_3553),
.B(n_3545),
.Y(n_3780)
);

NAND2xp33_ASAP7_75t_L g3781 ( 
.A(n_3444),
.B(n_3479),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3566),
.A2(n_158),
.B(n_159),
.Y(n_3782)
);

CKINVDCx20_ASAP7_75t_R g3783 ( 
.A(n_3396),
.Y(n_3783)
);

NOR2x1_ASAP7_75t_SL g3784 ( 
.A(n_3586),
.B(n_158),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3558),
.B(n_159),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3542),
.Y(n_3786)
);

OA21x2_ASAP7_75t_L g3787 ( 
.A1(n_3592),
.A2(n_3418),
.B(n_3503),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3595),
.B(n_160),
.Y(n_3788)
);

OAI21x1_ASAP7_75t_L g3789 ( 
.A1(n_3453),
.A2(n_161),
.B(n_162),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3595),
.B(n_161),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3595),
.B(n_163),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3503),
.B(n_163),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3586),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3503),
.A2(n_164),
.B(n_165),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3435),
.A2(n_164),
.B(n_166),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3479),
.B(n_166),
.Y(n_3796)
);

AND2x4_ASAP7_75t_L g3797 ( 
.A(n_3392),
.B(n_168),
.Y(n_3797)
);

OR2x6_ASAP7_75t_L g3798 ( 
.A(n_3392),
.B(n_168),
.Y(n_3798)
);

NOR2xp67_ASAP7_75t_L g3799 ( 
.A(n_3479),
.B(n_169),
.Y(n_3799)
);

OAI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3456),
.A2(n_169),
.B(n_170),
.Y(n_3800)
);

BUFx5_ASAP7_75t_L g3801 ( 
.A(n_3444),
.Y(n_3801)
);

O2A1O1Ixp5_ASAP7_75t_L g3802 ( 
.A1(n_3390),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3584),
.A2(n_172),
.B(n_173),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3443),
.B(n_173),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3398),
.Y(n_3805)
);

NOR2xp67_ASAP7_75t_SL g3806 ( 
.A(n_3487),
.B(n_174),
.Y(n_3806)
);

AO31x2_ASAP7_75t_L g3807 ( 
.A1(n_3521),
.A2(n_178),
.A3(n_176),
.B(n_177),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3584),
.A2(n_176),
.B(n_179),
.Y(n_3808)
);

OAI21x1_ASAP7_75t_L g3809 ( 
.A1(n_3584),
.A2(n_179),
.B(n_180),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3395),
.B(n_181),
.Y(n_3810)
);

AOI211x1_ASAP7_75t_L g3811 ( 
.A1(n_3432),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3429),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_3812)
);

O2A1O1Ixp5_ASAP7_75t_L g3813 ( 
.A1(n_3390),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3395),
.B(n_185),
.Y(n_3814)
);

AOI211x1_ASAP7_75t_L g3815 ( 
.A1(n_3432),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_3815)
);

OAI21x1_ASAP7_75t_L g3816 ( 
.A1(n_3584),
.A2(n_188),
.B(n_189),
.Y(n_3816)
);

OAI21x1_ASAP7_75t_L g3817 ( 
.A1(n_3584),
.A2(n_189),
.B(n_190),
.Y(n_3817)
);

OAI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3390),
.A2(n_191),
.B(n_192),
.Y(n_3818)
);

OAI21x1_ASAP7_75t_L g3819 ( 
.A1(n_3584),
.A2(n_191),
.B(n_192),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3584),
.A2(n_193),
.B(n_194),
.Y(n_3820)
);

AOI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3394),
.A2(n_193),
.B(n_194),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_L g3822 ( 
.A1(n_3584),
.A2(n_195),
.B(n_196),
.Y(n_3822)
);

OAI21x1_ASAP7_75t_L g3823 ( 
.A1(n_3584),
.A2(n_197),
.B(n_198),
.Y(n_3823)
);

INVx3_ASAP7_75t_L g3824 ( 
.A(n_3469),
.Y(n_3824)
);

AOI21xp33_ASAP7_75t_L g3825 ( 
.A1(n_3414),
.A2(n_199),
.B(n_200),
.Y(n_3825)
);

AND2x2_ASAP7_75t_SL g3826 ( 
.A(n_3439),
.B(n_201),
.Y(n_3826)
);

OAI21x1_ASAP7_75t_L g3827 ( 
.A1(n_3584),
.A2(n_202),
.B(n_203),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3429),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3443),
.B(n_204),
.Y(n_3829)
);

AO31x2_ASAP7_75t_L g3830 ( 
.A1(n_3521),
.A2(n_209),
.A3(n_205),
.B(n_206),
.Y(n_3830)
);

A2O1A1Ixp33_ASAP7_75t_L g3831 ( 
.A1(n_3722),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_3831)
);

BUFx8_ASAP7_75t_L g3832 ( 
.A(n_3724),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3603),
.A2(n_211),
.B(n_212),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3603),
.A2(n_213),
.B(n_214),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3644),
.Y(n_3835)
);

AOI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3660),
.A2(n_213),
.B(n_214),
.Y(n_3836)
);

AO32x2_ASAP7_75t_L g3837 ( 
.A1(n_3661),
.A2(n_3828),
.A3(n_3812),
.B1(n_3638),
.B2(n_3768),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3821),
.A2(n_215),
.B(n_216),
.Y(n_3838)
);

OAI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3632),
.A2(n_215),
.B(n_216),
.Y(n_3839)
);

OR2x6_ASAP7_75t_L g3840 ( 
.A(n_3766),
.B(n_217),
.Y(n_3840)
);

AOI21xp33_ASAP7_75t_L g3841 ( 
.A1(n_3633),
.A2(n_217),
.B(n_218),
.Y(n_3841)
);

AO31x2_ASAP7_75t_L g3842 ( 
.A1(n_3648),
.A2(n_3629),
.A3(n_3634),
.B(n_3729),
.Y(n_3842)
);

AO31x2_ASAP7_75t_L g3843 ( 
.A1(n_3708),
.A2(n_220),
.A3(n_218),
.B(n_219),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3649),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_SL g3845 ( 
.A(n_3612),
.B(n_219),
.Y(n_3845)
);

CKINVDCx5p33_ASAP7_75t_R g3846 ( 
.A(n_3712),
.Y(n_3846)
);

AOI21xp5_ASAP7_75t_L g3847 ( 
.A1(n_3699),
.A2(n_220),
.B(n_221),
.Y(n_3847)
);

AOI221xp5_ASAP7_75t_L g3848 ( 
.A1(n_3722),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.C(n_224),
.Y(n_3848)
);

INVx3_ASAP7_75t_L g3849 ( 
.A(n_3622),
.Y(n_3849)
);

INVx5_ASAP7_75t_L g3850 ( 
.A(n_3798),
.Y(n_3850)
);

INVx2_ASAP7_75t_SL g3851 ( 
.A(n_3652),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3699),
.A2(n_222),
.B(n_223),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_3614),
.Y(n_3853)
);

INVx3_ASAP7_75t_SL g3854 ( 
.A(n_3671),
.Y(n_3854)
);

NAND3xp33_ASAP7_75t_L g3855 ( 
.A(n_3753),
.B(n_224),
.C(n_225),
.Y(n_3855)
);

AOI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3700),
.A2(n_225),
.B(n_226),
.Y(n_3856)
);

AOI21xp33_ASAP7_75t_L g3857 ( 
.A1(n_3679),
.A2(n_227),
.B(n_228),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3645),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3695),
.Y(n_3859)
);

OAI21x1_ASAP7_75t_L g3860 ( 
.A1(n_3636),
.A2(n_228),
.B(n_229),
.Y(n_3860)
);

OR2x6_ASAP7_75t_L g3861 ( 
.A(n_3619),
.B(n_3635),
.Y(n_3861)
);

A2O1A1Ixp33_ASAP7_75t_L g3862 ( 
.A1(n_3818),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3758),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3805),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3688),
.B(n_230),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3745),
.Y(n_3866)
);

BUFx2_ASAP7_75t_L g3867 ( 
.A(n_3617),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3700),
.A2(n_3683),
.B(n_3680),
.Y(n_3868)
);

OAI21x1_ASAP7_75t_L g3869 ( 
.A1(n_3650),
.A2(n_232),
.B(n_233),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3683),
.A2(n_234),
.B(n_235),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3685),
.A2(n_234),
.B(n_235),
.Y(n_3871)
);

INVx1_ASAP7_75t_SL g3872 ( 
.A(n_3740),
.Y(n_3872)
);

OAI22xp5_ASAP7_75t_L g3873 ( 
.A1(n_3811),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3873)
);

OAI22xp5_ASAP7_75t_L g3874 ( 
.A1(n_3811),
.A2(n_240),
.B1(n_236),
.B2(n_239),
.Y(n_3874)
);

OAI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3802),
.A2(n_239),
.B(n_241),
.Y(n_3875)
);

AOI21xp5_ASAP7_75t_L g3876 ( 
.A1(n_3685),
.A2(n_241),
.B(n_242),
.Y(n_3876)
);

OAI21x1_ASAP7_75t_L g3877 ( 
.A1(n_3618),
.A2(n_243),
.B(n_244),
.Y(n_3877)
);

A2O1A1Ixp33_ASAP7_75t_L g3878 ( 
.A1(n_3687),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_3878)
);

A2O1A1Ixp33_ASAP7_75t_L g3879 ( 
.A1(n_3719),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_3879)
);

OAI22xp33_ASAP7_75t_L g3880 ( 
.A1(n_3628),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3605),
.B(n_249),
.Y(n_3881)
);

AOI21x1_ASAP7_75t_L g3882 ( 
.A1(n_3764),
.A2(n_251),
.B(n_252),
.Y(n_3882)
);

OR2x2_ASAP7_75t_L g3883 ( 
.A(n_3778),
.B(n_251),
.Y(n_3883)
);

AO21x2_ASAP7_75t_L g3884 ( 
.A1(n_3706),
.A2(n_252),
.B(n_253),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3690),
.Y(n_3885)
);

BUFx2_ASAP7_75t_L g3886 ( 
.A(n_3615),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3692),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3731),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3735),
.Y(n_3889)
);

NOR2xp33_ASAP7_75t_SL g3890 ( 
.A(n_3783),
.B(n_253),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3786),
.Y(n_3891)
);

AOI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3602),
.A2(n_254),
.B(n_255),
.Y(n_3892)
);

AOI31xp67_ASAP7_75t_L g3893 ( 
.A1(n_3785),
.A2(n_3705),
.A3(n_3697),
.B(n_3627),
.Y(n_3893)
);

AO32x2_ASAP7_75t_L g3894 ( 
.A1(n_3769),
.A2(n_257),
.A3(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_3894)
);

HB1xp67_ASAP7_75t_L g3895 ( 
.A(n_3662),
.Y(n_3895)
);

NAND3x1_ASAP7_75t_L g3896 ( 
.A(n_3605),
.B(n_256),
.C(n_257),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3706),
.A2(n_258),
.B(n_259),
.Y(n_3897)
);

OAI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3813),
.A2(n_3814),
.B(n_3810),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_3773),
.A2(n_259),
.B(n_260),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3693),
.B(n_262),
.Y(n_3900)
);

AND2x4_ASAP7_75t_L g3901 ( 
.A(n_3793),
.B(n_262),
.Y(n_3901)
);

AOI221xp5_ASAP7_75t_L g3902 ( 
.A1(n_3678),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_3902)
);

AOI221xp5_ASAP7_75t_L g3903 ( 
.A1(n_3815),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3642),
.A2(n_267),
.B(n_268),
.Y(n_3904)
);

AO31x2_ASAP7_75t_L g3905 ( 
.A1(n_3744),
.A2(n_271),
.A3(n_269),
.B(n_270),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3824),
.B(n_269),
.Y(n_3906)
);

OAI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3767),
.A2(n_271),
.B(n_272),
.Y(n_3907)
);

O2A1O1Ixp33_ASAP7_75t_L g3908 ( 
.A1(n_3825),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3746),
.A2(n_273),
.B(n_274),
.Y(n_3909)
);

AO31x2_ASAP7_75t_L g3910 ( 
.A1(n_3761),
.A2(n_277),
.A3(n_275),
.B(n_276),
.Y(n_3910)
);

INVxp67_ASAP7_75t_SL g3911 ( 
.A(n_3631),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_3637),
.A2(n_275),
.B(n_278),
.Y(n_3912)
);

BUFx6f_ASAP7_75t_L g3913 ( 
.A(n_3654),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3815),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_3914)
);

AO31x2_ASAP7_75t_L g3915 ( 
.A1(n_3748),
.A2(n_282),
.A3(n_279),
.B(n_280),
.Y(n_3915)
);

A2O1A1Ixp33_ASAP7_75t_L g3916 ( 
.A1(n_3772),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_3916)
);

O2A1O1Ixp33_ASAP7_75t_L g3917 ( 
.A1(n_3777),
.A2(n_286),
.B(n_283),
.C(n_285),
.Y(n_3917)
);

NAND3xp33_ASAP7_75t_L g3918 ( 
.A(n_3728),
.B(n_285),
.C(n_286),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3779),
.Y(n_3919)
);

CKINVDCx20_ASAP7_75t_R g3920 ( 
.A(n_3623),
.Y(n_3920)
);

NOR2xp67_ASAP7_75t_L g3921 ( 
.A(n_3631),
.B(n_287),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3667),
.A2(n_287),
.B(n_288),
.Y(n_3922)
);

OAI21x1_ASAP7_75t_L g3923 ( 
.A1(n_3604),
.A2(n_288),
.B(n_289),
.Y(n_3923)
);

OAI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3646),
.A2(n_289),
.B(n_290),
.Y(n_3924)
);

OAI21x1_ASAP7_75t_L g3925 ( 
.A1(n_3702),
.A2(n_290),
.B(n_291),
.Y(n_3925)
);

OAI21x1_ASAP7_75t_L g3926 ( 
.A1(n_3713),
.A2(n_292),
.B(n_293),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3639),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3607),
.B(n_292),
.Y(n_3928)
);

AO31x2_ASAP7_75t_L g3929 ( 
.A1(n_3755),
.A2(n_296),
.A3(n_294),
.B(n_295),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3609),
.B(n_294),
.Y(n_3930)
);

OR2x2_ASAP7_75t_L g3931 ( 
.A(n_3778),
.B(n_295),
.Y(n_3931)
);

OAI21x1_ASAP7_75t_L g3932 ( 
.A1(n_3611),
.A2(n_3608),
.B(n_3616),
.Y(n_3932)
);

HB1xp67_ASAP7_75t_L g3933 ( 
.A(n_3610),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3728),
.B(n_296),
.Y(n_3934)
);

NOR2xp33_ASAP7_75t_L g3935 ( 
.A(n_3682),
.B(n_298),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3643),
.A2(n_3653),
.B(n_3694),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3606),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3681),
.A2(n_299),
.B(n_300),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3672),
.A2(n_299),
.B(n_300),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3675),
.A2(n_301),
.B(n_302),
.Y(n_3940)
);

AO21x1_ASAP7_75t_L g3941 ( 
.A1(n_3703),
.A2(n_301),
.B(n_302),
.Y(n_3941)
);

NOR2xp33_ASAP7_75t_SL g3942 ( 
.A(n_3826),
.B(n_303),
.Y(n_3942)
);

CKINVDCx5p33_ASAP7_75t_R g3943 ( 
.A(n_3738),
.Y(n_3943)
);

BUFx10_ASAP7_75t_L g3944 ( 
.A(n_3798),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3621),
.Y(n_3945)
);

OR2x2_ASAP7_75t_L g3946 ( 
.A(n_3651),
.B(n_303),
.Y(n_3946)
);

AOI221x1_ASAP7_75t_L g3947 ( 
.A1(n_3711),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.C(n_307),
.Y(n_3947)
);

OAI21x1_ASAP7_75t_L g3948 ( 
.A1(n_3668),
.A2(n_304),
.B(n_305),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3615),
.B(n_308),
.Y(n_3949)
);

OAI21x1_ASAP7_75t_L g3950 ( 
.A1(n_3677),
.A2(n_308),
.B(n_309),
.Y(n_3950)
);

AO31x2_ASAP7_75t_L g3951 ( 
.A1(n_3757),
.A2(n_312),
.A3(n_310),
.B(n_311),
.Y(n_3951)
);

BUFx2_ASAP7_75t_L g3952 ( 
.A(n_3622),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3824),
.B(n_311),
.Y(n_3953)
);

AO31x2_ASAP7_75t_L g3954 ( 
.A1(n_3760),
.A2(n_3691),
.A3(n_3770),
.B(n_3784),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3733),
.B(n_3625),
.Y(n_3955)
);

OAI21x1_ASAP7_75t_L g3956 ( 
.A1(n_3780),
.A2(n_313),
.B(n_314),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3727),
.B(n_313),
.Y(n_3957)
);

CKINVDCx5p33_ASAP7_75t_R g3958 ( 
.A(n_3641),
.Y(n_3958)
);

INVx3_ASAP7_75t_L g3959 ( 
.A(n_3641),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3715),
.Y(n_3960)
);

AO21x2_ASAP7_75t_L g3961 ( 
.A1(n_3716),
.A2(n_315),
.B(n_316),
.Y(n_3961)
);

OA21x2_ASAP7_75t_L g3962 ( 
.A1(n_3626),
.A2(n_316),
.B(n_317),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3721),
.A2(n_317),
.B(n_318),
.Y(n_3963)
);

CKINVDCx20_ASAP7_75t_R g3964 ( 
.A(n_3620),
.Y(n_3964)
);

CKINVDCx5p33_ASAP7_75t_R g3965 ( 
.A(n_3647),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3630),
.Y(n_3966)
);

AOI21x1_ASAP7_75t_L g3967 ( 
.A1(n_3764),
.A2(n_319),
.B(n_320),
.Y(n_3967)
);

A2O1A1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3698),
.A2(n_322),
.B(n_319),
.C(n_321),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3717),
.Y(n_3969)
);

AO21x1_ASAP7_75t_L g3970 ( 
.A1(n_3718),
.A2(n_322),
.B(n_323),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3669),
.B(n_324),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3630),
.Y(n_3972)
);

A2O1A1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_3795),
.A2(n_328),
.B(n_325),
.C(n_326),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3670),
.A2(n_325),
.B(n_326),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3647),
.B(n_328),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3630),
.Y(n_3976)
);

AO31x2_ASAP7_75t_L g3977 ( 
.A1(n_3732),
.A2(n_332),
.A3(n_330),
.B(n_331),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3767),
.A2(n_330),
.B(n_331),
.Y(n_3978)
);

AOI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3775),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3613),
.B(n_333),
.Y(n_3980)
);

AOI221x1_ASAP7_75t_L g3981 ( 
.A1(n_3750),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.C(n_337),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3720),
.Y(n_3982)
);

NOR2xp33_ASAP7_75t_L g3983 ( 
.A(n_3797),
.B(n_335),
.Y(n_3983)
);

INVx1_ASAP7_75t_SL g3984 ( 
.A(n_3797),
.Y(n_3984)
);

AO31x2_ASAP7_75t_L g3985 ( 
.A1(n_3658),
.A2(n_339),
.A3(n_337),
.B(n_338),
.Y(n_3985)
);

OAI21x1_ASAP7_75t_L g3986 ( 
.A1(n_3674),
.A2(n_338),
.B(n_339),
.Y(n_3986)
);

A2O1A1Ixp33_ASAP7_75t_L g3987 ( 
.A1(n_3751),
.A2(n_343),
.B(n_340),
.C(n_341),
.Y(n_3987)
);

BUFx12f_ASAP7_75t_L g3988 ( 
.A(n_3798),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3730),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3756),
.B(n_340),
.Y(n_3990)
);

A2O1A1Ixp33_ASAP7_75t_L g3991 ( 
.A1(n_3707),
.A2(n_344),
.B(n_341),
.C(n_343),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3665),
.Y(n_3992)
);

INVx4_ASAP7_75t_L g3993 ( 
.A(n_3654),
.Y(n_3993)
);

A2O1A1Ixp33_ASAP7_75t_L g3994 ( 
.A1(n_3762),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_3994)
);

AOI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3800),
.A2(n_345),
.B(n_346),
.Y(n_3995)
);

AO21x2_ASAP7_75t_L g3996 ( 
.A1(n_3709),
.A2(n_347),
.B(n_348),
.Y(n_3996)
);

OAI21x1_ASAP7_75t_L g3997 ( 
.A1(n_3657),
.A2(n_348),
.B(n_349),
.Y(n_3997)
);

INVxp67_ASAP7_75t_L g3998 ( 
.A(n_3804),
.Y(n_3998)
);

OAI21x1_ASAP7_75t_L g3999 ( 
.A1(n_3666),
.A2(n_349),
.B(n_350),
.Y(n_3999)
);

INVx4_ASAP7_75t_L g4000 ( 
.A(n_3654),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3659),
.Y(n_4001)
);

AOI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_3800),
.A2(n_351),
.B(n_353),
.Y(n_4002)
);

AND2x4_ASAP7_75t_L g4003 ( 
.A(n_3659),
.B(n_354),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3759),
.A2(n_355),
.B(n_356),
.Y(n_4004)
);

AND2x6_ASAP7_75t_SL g4005 ( 
.A(n_3829),
.B(n_355),
.Y(n_4005)
);

NAND2xp33_ASAP7_75t_L g4006 ( 
.A(n_3801),
.B(n_356),
.Y(n_4006)
);

BUFx3_ASAP7_75t_L g4007 ( 
.A(n_3664),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3743),
.Y(n_4008)
);

BUFx3_ASAP7_75t_L g4009 ( 
.A(n_3664),
.Y(n_4009)
);

INVx1_ASAP7_75t_SL g4010 ( 
.A(n_3737),
.Y(n_4010)
);

A2O1A1Ixp33_ASAP7_75t_L g4011 ( 
.A1(n_3799),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_4011)
);

AO21x1_ASAP7_75t_SL g4012 ( 
.A1(n_3792),
.A2(n_357),
.B(n_359),
.Y(n_4012)
);

OAI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3868),
.A2(n_3759),
.B(n_3676),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3835),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_L g4015 ( 
.A(n_3928),
.B(n_3788),
.Y(n_4015)
);

O2A1O1Ixp33_ASAP7_75t_L g4016 ( 
.A1(n_3862),
.A2(n_3796),
.B(n_3734),
.C(n_3723),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3919),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3844),
.Y(n_4018)
);

NAND2x1p5_ASAP7_75t_L g4019 ( 
.A(n_3850),
.B(n_3787),
.Y(n_4019)
);

A2O1A1Ixp33_ASAP7_75t_L g4020 ( 
.A1(n_3855),
.A2(n_3709),
.B(n_3799),
.C(n_3624),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3885),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3857),
.A2(n_3749),
.B1(n_3725),
.B2(n_3742),
.Y(n_4022)
);

OAI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3932),
.A2(n_3787),
.B(n_3696),
.Y(n_4023)
);

CKINVDCx20_ASAP7_75t_R g4024 ( 
.A(n_3920),
.Y(n_4024)
);

AO21x2_ASAP7_75t_L g4025 ( 
.A1(n_4008),
.A2(n_3701),
.B(n_3790),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_3891),
.B(n_3807),
.Y(n_4026)
);

OAI21x1_ASAP7_75t_L g4027 ( 
.A1(n_3966),
.A2(n_3808),
.B(n_3803),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3887),
.B(n_3807),
.Y(n_4028)
);

NOR2x1_ASAP7_75t_R g4029 ( 
.A(n_3850),
.B(n_3684),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3866),
.Y(n_4030)
);

NAND2x1p5_ASAP7_75t_L g4031 ( 
.A(n_3850),
.B(n_3684),
.Y(n_4031)
);

OAI21x1_ASAP7_75t_L g4032 ( 
.A1(n_3972),
.A2(n_3816),
.B(n_3809),
.Y(n_4032)
);

OAI21x1_ASAP7_75t_L g4033 ( 
.A1(n_3976),
.A2(n_3819),
.B(n_3817),
.Y(n_4033)
);

BUFx12f_ASAP7_75t_SL g4034 ( 
.A(n_3840),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3888),
.B(n_3807),
.Y(n_4035)
);

OR2x2_ASAP7_75t_L g4036 ( 
.A(n_3933),
.B(n_3743),
.Y(n_4036)
);

OA21x2_ASAP7_75t_L g4037 ( 
.A1(n_3911),
.A2(n_3936),
.B(n_3934),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3889),
.B(n_3830),
.Y(n_4038)
);

AND2x4_ASAP7_75t_L g4039 ( 
.A(n_3867),
.B(n_3895),
.Y(n_4039)
);

INVx3_ASAP7_75t_L g4040 ( 
.A(n_3849),
.Y(n_4040)
);

OAI21x1_ASAP7_75t_L g4041 ( 
.A1(n_3882),
.A2(n_3822),
.B(n_3820),
.Y(n_4041)
);

OAI21x1_ASAP7_75t_L g4042 ( 
.A1(n_3967),
.A2(n_3956),
.B(n_3845),
.Y(n_4042)
);

BUFx3_ASAP7_75t_L g4043 ( 
.A(n_3832),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_3858),
.Y(n_4044)
);

AO31x2_ASAP7_75t_L g4045 ( 
.A1(n_3873),
.A2(n_3791),
.A3(n_3782),
.B(n_3794),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3859),
.Y(n_4046)
);

O2A1O1Ixp33_ASAP7_75t_L g4047 ( 
.A1(n_3879),
.A2(n_3739),
.B(n_3736),
.C(n_3774),
.Y(n_4047)
);

OAI21x1_ASAP7_75t_L g4048 ( 
.A1(n_3923),
.A2(n_3827),
.B(n_3823),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3927),
.Y(n_4049)
);

CKINVDCx20_ASAP7_75t_R g4050 ( 
.A(n_3832),
.Y(n_4050)
);

BUFx3_ASAP7_75t_L g4051 ( 
.A(n_3846),
.Y(n_4051)
);

BUFx3_ASAP7_75t_L g4052 ( 
.A(n_3853),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3945),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3872),
.B(n_3684),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3886),
.B(n_3754),
.Y(n_4055)
);

OAI22xp5_ASAP7_75t_SL g4056 ( 
.A1(n_3988),
.A2(n_3776),
.B1(n_3806),
.B2(n_3673),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3937),
.B(n_3830),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3952),
.B(n_3754),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3960),
.Y(n_4059)
);

A2O1A1Ixp33_ASAP7_75t_L g4060 ( 
.A1(n_3942),
.A2(n_3870),
.B(n_3847),
.C(n_3856),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_3924),
.A2(n_3655),
.B(n_3663),
.Y(n_4061)
);

OA21x2_ASAP7_75t_L g4062 ( 
.A1(n_3865),
.A2(n_3686),
.B(n_3689),
.Y(n_4062)
);

BUFx12f_ASAP7_75t_L g4063 ( 
.A(n_3944),
.Y(n_4063)
);

AND2x2_ASAP7_75t_SL g4064 ( 
.A(n_4003),
.B(n_3781),
.Y(n_4064)
);

OAI21x1_ASAP7_75t_L g4065 ( 
.A1(n_3860),
.A2(n_3704),
.B(n_3741),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3925),
.A2(n_3763),
.B(n_3789),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3969),
.B(n_3830),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3848),
.A2(n_3765),
.B1(n_3710),
.B2(n_3726),
.Y(n_4068)
);

OAI21x1_ASAP7_75t_L g4069 ( 
.A1(n_3926),
.A2(n_3747),
.B(n_3771),
.Y(n_4069)
);

INVx4_ASAP7_75t_L g4070 ( 
.A(n_3854),
.Y(n_4070)
);

OAI21x1_ASAP7_75t_L g4071 ( 
.A1(n_3959),
.A2(n_3640),
.B(n_3656),
.Y(n_4071)
);

NOR2xp67_ASAP7_75t_L g4072 ( 
.A(n_3921),
.B(n_3664),
.Y(n_4072)
);

INVx2_ASAP7_75t_L g4073 ( 
.A(n_3863),
.Y(n_4073)
);

AO31x2_ASAP7_75t_L g4074 ( 
.A1(n_3874),
.A2(n_3726),
.A3(n_3743),
.B(n_3656),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3864),
.Y(n_4075)
);

OAI21x1_ASAP7_75t_L g4076 ( 
.A1(n_3948),
.A2(n_3962),
.B(n_3949),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3982),
.Y(n_4077)
);

CKINVDCx11_ASAP7_75t_R g4078 ( 
.A(n_4005),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3989),
.Y(n_4079)
);

AND2x4_ASAP7_75t_L g4080 ( 
.A(n_3861),
.B(n_3726),
.Y(n_4080)
);

AOI21x1_ASAP7_75t_L g4081 ( 
.A1(n_3962),
.A2(n_3754),
.B(n_3801),
.Y(n_4081)
);

AOI21x1_ASAP7_75t_L g4082 ( 
.A1(n_3953),
.A2(n_3754),
.B(n_3801),
.Y(n_4082)
);

BUFx10_ASAP7_75t_L g4083 ( 
.A(n_3983),
.Y(n_4083)
);

OAI21x1_ASAP7_75t_L g4084 ( 
.A1(n_3896),
.A2(n_3754),
.B(n_3801),
.Y(n_4084)
);

OAI21x1_ASAP7_75t_L g4085 ( 
.A1(n_3992),
.A2(n_3801),
.B(n_3752),
.Y(n_4085)
);

OAI21x1_ASAP7_75t_L g4086 ( 
.A1(n_3877),
.A2(n_3752),
.B(n_3714),
.Y(n_4086)
);

AOI21x1_ASAP7_75t_L g4087 ( 
.A1(n_3930),
.A2(n_3752),
.B(n_3714),
.Y(n_4087)
);

OA21x2_ASAP7_75t_L g4088 ( 
.A1(n_4001),
.A2(n_3714),
.B(n_360),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_4012),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3883),
.Y(n_4090)
);

OA21x2_ASAP7_75t_L g4091 ( 
.A1(n_3998),
.A2(n_360),
.B(n_361),
.Y(n_4091)
);

A2O1A1Ixp33_ASAP7_75t_L g4092 ( 
.A1(n_3852),
.A2(n_363),
.B(n_361),
.C(n_362),
.Y(n_4092)
);

AOI21xp33_ASAP7_75t_SL g4093 ( 
.A1(n_3898),
.A2(n_363),
.B(n_364),
.Y(n_4093)
);

OR2x6_ASAP7_75t_L g4094 ( 
.A(n_3861),
.B(n_4003),
.Y(n_4094)
);

INVx3_ASAP7_75t_L g4095 ( 
.A(n_4007),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3893),
.Y(n_4096)
);

BUFx6f_ASAP7_75t_L g4097 ( 
.A(n_3913),
.Y(n_4097)
);

A2O1A1Ixp33_ASAP7_75t_L g4098 ( 
.A1(n_3871),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_4098)
);

NAND2x1_ASAP7_75t_L g4099 ( 
.A(n_3851),
.B(n_365),
.Y(n_4099)
);

OR2x2_ASAP7_75t_L g4100 ( 
.A(n_3955),
.B(n_367),
.Y(n_4100)
);

BUFx2_ASAP7_75t_L g4101 ( 
.A(n_3958),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3931),
.Y(n_4102)
);

O2A1O1Ixp33_ASAP7_75t_L g4103 ( 
.A1(n_3831),
.A2(n_3991),
.B(n_3907),
.C(n_3916),
.Y(n_4103)
);

NAND2x1p5_ASAP7_75t_L g4104 ( 
.A(n_4009),
.B(n_368),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3915),
.Y(n_4105)
);

OAI21x1_ASAP7_75t_L g4106 ( 
.A1(n_3869),
.A2(n_368),
.B(n_369),
.Y(n_4106)
);

INVx1_ASAP7_75t_SL g4107 ( 
.A(n_3984),
.Y(n_4107)
);

AOI21xp33_ASAP7_75t_SL g4108 ( 
.A1(n_3935),
.A2(n_3914),
.B(n_3943),
.Y(n_4108)
);

NAND2x1p5_ASAP7_75t_L g4109 ( 
.A(n_3913),
.B(n_369),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3915),
.Y(n_4110)
);

INVx4_ASAP7_75t_SL g4111 ( 
.A(n_3954),
.Y(n_4111)
);

OAI21x1_ASAP7_75t_L g4112 ( 
.A1(n_3899),
.A2(n_370),
.B(n_371),
.Y(n_4112)
);

OAI21x1_ASAP7_75t_L g4113 ( 
.A1(n_3892),
.A2(n_3839),
.B(n_3912),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4010),
.B(n_370),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3915),
.Y(n_4115)
);

OAI21x1_ASAP7_75t_L g4116 ( 
.A1(n_3950),
.A2(n_371),
.B(n_372),
.Y(n_4116)
);

OAI21x1_ASAP7_75t_L g4117 ( 
.A1(n_3975),
.A2(n_372),
.B(n_373),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_3954),
.Y(n_4118)
);

INVx4_ASAP7_75t_L g4119 ( 
.A(n_3944),
.Y(n_4119)
);

CKINVDCx5p33_ASAP7_75t_R g4120 ( 
.A(n_3965),
.Y(n_4120)
);

OAI21x1_ASAP7_75t_L g4121 ( 
.A1(n_3909),
.A2(n_373),
.B(n_375),
.Y(n_4121)
);

BUFx12f_ASAP7_75t_L g4122 ( 
.A(n_3980),
.Y(n_4122)
);

OA21x2_ASAP7_75t_L g4123 ( 
.A1(n_3900),
.A2(n_3841),
.B(n_3957),
.Y(n_4123)
);

AO21x2_ASAP7_75t_L g4124 ( 
.A1(n_3833),
.A2(n_375),
.B(n_376),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_3964),
.B(n_377),
.Y(n_4125)
);

OR2x2_ASAP7_75t_L g4126 ( 
.A(n_3946),
.B(n_378),
.Y(n_4126)
);

OAI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3938),
.A2(n_378),
.B(n_380),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3929),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_4006),
.A2(n_380),
.B(n_382),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3929),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3929),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_3978),
.A2(n_383),
.B(n_384),
.Y(n_4132)
);

OAI21x1_ASAP7_75t_L g4133 ( 
.A1(n_3836),
.A2(n_385),
.B(n_386),
.Y(n_4133)
);

INVx4_ASAP7_75t_L g4134 ( 
.A(n_3840),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_3954),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3985),
.B(n_3961),
.Y(n_4136)
);

BUFx8_ASAP7_75t_L g4137 ( 
.A(n_3881),
.Y(n_4137)
);

NAND2x1p5_ASAP7_75t_L g4138 ( 
.A(n_3913),
.B(n_385),
.Y(n_4138)
);

NOR4xp25_ASAP7_75t_L g4139 ( 
.A(n_3971),
.B(n_389),
.C(n_387),
.D(n_388),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3985),
.B(n_388),
.Y(n_4140)
);

CKINVDCx5p33_ASAP7_75t_R g4141 ( 
.A(n_3990),
.Y(n_4141)
);

OAI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_3897),
.A2(n_3918),
.B1(n_4002),
.B2(n_3995),
.Y(n_4142)
);

AO21x2_ASAP7_75t_L g4143 ( 
.A1(n_3834),
.A2(n_389),
.B(n_390),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3985),
.B(n_390),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3951),
.Y(n_4145)
);

OAI21x1_ASAP7_75t_L g4146 ( 
.A1(n_3940),
.A2(n_391),
.B(n_392),
.Y(n_4146)
);

BUFx2_ASAP7_75t_L g4147 ( 
.A(n_3993),
.Y(n_4147)
);

OAI21x1_ASAP7_75t_L g4148 ( 
.A1(n_3986),
.A2(n_4004),
.B(n_3974),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3951),
.Y(n_4149)
);

OAI21x1_ASAP7_75t_L g4150 ( 
.A1(n_3963),
.A2(n_393),
.B(n_394),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3951),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3842),
.Y(n_4152)
);

AND2x4_ASAP7_75t_L g4153 ( 
.A(n_3901),
.B(n_393),
.Y(n_4153)
);

INVx3_ASAP7_75t_SL g4154 ( 
.A(n_3901),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3842),
.Y(n_4155)
);

OAI21x1_ASAP7_75t_L g4156 ( 
.A1(n_3939),
.A2(n_395),
.B(n_396),
.Y(n_4156)
);

OAI21x1_ASAP7_75t_L g4157 ( 
.A1(n_3922),
.A2(n_395),
.B(n_396),
.Y(n_4157)
);

INVx4_ASAP7_75t_SL g4158 ( 
.A(n_3842),
.Y(n_4158)
);

AO21x2_ASAP7_75t_L g4159 ( 
.A1(n_3970),
.A2(n_397),
.B(n_398),
.Y(n_4159)
);

BUFx2_ASAP7_75t_L g4160 ( 
.A(n_4000),
.Y(n_4160)
);

AND2x4_ASAP7_75t_L g4161 ( 
.A(n_3906),
.B(n_3996),
.Y(n_4161)
);

AND2x4_ASAP7_75t_L g4162 ( 
.A(n_3884),
.B(n_397),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3905),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3997),
.Y(n_4164)
);

OAI21x1_ASAP7_75t_SL g4165 ( 
.A1(n_3941),
.A2(n_398),
.B(n_400),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4028),
.Y(n_4166)
);

AOI21xp5_ASAP7_75t_L g4167 ( 
.A1(n_4013),
.A2(n_4142),
.B(n_4060),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_4037),
.B(n_3903),
.Y(n_4168)
);

AND2x4_ASAP7_75t_L g4169 ( 
.A(n_4094),
.B(n_3905),
.Y(n_4169)
);

AOI21xp5_ASAP7_75t_L g4170 ( 
.A1(n_4013),
.A2(n_3880),
.B(n_3876),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_4142),
.A2(n_3875),
.B(n_3917),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4037),
.B(n_3905),
.Y(n_4172)
);

BUFx6f_ASAP7_75t_L g4173 ( 
.A(n_4043),
.Y(n_4173)
);

AND2x4_ASAP7_75t_L g4174 ( 
.A(n_4094),
.B(n_3977),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_4107),
.B(n_3977),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_4096),
.B(n_3977),
.Y(n_4176)
);

OAI21x1_ASAP7_75t_L g4177 ( 
.A1(n_4118),
.A2(n_3999),
.B(n_3904),
.Y(n_4177)
);

AO21x1_ASAP7_75t_L g4178 ( 
.A1(n_4152),
.A2(n_3890),
.B(n_3908),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4053),
.B(n_3902),
.Y(n_4179)
);

OAI21xp33_ASAP7_75t_SL g4180 ( 
.A1(n_4094),
.A2(n_3979),
.B(n_3838),
.Y(n_4180)
);

OA21x2_ASAP7_75t_L g4181 ( 
.A1(n_4135),
.A2(n_3947),
.B(n_3981),
.Y(n_4181)
);

AOI21xp5_ASAP7_75t_L g4182 ( 
.A1(n_4060),
.A2(n_3973),
.B(n_4011),
.Y(n_4182)
);

NAND2x1p5_ASAP7_75t_L g4183 ( 
.A(n_4064),
.B(n_4072),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4049),
.Y(n_4184)
);

OA21x2_ASAP7_75t_L g4185 ( 
.A1(n_4155),
.A2(n_3968),
.B(n_3878),
.Y(n_4185)
);

NAND2x1p5_ASAP7_75t_L g4186 ( 
.A(n_4072),
.B(n_3837),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4014),
.Y(n_4187)
);

AO21x2_ASAP7_75t_L g4188 ( 
.A1(n_4136),
.A2(n_3994),
.B(n_3987),
.Y(n_4188)
);

AO31x2_ASAP7_75t_L g4189 ( 
.A1(n_4136),
.A2(n_3837),
.A3(n_3894),
.B(n_3843),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_4088),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_4039),
.B(n_3837),
.Y(n_4191)
);

AO21x2_ASAP7_75t_L g4192 ( 
.A1(n_4140),
.A2(n_3894),
.B(n_3843),
.Y(n_4192)
);

INVx1_ASAP7_75t_SL g4193 ( 
.A(n_4024),
.Y(n_4193)
);

AOI22x1_ASAP7_75t_L g4194 ( 
.A1(n_4089),
.A2(n_3894),
.B1(n_3910),
.B2(n_3843),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_4088),
.Y(n_4195)
);

CKINVDCx5p33_ASAP7_75t_R g4196 ( 
.A(n_4050),
.Y(n_4196)
);

AOI21x1_ASAP7_75t_L g4197 ( 
.A1(n_4081),
.A2(n_3910),
.B(n_401),
.Y(n_4197)
);

AND2x4_ASAP7_75t_L g4198 ( 
.A(n_4111),
.B(n_3910),
.Y(n_4198)
);

OAI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_4134),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_4199)
);

HB1xp67_ASAP7_75t_L g4200 ( 
.A(n_4026),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4028),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4018),
.Y(n_4202)
);

AO21x2_ASAP7_75t_L g4203 ( 
.A1(n_4140),
.A2(n_404),
.B(n_405),
.Y(n_4203)
);

A2O1A1Ixp33_ASAP7_75t_L g4204 ( 
.A1(n_4103),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4021),
.Y(n_4205)
);

AO31x2_ASAP7_75t_L g4206 ( 
.A1(n_4067),
.A2(n_410),
.A3(n_408),
.B(n_409),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_4059),
.Y(n_4207)
);

AOI21xp5_ASAP7_75t_L g4208 ( 
.A1(n_4129),
.A2(n_408),
.B(n_409),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4161),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_4129),
.A2(n_411),
.B(n_412),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_4070),
.B(n_412),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4077),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4057),
.B(n_413),
.Y(n_4213)
);

AOI21xp5_ASAP7_75t_L g4214 ( 
.A1(n_4029),
.A2(n_4103),
.B(n_4139),
.Y(n_4214)
);

OR2x2_ASAP7_75t_L g4215 ( 
.A(n_4107),
.B(n_413),
.Y(n_4215)
);

OA21x2_ASAP7_75t_L g4216 ( 
.A1(n_4057),
.A2(n_414),
.B(n_415),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4079),
.Y(n_4217)
);

HB1xp67_ASAP7_75t_L g4218 ( 
.A(n_4026),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4161),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_4029),
.A2(n_414),
.B(n_415),
.Y(n_4220)
);

OA21x2_ASAP7_75t_L g4221 ( 
.A1(n_4067),
.A2(n_416),
.B(n_417),
.Y(n_4221)
);

OA21x2_ASAP7_75t_L g4222 ( 
.A1(n_4023),
.A2(n_416),
.B(n_417),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_4111),
.B(n_420),
.Y(n_4223)
);

INVx5_ASAP7_75t_L g4224 ( 
.A(n_4089),
.Y(n_4224)
);

OAI21x1_ASAP7_75t_L g4225 ( 
.A1(n_4019),
.A2(n_421),
.B(n_422),
.Y(n_4225)
);

OA21x2_ASAP7_75t_L g4226 ( 
.A1(n_4035),
.A2(n_4038),
.B(n_4017),
.Y(n_4226)
);

AO21x2_ASAP7_75t_L g4227 ( 
.A1(n_4144),
.A2(n_421),
.B(n_422),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4015),
.B(n_423),
.Y(n_4228)
);

A2O1A1Ixp33_ASAP7_75t_L g4229 ( 
.A1(n_4108),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_4229)
);

AND2x2_ASAP7_75t_L g4230 ( 
.A(n_4039),
.B(n_426),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_4030),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4015),
.B(n_426),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_SL g4233 ( 
.A(n_4119),
.B(n_427),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4139),
.A2(n_427),
.B(n_428),
.Y(n_4234)
);

BUFx2_ASAP7_75t_R g4235 ( 
.A(n_4141),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4044),
.Y(n_4236)
);

OAI21x1_ASAP7_75t_SL g4237 ( 
.A1(n_4119),
.A2(n_428),
.B(n_429),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_4144),
.A2(n_429),
.B(n_430),
.Y(n_4238)
);

NAND2x1p5_ASAP7_75t_L g4239 ( 
.A(n_4153),
.B(n_430),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4054),
.B(n_431),
.Y(n_4240)
);

AOI21x1_ASAP7_75t_L g4241 ( 
.A1(n_4087),
.A2(n_4101),
.B(n_4082),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4158),
.B(n_431),
.Y(n_4242)
);

OAI21x1_ASAP7_75t_L g4243 ( 
.A1(n_4019),
.A2(n_432),
.B(n_433),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4035),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4038),
.Y(n_4245)
);

OAI21x1_ASAP7_75t_L g4246 ( 
.A1(n_4085),
.A2(n_432),
.B(n_435),
.Y(n_4246)
);

INVx4_ASAP7_75t_L g4247 ( 
.A(n_4089),
.Y(n_4247)
);

OAI21x1_ASAP7_75t_L g4248 ( 
.A1(n_4036),
.A2(n_4031),
.B(n_4076),
.Y(n_4248)
);

AND2x4_ASAP7_75t_L g4249 ( 
.A(n_4111),
.B(n_435),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4158),
.B(n_436),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4163),
.Y(n_4251)
);

OAI21x1_ASAP7_75t_SL g4252 ( 
.A1(n_4134),
.A2(n_436),
.B(n_437),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_SL g4253 ( 
.A1(n_4091),
.A2(n_438),
.B(n_439),
.Y(n_4253)
);

CKINVDCx5p33_ASAP7_75t_R g4254 ( 
.A(n_4120),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_4020),
.A2(n_438),
.B(n_440),
.Y(n_4255)
);

INVx3_ASAP7_75t_L g4256 ( 
.A(n_4070),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_4095),
.B(n_441),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4105),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4046),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4158),
.B(n_441),
.Y(n_4260)
);

OAI21x1_ASAP7_75t_L g4261 ( 
.A1(n_4031),
.A2(n_442),
.B(n_443),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4110),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4123),
.B(n_443),
.Y(n_4263)
);

OAI21x1_ASAP7_75t_L g4264 ( 
.A1(n_4115),
.A2(n_444),
.B(n_446),
.Y(n_4264)
);

HB1xp67_ASAP7_75t_L g4265 ( 
.A(n_4091),
.Y(n_4265)
);

AO21x2_ASAP7_75t_L g4266 ( 
.A1(n_4128),
.A2(n_447),
.B(n_448),
.Y(n_4266)
);

AOI22xp33_ASAP7_75t_L g4267 ( 
.A1(n_4080),
.A2(n_4078),
.B1(n_4143),
.B2(n_4124),
.Y(n_4267)
);

INVx3_ASAP7_75t_L g4268 ( 
.A(n_4063),
.Y(n_4268)
);

NOR2xp33_ASAP7_75t_R g4269 ( 
.A(n_4034),
.B(n_447),
.Y(n_4269)
);

AOI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_4124),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_4270)
);

AO21x2_ASAP7_75t_L g4271 ( 
.A1(n_4130),
.A2(n_449),
.B(n_451),
.Y(n_4271)
);

AO31x2_ASAP7_75t_L g4272 ( 
.A1(n_4131),
.A2(n_454),
.A3(n_452),
.B(n_453),
.Y(n_4272)
);

INVx4_ASAP7_75t_L g4273 ( 
.A(n_4104),
.Y(n_4273)
);

OAI21x1_ASAP7_75t_L g4274 ( 
.A1(n_4145),
.A2(n_452),
.B(n_454),
.Y(n_4274)
);

BUFx2_ASAP7_75t_R g4275 ( 
.A(n_4051),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4095),
.B(n_455),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4149),
.Y(n_4277)
);

HB1xp67_ASAP7_75t_L g4278 ( 
.A(n_4123),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4151),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4090),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4080),
.B(n_4062),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_4020),
.A2(n_455),
.B(n_456),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4073),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4025),
.B(n_456),
.Y(n_4284)
);

AOI21xp5_ASAP7_75t_L g4285 ( 
.A1(n_4132),
.A2(n_457),
.B(n_458),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4132),
.A2(n_457),
.B(n_458),
.Y(n_4286)
);

AOI21x1_ASAP7_75t_L g4287 ( 
.A1(n_4147),
.A2(n_459),
.B(n_460),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_4092),
.A2(n_460),
.B(n_462),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4062),
.B(n_463),
.Y(n_4289)
);

AOI21xp5_ASAP7_75t_L g4290 ( 
.A1(n_4092),
.A2(n_464),
.B(n_465),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4164),
.B(n_465),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4075),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4102),
.B(n_466),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_4160),
.B(n_466),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4025),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_4055),
.B(n_467),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4086),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_4100),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4074),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_SL g4300 ( 
.A(n_4052),
.B(n_467),
.Y(n_4300)
);

OAI21x1_ASAP7_75t_L g4301 ( 
.A1(n_4040),
.A2(n_468),
.B(n_469),
.Y(n_4301)
);

BUFx8_ASAP7_75t_L g4302 ( 
.A(n_4125),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_4114),
.B(n_469),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4074),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_4122),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_4042),
.Y(n_4306)
);

INVxp33_ASAP7_75t_L g4307 ( 
.A(n_4099),
.Y(n_4307)
);

AOI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_4108),
.A2(n_4084),
.B(n_4056),
.Y(n_4308)
);

OAI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4093),
.A2(n_4098),
.B(n_4113),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4027),
.Y(n_4310)
);

AO21x2_ASAP7_75t_L g4311 ( 
.A1(n_4093),
.A2(n_470),
.B(n_471),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4032),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4069),
.Y(n_4313)
);

AO31x2_ASAP7_75t_L g4314 ( 
.A1(n_4098),
.A2(n_472),
.A3(n_470),
.B(n_471),
.Y(n_4314)
);

OR2x2_ASAP7_75t_L g4315 ( 
.A(n_4040),
.B(n_472),
.Y(n_4315)
);

A2O1A1Ixp33_ASAP7_75t_L g4316 ( 
.A1(n_4047),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_4316)
);

AOI22xp33_ASAP7_75t_SL g4317 ( 
.A1(n_4168),
.A2(n_4162),
.B1(n_4159),
.B2(n_4165),
.Y(n_4317)
);

CKINVDCx5p33_ASAP7_75t_R g4318 ( 
.A(n_4196),
.Y(n_4318)
);

OAI22xp5_ASAP7_75t_L g4319 ( 
.A1(n_4167),
.A2(n_4154),
.B1(n_4056),
.B2(n_4068),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_4178),
.A2(n_4159),
.B1(n_4143),
.B2(n_4068),
.Y(n_4320)
);

OAI21xp33_ASAP7_75t_L g4321 ( 
.A1(n_4214),
.A2(n_4022),
.B(n_4104),
.Y(n_4321)
);

HB1xp67_ASAP7_75t_L g4322 ( 
.A(n_4222),
.Y(n_4322)
);

AOI22xp33_ASAP7_75t_L g4323 ( 
.A1(n_4192),
.A2(n_4162),
.B1(n_4022),
.B2(n_4148),
.Y(n_4323)
);

AOI22xp33_ASAP7_75t_L g4324 ( 
.A1(n_4192),
.A2(n_4133),
.B1(n_4121),
.B2(n_4146),
.Y(n_4324)
);

OAI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_4182),
.A2(n_4126),
.B1(n_4138),
.B2(n_4109),
.Y(n_4325)
);

NOR2xp33_ASAP7_75t_L g4326 ( 
.A(n_4235),
.B(n_4083),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_SL g4327 ( 
.A1(n_4171),
.A2(n_4047),
.B(n_4016),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4187),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_4191),
.B(n_4058),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4202),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4186),
.Y(n_4331)
);

AOI222xp33_ASAP7_75t_L g4332 ( 
.A1(n_4309),
.A2(n_4153),
.B1(n_4150),
.B2(n_4083),
.C1(n_4112),
.C2(n_4157),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4190),
.Y(n_4333)
);

CKINVDCx20_ASAP7_75t_R g4334 ( 
.A(n_4302),
.Y(n_4334)
);

BUFx12f_ASAP7_75t_L g4335 ( 
.A(n_4173),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4205),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_SL g4337 ( 
.A1(n_4194),
.A2(n_4137),
.B1(n_4138),
.B2(n_4109),
.Y(n_4337)
);

AOI22xp5_ASAP7_75t_L g4338 ( 
.A1(n_4170),
.A2(n_4065),
.B1(n_4127),
.B2(n_4156),
.Y(n_4338)
);

CKINVDCx5p33_ASAP7_75t_R g4339 ( 
.A(n_4254),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4195),
.Y(n_4340)
);

AOI22xp5_ASAP7_75t_L g4341 ( 
.A1(n_4188),
.A2(n_4117),
.B1(n_4066),
.B2(n_4137),
.Y(n_4341)
);

AOI22xp33_ASAP7_75t_L g4342 ( 
.A1(n_4188),
.A2(n_4106),
.B1(n_4116),
.B2(n_4061),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4229),
.A2(n_4016),
.B1(n_4097),
.B2(n_4045),
.Y(n_4343)
);

AOI22xp33_ASAP7_75t_L g4344 ( 
.A1(n_4185),
.A2(n_4041),
.B1(n_4097),
.B2(n_4048),
.Y(n_4344)
);

AOI22xp33_ASAP7_75t_SL g4345 ( 
.A1(n_4278),
.A2(n_4074),
.B1(n_4097),
.B2(n_4045),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_SL g4346 ( 
.A(n_4183),
.B(n_4071),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4223),
.Y(n_4347)
);

OAI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_4172),
.A2(n_4045),
.B1(n_4033),
.B2(n_476),
.Y(n_4348)
);

OAI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4265),
.A2(n_477),
.B1(n_473),
.B2(n_475),
.Y(n_4349)
);

OAI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4289),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_4350)
);

OAI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_4204),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_4351)
);

AOI22xp33_ASAP7_75t_L g4352 ( 
.A1(n_4185),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_4352)
);

AOI22xp5_ASAP7_75t_L g4353 ( 
.A1(n_4180),
.A2(n_485),
.B1(n_481),
.B2(n_483),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4255),
.A2(n_488),
.B1(n_485),
.B2(n_486),
.Y(n_4354)
);

OR2x2_ASAP7_75t_L g4355 ( 
.A(n_4298),
.B(n_486),
.Y(n_4355)
);

OAI21xp33_ASAP7_75t_L g4356 ( 
.A1(n_4176),
.A2(n_489),
.B(n_490),
.Y(n_4356)
);

AOI22xp33_ASAP7_75t_L g4357 ( 
.A1(n_4181),
.A2(n_490),
.B1(n_491),
.B2(n_492),
.Y(n_4357)
);

AOI22xp33_ASAP7_75t_L g4358 ( 
.A1(n_4181),
.A2(n_491),
.B1(n_492),
.B2(n_493),
.Y(n_4358)
);

OAI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4282),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_4359)
);

AOI22xp33_ASAP7_75t_L g4360 ( 
.A1(n_4234),
.A2(n_4267),
.B1(n_4284),
.B2(n_4174),
.Y(n_4360)
);

BUFx4f_ASAP7_75t_SL g4361 ( 
.A(n_4173),
.Y(n_4361)
);

AOI222xp33_ASAP7_75t_L g4362 ( 
.A1(n_4179),
.A2(n_494),
.B1(n_496),
.B2(n_497),
.C1(n_498),
.C2(n_500),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4256),
.B(n_496),
.Y(n_4363)
);

OAI222xp33_ASAP7_75t_L g4364 ( 
.A1(n_4175),
.A2(n_497),
.B1(n_500),
.B2(n_501),
.C1(n_502),
.C2(n_503),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4263),
.B(n_502),
.Y(n_4365)
);

BUFx3_ASAP7_75t_L g4366 ( 
.A(n_4302),
.Y(n_4366)
);

AND2x4_ASAP7_75t_L g4367 ( 
.A(n_4256),
.B(n_503),
.Y(n_4367)
);

BUFx2_ASAP7_75t_L g4368 ( 
.A(n_4268),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4280),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_4275),
.B(n_504),
.Y(n_4370)
);

AOI22xp33_ASAP7_75t_L g4371 ( 
.A1(n_4284),
.A2(n_505),
.B1(n_507),
.B2(n_509),
.Y(n_4371)
);

AOI22xp33_ASAP7_75t_SL g4372 ( 
.A1(n_4198),
.A2(n_505),
.B1(n_507),
.B2(n_509),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4184),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4221),
.B(n_510),
.Y(n_4374)
);

INVx5_ASAP7_75t_SL g4375 ( 
.A(n_4173),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_4174),
.A2(n_510),
.B1(n_512),
.B2(n_513),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_SL g4377 ( 
.A1(n_4198),
.A2(n_4169),
.B1(n_4216),
.B2(n_4221),
.Y(n_4377)
);

BUFx2_ASAP7_75t_L g4378 ( 
.A(n_4268),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4169),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4273),
.B(n_515),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4223),
.Y(n_4381)
);

INVx4_ASAP7_75t_L g4382 ( 
.A(n_4224),
.Y(n_4382)
);

AOI22xp33_ASAP7_75t_L g4383 ( 
.A1(n_4216),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.Y(n_4383)
);

OAI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_4316),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4189),
.B(n_518),
.Y(n_4385)
);

AOI22xp33_ASAP7_75t_SL g4386 ( 
.A1(n_4281),
.A2(n_520),
.B1(n_522),
.B2(n_523),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_4222),
.A2(n_520),
.B1(n_524),
.B2(n_525),
.Y(n_4387)
);

NOR2xp33_ASAP7_75t_L g4388 ( 
.A(n_4247),
.B(n_4193),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_4269),
.Y(n_4389)
);

AOI22xp33_ASAP7_75t_SL g4390 ( 
.A1(n_4203),
.A2(n_524),
.B1(n_526),
.B2(n_527),
.Y(n_4390)
);

INVxp67_ASAP7_75t_L g4391 ( 
.A(n_4242),
.Y(n_4391)
);

OAI21xp33_ASAP7_75t_L g4392 ( 
.A1(n_4313),
.A2(n_4308),
.B(n_4306),
.Y(n_4392)
);

OAI222xp33_ASAP7_75t_L g4393 ( 
.A1(n_4270),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.C1(n_529),
.C2(n_530),
.Y(n_4393)
);

AND2x2_ASAP7_75t_L g4394 ( 
.A(n_4273),
.B(n_528),
.Y(n_4394)
);

INVx1_ASAP7_75t_SL g4395 ( 
.A(n_4250),
.Y(n_4395)
);

INVx3_ASAP7_75t_L g4396 ( 
.A(n_4247),
.Y(n_4396)
);

OAI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_4307),
.A2(n_529),
.B1(n_531),
.B2(n_534),
.Y(n_4397)
);

NOR2xp33_ASAP7_75t_L g4398 ( 
.A(n_4224),
.B(n_531),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_L g4399 ( 
.A1(n_4288),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4207),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4249),
.Y(n_4401)
);

AOI22xp33_ASAP7_75t_L g4402 ( 
.A1(n_4290),
.A2(n_536),
.B1(n_537),
.B2(n_538),
.Y(n_4402)
);

OAI21xp33_ASAP7_75t_L g4403 ( 
.A1(n_4310),
.A2(n_4312),
.B(n_4253),
.Y(n_4403)
);

OAI22xp5_ASAP7_75t_L g4404 ( 
.A1(n_4213),
.A2(n_537),
.B1(n_538),
.B2(n_539),
.Y(n_4404)
);

AOI22xp5_ASAP7_75t_L g4405 ( 
.A1(n_4203),
.A2(n_539),
.B1(n_541),
.B2(n_542),
.Y(n_4405)
);

OAI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4215),
.A2(n_541),
.B1(n_542),
.B2(n_543),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4212),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_4305),
.Y(n_4408)
);

OAI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_4224),
.A2(n_4260),
.B1(n_4315),
.B2(n_4249),
.Y(n_4409)
);

HB1xp67_ASAP7_75t_L g4410 ( 
.A(n_4217),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4227),
.A2(n_544),
.B1(n_545),
.B2(n_546),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4206),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4206),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4206),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4228),
.A2(n_544),
.B1(n_545),
.B2(n_546),
.Y(n_4415)
);

AOI22xp33_ASAP7_75t_SL g4416 ( 
.A1(n_4227),
.A2(n_547),
.B1(n_548),
.B2(n_549),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4189),
.B(n_547),
.Y(n_4417)
);

AOI22xp33_ASAP7_75t_SL g4418 ( 
.A1(n_4266),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_4230),
.B(n_550),
.Y(n_4419)
);

OAI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4209),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.Y(n_4420)
);

BUFx3_ASAP7_75t_L g4421 ( 
.A(n_4239),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4219),
.Y(n_4422)
);

CKINVDCx20_ASAP7_75t_R g4423 ( 
.A(n_4240),
.Y(n_4423)
);

OAI21xp5_ASAP7_75t_SL g4424 ( 
.A1(n_4220),
.A2(n_551),
.B(n_552),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_4297),
.Y(n_4425)
);

OAI222xp33_ASAP7_75t_L g4426 ( 
.A1(n_4238),
.A2(n_553),
.B1(n_555),
.B2(n_557),
.C1(n_558),
.C2(n_559),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_L g4427 ( 
.A1(n_4266),
.A2(n_4271),
.B1(n_4304),
.B2(n_4299),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4241),
.B(n_557),
.Y(n_4428)
);

AOI22xp33_ASAP7_75t_L g4429 ( 
.A1(n_4271),
.A2(n_558),
.B1(n_560),
.B2(n_561),
.Y(n_4429)
);

INVx3_ASAP7_75t_L g4430 ( 
.A(n_4248),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4177),
.Y(n_4431)
);

AO22x1_ASAP7_75t_L g4432 ( 
.A1(n_4257),
.A2(n_560),
.B1(n_561),
.B2(n_562),
.Y(n_4432)
);

AOI22xp33_ASAP7_75t_SL g4433 ( 
.A1(n_4300),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4433)
);

AOI22xp33_ASAP7_75t_SL g4434 ( 
.A1(n_4226),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4258),
.Y(n_4435)
);

AOI21xp5_ASAP7_75t_SL g4436 ( 
.A1(n_4296),
.A2(n_566),
.B(n_567),
.Y(n_4436)
);

AOI22xp33_ASAP7_75t_L g4437 ( 
.A1(n_4285),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.Y(n_4437)
);

OAI22xp5_ASAP7_75t_L g4438 ( 
.A1(n_4232),
.A2(n_570),
.B1(n_571),
.B2(n_572),
.Y(n_4438)
);

OAI22xp5_ASAP7_75t_L g4439 ( 
.A1(n_4208),
.A2(n_4210),
.B1(n_4286),
.B2(n_4293),
.Y(n_4439)
);

CKINVDCx16_ASAP7_75t_R g4440 ( 
.A(n_4294),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4246),
.Y(n_4441)
);

INVxp67_ASAP7_75t_SL g4442 ( 
.A(n_4226),
.Y(n_4442)
);

OR2x2_ASAP7_75t_L g4443 ( 
.A(n_4189),
.B(n_573),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4258),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_4236),
.Y(n_4445)
);

BUFx6f_ASAP7_75t_L g4446 ( 
.A(n_4287),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_SL g4447 ( 
.A(n_4291),
.B(n_573),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4200),
.B(n_4218),
.Y(n_4448)
);

AOI22xp5_ASAP7_75t_L g4449 ( 
.A1(n_4311),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.Y(n_4449)
);

CKINVDCx5p33_ASAP7_75t_R g4450 ( 
.A(n_4211),
.Y(n_4450)
);

HB1xp67_ASAP7_75t_L g4451 ( 
.A(n_4310),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_4259),
.Y(n_4452)
);

AOI22xp5_ASAP7_75t_L g4453 ( 
.A1(n_4311),
.A2(n_574),
.B1(n_575),
.B2(n_577),
.Y(n_4453)
);

AOI22xp33_ASAP7_75t_SL g4454 ( 
.A1(n_4295),
.A2(n_577),
.B1(n_578),
.B2(n_579),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4262),
.Y(n_4455)
);

INVx3_ASAP7_75t_L g4456 ( 
.A(n_4312),
.Y(n_4456)
);

BUFx6f_ASAP7_75t_L g4457 ( 
.A(n_4264),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4262),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4251),
.Y(n_4459)
);

OAI22xp5_ASAP7_75t_L g4460 ( 
.A1(n_4199),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.Y(n_4460)
);

AOI22xp33_ASAP7_75t_SL g4461 ( 
.A1(n_4295),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_4461)
);

OAI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4233),
.A2(n_582),
.B1(n_583),
.B2(n_584),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4283),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4251),
.Y(n_4464)
);

INVx2_ASAP7_75t_L g4465 ( 
.A(n_4292),
.Y(n_4465)
);

HB1xp67_ASAP7_75t_L g4466 ( 
.A(n_4166),
.Y(n_4466)
);

HB1xp67_ASAP7_75t_L g4467 ( 
.A(n_4166),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4276),
.B(n_583),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_4443),
.Y(n_4469)
);

HB1xp67_ASAP7_75t_L g4470 ( 
.A(n_4322),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4317),
.B(n_4395),
.Y(n_4471)
);

AOI21x1_ASAP7_75t_L g4472 ( 
.A1(n_4428),
.A2(n_4303),
.B(n_4197),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4329),
.B(n_4201),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4410),
.Y(n_4474)
);

INVx2_ASAP7_75t_L g4475 ( 
.A(n_4457),
.Y(n_4475)
);

AO21x2_ASAP7_75t_L g4476 ( 
.A1(n_4385),
.A2(n_4201),
.B(n_4244),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4417),
.Y(n_4477)
);

INVxp33_ASAP7_75t_L g4478 ( 
.A(n_4326),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4328),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4396),
.B(n_4244),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4330),
.Y(n_4481)
);

OR2x6_ASAP7_75t_L g4482 ( 
.A(n_4382),
.B(n_4252),
.Y(n_4482)
);

AO31x2_ASAP7_75t_L g4483 ( 
.A1(n_4412),
.A2(n_4279),
.A3(n_4277),
.B(n_4245),
.Y(n_4483)
);

BUFx3_ASAP7_75t_L g4484 ( 
.A(n_4334),
.Y(n_4484)
);

AND2x4_ASAP7_75t_L g4485 ( 
.A(n_4368),
.B(n_4245),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4336),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4457),
.Y(n_4487)
);

AO21x2_ASAP7_75t_L g4488 ( 
.A1(n_4442),
.A2(n_4237),
.B(n_4274),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4457),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4373),
.Y(n_4490)
);

AND3x2_ASAP7_75t_L g4491 ( 
.A(n_4436),
.B(n_4231),
.C(n_4243),
.Y(n_4491)
);

OR2x6_ASAP7_75t_L g4492 ( 
.A(n_4382),
.B(n_4225),
.Y(n_4492)
);

BUFx3_ASAP7_75t_L g4493 ( 
.A(n_4366),
.Y(n_4493)
);

HB1xp67_ASAP7_75t_L g4494 ( 
.A(n_4441),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4400),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4446),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4396),
.B(n_4301),
.Y(n_4497)
);

HB1xp67_ASAP7_75t_L g4498 ( 
.A(n_4407),
.Y(n_4498)
);

AO21x2_ASAP7_75t_L g4499 ( 
.A1(n_4392),
.A2(n_4261),
.B(n_4272),
.Y(n_4499)
);

AND2x4_ASAP7_75t_L g4500 ( 
.A(n_4378),
.B(n_4272),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4395),
.B(n_4314),
.Y(n_4501)
);

HB1xp67_ASAP7_75t_L g4502 ( 
.A(n_4446),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4446),
.Y(n_4503)
);

AND2x4_ASAP7_75t_L g4504 ( 
.A(n_4331),
.B(n_4272),
.Y(n_4504)
);

HB1xp67_ASAP7_75t_L g4505 ( 
.A(n_4451),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4369),
.Y(n_4506)
);

INVx2_ASAP7_75t_L g4507 ( 
.A(n_4456),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4374),
.Y(n_4508)
);

INVx3_ASAP7_75t_L g4509 ( 
.A(n_4335),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_4431),
.B(n_4314),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4435),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_4448),
.B(n_4314),
.Y(n_4512)
);

INVxp67_ASAP7_75t_L g4513 ( 
.A(n_4388),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4444),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4455),
.Y(n_4515)
);

HB1xp67_ASAP7_75t_L g4516 ( 
.A(n_4466),
.Y(n_4516)
);

BUFx4f_ASAP7_75t_SL g4517 ( 
.A(n_4367),
.Y(n_4517)
);

INVx3_ASAP7_75t_L g4518 ( 
.A(n_4375),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4456),
.Y(n_4519)
);

BUFx2_ASAP7_75t_L g4520 ( 
.A(n_4408),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4467),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4333),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4458),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4340),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_4413),
.Y(n_4525)
);

HB1xp67_ASAP7_75t_L g4526 ( 
.A(n_4391),
.Y(n_4526)
);

AO21x2_ASAP7_75t_L g4527 ( 
.A1(n_4348),
.A2(n_584),
.B(n_585),
.Y(n_4527)
);

INVx1_ASAP7_75t_SL g4528 ( 
.A(n_4423),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_4414),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_4422),
.Y(n_4530)
);

AND2x4_ASAP7_75t_L g4531 ( 
.A(n_4347),
.B(n_586),
.Y(n_4531)
);

OA21x2_ASAP7_75t_L g4532 ( 
.A1(n_4327),
.A2(n_587),
.B(n_589),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4459),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4464),
.Y(n_4534)
);

HB1xp67_ASAP7_75t_L g4535 ( 
.A(n_4439),
.Y(n_4535)
);

AO21x2_ASAP7_75t_L g4536 ( 
.A1(n_4365),
.A2(n_587),
.B(n_589),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4440),
.B(n_590),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4355),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4425),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4344),
.B(n_590),
.Y(n_4540)
);

AND2x4_ASAP7_75t_L g4541 ( 
.A(n_4381),
.B(n_591),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4375),
.B(n_592),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4375),
.B(n_592),
.Y(n_4543)
);

NOR3xp33_ASAP7_75t_L g4544 ( 
.A(n_4343),
.B(n_594),
.C(n_595),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4338),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4380),
.Y(n_4546)
);

INVx3_ASAP7_75t_L g4547 ( 
.A(n_4430),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_4394),
.Y(n_4548)
);

HB1xp67_ASAP7_75t_L g4549 ( 
.A(n_4439),
.Y(n_4549)
);

AO21x2_ASAP7_75t_L g4550 ( 
.A1(n_4403),
.A2(n_594),
.B(n_596),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4405),
.Y(n_4551)
);

HB1xp67_ASAP7_75t_L g4552 ( 
.A(n_4343),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4360),
.B(n_596),
.Y(n_4553)
);

NOR2xp33_ASAP7_75t_L g4554 ( 
.A(n_4361),
.B(n_597),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4341),
.B(n_598),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4409),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4401),
.Y(n_4557)
);

OA21x2_ASAP7_75t_L g4558 ( 
.A1(n_4321),
.A2(n_599),
.B(n_600),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4445),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4346),
.B(n_4323),
.Y(n_4560)
);

OR2x2_ASAP7_75t_L g4561 ( 
.A(n_4342),
.B(n_599),
.Y(n_4561)
);

AO21x2_ASAP7_75t_L g4562 ( 
.A1(n_4319),
.A2(n_602),
.B(n_603),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4452),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4325),
.Y(n_4564)
);

HB1xp67_ASAP7_75t_L g4565 ( 
.A(n_4397),
.Y(n_4565)
);

AO21x2_ASAP7_75t_L g4566 ( 
.A1(n_4349),
.A2(n_603),
.B(n_604),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_4363),
.Y(n_4567)
);

INVx3_ASAP7_75t_L g4568 ( 
.A(n_4430),
.Y(n_4568)
);

INVxp67_ASAP7_75t_L g4569 ( 
.A(n_4370),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4463),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4325),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4465),
.Y(n_4572)
);

BUFx6f_ASAP7_75t_L g4573 ( 
.A(n_4367),
.Y(n_4573)
);

AOI222xp33_ASAP7_75t_L g4574 ( 
.A1(n_4320),
.A2(n_690),
.B1(n_605),
.B2(n_606),
.C1(n_608),
.C2(n_610),
.Y(n_4574)
);

OR2x6_ASAP7_75t_L g4575 ( 
.A(n_4432),
.B(n_604),
.Y(n_4575)
);

NOR2xp33_ASAP7_75t_L g4576 ( 
.A(n_4450),
.B(n_605),
.Y(n_4576)
);

INVx2_ASAP7_75t_SL g4577 ( 
.A(n_4421),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4449),
.Y(n_4578)
);

BUFx6f_ASAP7_75t_L g4579 ( 
.A(n_4398),
.Y(n_4579)
);

AO21x2_ASAP7_75t_L g4580 ( 
.A1(n_4350),
.A2(n_608),
.B(n_610),
.Y(n_4580)
);

OA21x2_ASAP7_75t_L g4581 ( 
.A1(n_4427),
.A2(n_611),
.B(n_612),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4453),
.Y(n_4582)
);

AO21x2_ASAP7_75t_L g4583 ( 
.A1(n_4353),
.A2(n_611),
.B(n_613),
.Y(n_4583)
);

HB1xp67_ASAP7_75t_L g4584 ( 
.A(n_4332),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4434),
.B(n_613),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4468),
.Y(n_4586)
);

HB1xp67_ASAP7_75t_L g4587 ( 
.A(n_4332),
.Y(n_4587)
);

OR2x2_ASAP7_75t_L g4588 ( 
.A(n_4324),
.B(n_614),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4419),
.Y(n_4589)
);

HB1xp67_ASAP7_75t_L g4590 ( 
.A(n_4438),
.Y(n_4590)
);

OA21x2_ASAP7_75t_L g4591 ( 
.A1(n_4356),
.A2(n_614),
.B(n_615),
.Y(n_4591)
);

INVx3_ASAP7_75t_L g4592 ( 
.A(n_4318),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4377),
.B(n_615),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4447),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4345),
.B(n_616),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4406),
.Y(n_4596)
);

INVx4_ASAP7_75t_L g4597 ( 
.A(n_4339),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4406),
.Y(n_4598)
);

OAI21xp33_ASAP7_75t_SL g4599 ( 
.A1(n_4362),
.A2(n_690),
.B(n_617),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4357),
.B(n_616),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4438),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4404),
.Y(n_4602)
);

BUFx2_ASAP7_75t_L g4603 ( 
.A(n_4389),
.Y(n_4603)
);

AOI22xp33_ASAP7_75t_L g4604 ( 
.A1(n_4351),
.A2(n_618),
.B1(n_619),
.B2(n_620),
.Y(n_4604)
);

NAND2x1_ASAP7_75t_L g4605 ( 
.A(n_4379),
.B(n_619),
.Y(n_4605)
);

AO21x2_ASAP7_75t_L g4606 ( 
.A1(n_4364),
.A2(n_620),
.B(n_621),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4470),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4525),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4525),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4535),
.B(n_4337),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4549),
.B(n_4358),
.Y(n_4611)
);

NAND2x1_ASAP7_75t_L g4612 ( 
.A(n_4573),
.B(n_4352),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4577),
.B(n_4386),
.Y(n_4613)
);

AND2x2_ASAP7_75t_L g4614 ( 
.A(n_4577),
.B(n_4415),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4573),
.B(n_4376),
.Y(n_4615)
);

INVx2_ASAP7_75t_SL g4616 ( 
.A(n_4484),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4529),
.Y(n_4617)
);

OR2x2_ASAP7_75t_L g4618 ( 
.A(n_4590),
.B(n_4387),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4529),
.Y(n_4619)
);

OA21x2_ASAP7_75t_L g4620 ( 
.A1(n_4595),
.A2(n_4471),
.B(n_4552),
.Y(n_4620)
);

AO21x2_ASAP7_75t_L g4621 ( 
.A1(n_4584),
.A2(n_4420),
.B(n_4354),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4573),
.B(n_4424),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4573),
.B(n_4372),
.Y(n_4623)
);

NAND2x1p5_ASAP7_75t_L g4624 ( 
.A(n_4532),
.B(n_4418),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4526),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4532),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_4518),
.B(n_4362),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4498),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4505),
.Y(n_4629)
);

BUFx2_ASAP7_75t_L g4630 ( 
.A(n_4520),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4593),
.B(n_4390),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4516),
.Y(n_4632)
);

HB1xp67_ASAP7_75t_L g4633 ( 
.A(n_4567),
.Y(n_4633)
);

AOI22xp5_ASAP7_75t_SL g4634 ( 
.A1(n_4593),
.A2(n_4462),
.B1(n_4354),
.B2(n_4359),
.Y(n_4634)
);

AND2x2_ASAP7_75t_L g4635 ( 
.A(n_4518),
.B(n_4462),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4532),
.Y(n_4636)
);

AO21x2_ASAP7_75t_L g4637 ( 
.A1(n_4587),
.A2(n_4359),
.B(n_4426),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4518),
.B(n_4383),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4521),
.Y(n_4639)
);

OR2x2_ASAP7_75t_L g4640 ( 
.A(n_4601),
.B(n_4596),
.Y(n_4640)
);

HB1xp67_ASAP7_75t_L g4641 ( 
.A(n_4502),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4575),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4511),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4544),
.B(n_4416),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4497),
.B(n_4371),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4586),
.B(n_4589),
.Y(n_4646)
);

HB1xp67_ASAP7_75t_L g4647 ( 
.A(n_4528),
.Y(n_4647)
);

AND2x2_ASAP7_75t_L g4648 ( 
.A(n_4497),
.B(n_4411),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4514),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4575),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4575),
.Y(n_4651)
);

HB1xp67_ASAP7_75t_L g4652 ( 
.A(n_4589),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4473),
.B(n_4433),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4515),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4473),
.B(n_4454),
.Y(n_4655)
);

AND2x4_ASAP7_75t_L g4656 ( 
.A(n_4546),
.B(n_4548),
.Y(n_4656)
);

AND2x2_ASAP7_75t_L g4657 ( 
.A(n_4520),
.B(n_4461),
.Y(n_4657)
);

OR2x2_ASAP7_75t_L g4658 ( 
.A(n_4598),
.B(n_4384),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4523),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4533),
.Y(n_4660)
);

INVx2_ASAP7_75t_SL g4661 ( 
.A(n_4484),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4483),
.Y(n_4662)
);

HB1xp67_ASAP7_75t_L g4663 ( 
.A(n_4488),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4474),
.B(n_4384),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4513),
.B(n_4429),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4534),
.Y(n_4666)
);

NAND3xp33_ASAP7_75t_L g4667 ( 
.A(n_4599),
.B(n_4351),
.C(n_4402),
.Y(n_4667)
);

INVx2_ASAP7_75t_L g4668 ( 
.A(n_4575),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4479),
.Y(n_4669)
);

OAI21xp5_ASAP7_75t_SL g4670 ( 
.A1(n_4478),
.A2(n_4393),
.B(n_4399),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4481),
.Y(n_4671)
);

BUFx3_ASAP7_75t_L g4672 ( 
.A(n_4493),
.Y(n_4672)
);

INVx2_ASAP7_75t_L g4673 ( 
.A(n_4581),
.Y(n_4673)
);

AOI322xp5_ASAP7_75t_L g4674 ( 
.A1(n_4551),
.A2(n_4437),
.A3(n_4460),
.B1(n_623),
.B2(n_624),
.C1(n_625),
.C2(n_627),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4486),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4586),
.B(n_4460),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4556),
.B(n_685),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4546),
.B(n_685),
.Y(n_4678)
);

AO21x2_ASAP7_75t_L g4679 ( 
.A1(n_4560),
.A2(n_621),
.B(n_622),
.Y(n_4679)
);

NOR2xp33_ASAP7_75t_L g4680 ( 
.A(n_4478),
.B(n_622),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4581),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4483),
.Y(n_4682)
);

INVxp67_ASAP7_75t_SL g4683 ( 
.A(n_4592),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4536),
.B(n_623),
.Y(n_4684)
);

INVx5_ASAP7_75t_SL g4685 ( 
.A(n_4580),
.Y(n_4685)
);

OR2x2_ASAP7_75t_L g4686 ( 
.A(n_4490),
.B(n_625),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4495),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4536),
.B(n_629),
.Y(n_4688)
);

AND2x2_ASAP7_75t_L g4689 ( 
.A(n_4548),
.B(n_4485),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4581),
.Y(n_4690)
);

INVx4_ASAP7_75t_L g4691 ( 
.A(n_4509),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4506),
.Y(n_4692)
);

HB1xp67_ASAP7_75t_L g4693 ( 
.A(n_4488),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4469),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4485),
.B(n_4480),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4558),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4558),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4469),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4538),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4508),
.Y(n_4700)
);

NOR2x1_ASAP7_75t_SL g4701 ( 
.A(n_4482),
.B(n_632),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4494),
.Y(n_4702)
);

AOI22xp33_ASAP7_75t_L g4703 ( 
.A1(n_4545),
.A2(n_633),
.B1(n_634),
.B2(n_635),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4501),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4485),
.B(n_633),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4558),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4536),
.B(n_634),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4483),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4480),
.B(n_635),
.Y(n_4709)
);

AOI22xp33_ASAP7_75t_L g4710 ( 
.A1(n_4527),
.A2(n_637),
.B1(n_638),
.B2(n_639),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4483),
.Y(n_4711)
);

INVx2_ASAP7_75t_L g4712 ( 
.A(n_4580),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4580),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4496),
.B(n_638),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4483),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4527),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4527),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4657),
.B(n_4496),
.Y(n_4718)
);

HB1xp67_ASAP7_75t_L g4719 ( 
.A(n_4663),
.Y(n_4719)
);

BUFx2_ASAP7_75t_L g4720 ( 
.A(n_4672),
.Y(n_4720)
);

INVx4_ASAP7_75t_L g4721 ( 
.A(n_4672),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4693),
.Y(n_4722)
);

AND2x4_ASAP7_75t_L g4723 ( 
.A(n_4616),
.B(n_4661),
.Y(n_4723)
);

INVx3_ASAP7_75t_L g4724 ( 
.A(n_4715),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4662),
.Y(n_4725)
);

AND2x2_ASAP7_75t_L g4726 ( 
.A(n_4657),
.B(n_4503),
.Y(n_4726)
);

BUFx2_ASAP7_75t_L g4727 ( 
.A(n_4677),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4653),
.B(n_4630),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4630),
.B(n_4603),
.Y(n_4729)
);

INVx3_ASAP7_75t_L g4730 ( 
.A(n_4715),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4647),
.B(n_4603),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4662),
.Y(n_4732)
);

NAND2x1p5_ASAP7_75t_L g4733 ( 
.A(n_4677),
.B(n_4542),
.Y(n_4733)
);

OR2x2_ASAP7_75t_L g4734 ( 
.A(n_4640),
.B(n_4512),
.Y(n_4734)
);

BUFx2_ASAP7_75t_L g4735 ( 
.A(n_4616),
.Y(n_4735)
);

INVx1_ASAP7_75t_SL g4736 ( 
.A(n_4661),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4682),
.Y(n_4737)
);

INVx2_ASAP7_75t_L g4738 ( 
.A(n_4685),
.Y(n_4738)
);

BUFx2_ASAP7_75t_L g4739 ( 
.A(n_4683),
.Y(n_4739)
);

AND2x2_ASAP7_75t_L g4740 ( 
.A(n_4695),
.B(n_4509),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4640),
.B(n_4512),
.Y(n_4741)
);

INVx3_ASAP7_75t_L g4742 ( 
.A(n_4682),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4685),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_4685),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4653),
.B(n_4503),
.Y(n_4745)
);

OR2x2_ASAP7_75t_L g4746 ( 
.A(n_4658),
.B(n_4477),
.Y(n_4746)
);

INVxp67_ASAP7_75t_SL g4747 ( 
.A(n_4680),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4695),
.B(n_4500),
.Y(n_4748)
);

AND2x4_ASAP7_75t_L g4749 ( 
.A(n_4689),
.B(n_4500),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4708),
.Y(n_4750)
);

INVx3_ASAP7_75t_L g4751 ( 
.A(n_4624),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4689),
.B(n_4500),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_L g4753 ( 
.A(n_4634),
.B(n_4565),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4655),
.B(n_4560),
.Y(n_4754)
);

INVx4_ASAP7_75t_L g4755 ( 
.A(n_4691),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4701),
.B(n_4509),
.Y(n_4756)
);

HB1xp67_ASAP7_75t_L g4757 ( 
.A(n_4711),
.Y(n_4757)
);

OR2x2_ASAP7_75t_L g4758 ( 
.A(n_4658),
.B(n_4476),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4685),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4716),
.Y(n_4760)
);

AND2x4_ASAP7_75t_L g4761 ( 
.A(n_4656),
.B(n_4493),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4611),
.B(n_4476),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4701),
.B(n_4592),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_4635),
.B(n_4592),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4635),
.B(n_4597),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4614),
.B(n_4597),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4712),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4611),
.B(n_4476),
.Y(n_4768)
);

AND2x4_ASAP7_75t_L g4769 ( 
.A(n_4656),
.B(n_4475),
.Y(n_4769)
);

AND2x2_ASAP7_75t_L g4770 ( 
.A(n_4614),
.B(n_4597),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4716),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4712),
.Y(n_4772)
);

AND2x2_ASAP7_75t_L g4773 ( 
.A(n_4709),
.B(n_4488),
.Y(n_4773)
);

INVx2_ASAP7_75t_SL g4774 ( 
.A(n_4622),
.Y(n_4774)
);

AND2x2_ASAP7_75t_L g4775 ( 
.A(n_4655),
.B(n_4507),
.Y(n_4775)
);

BUFx3_ASAP7_75t_L g4776 ( 
.A(n_4705),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4713),
.Y(n_4777)
);

INVx2_ASAP7_75t_L g4778 ( 
.A(n_4717),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4713),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4717),
.Y(n_4780)
);

INVxp67_ASAP7_75t_L g4781 ( 
.A(n_4641),
.Y(n_4781)
);

INVx5_ASAP7_75t_L g4782 ( 
.A(n_4691),
.Y(n_4782)
);

INVx3_ASAP7_75t_L g4783 ( 
.A(n_4624),
.Y(n_4783)
);

INVxp33_ASAP7_75t_L g4784 ( 
.A(n_4613),
.Y(n_4784)
);

INVx3_ASAP7_75t_L g4785 ( 
.A(n_4624),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4727),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4731),
.B(n_4709),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4761),
.B(n_4691),
.Y(n_4788)
);

AND2x2_ASAP7_75t_L g4789 ( 
.A(n_4761),
.B(n_4633),
.Y(n_4789)
);

NAND3xp33_ASAP7_75t_L g4790 ( 
.A(n_4751),
.B(n_4620),
.C(n_4626),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4727),
.Y(n_4791)
);

HB1xp67_ASAP7_75t_L g4792 ( 
.A(n_4764),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_4761),
.B(n_4728),
.Y(n_4793)
);

OR2x2_ASAP7_75t_L g4794 ( 
.A(n_4753),
.B(n_4664),
.Y(n_4794)
);

INVxp67_ASAP7_75t_SL g4795 ( 
.A(n_4733),
.Y(n_4795)
);

INVx3_ASAP7_75t_L g4796 ( 
.A(n_4751),
.Y(n_4796)
);

OR2x2_ASAP7_75t_L g4797 ( 
.A(n_4753),
.B(n_4664),
.Y(n_4797)
);

AND2x2_ASAP7_75t_L g4798 ( 
.A(n_4761),
.B(n_4610),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4731),
.B(n_4627),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4751),
.Y(n_4800)
);

NOR2x1_ASAP7_75t_L g4801 ( 
.A(n_4721),
.B(n_4705),
.Y(n_4801)
);

NOR2xp33_ASAP7_75t_L g4802 ( 
.A(n_4751),
.B(n_4517),
.Y(n_4802)
);

INVxp67_ASAP7_75t_L g4803 ( 
.A(n_4720),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4783),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4739),
.Y(n_4805)
);

HB1xp67_ASAP7_75t_L g4806 ( 
.A(n_4764),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_SL g4807 ( 
.A(n_4783),
.B(n_4626),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4783),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4739),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4773),
.B(n_4627),
.Y(n_4810)
);

OR2x2_ASAP7_75t_L g4811 ( 
.A(n_4728),
.B(n_4625),
.Y(n_4811)
);

HB1xp67_ASAP7_75t_L g4812 ( 
.A(n_4720),
.Y(n_4812)
);

AND2x4_ASAP7_75t_L g4813 ( 
.A(n_4723),
.B(n_4656),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4757),
.Y(n_4814)
);

OR2x2_ASAP7_75t_L g4815 ( 
.A(n_4728),
.B(n_4646),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4773),
.B(n_4678),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4765),
.B(n_4610),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4729),
.B(n_4678),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4757),
.Y(n_4819)
);

BUFx3_ASAP7_75t_L g4820 ( 
.A(n_4735),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4729),
.B(n_4735),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4723),
.B(n_4714),
.Y(n_4822)
);

HB1xp67_ASAP7_75t_L g4823 ( 
.A(n_4765),
.Y(n_4823)
);

AND2x4_ASAP7_75t_SL g4824 ( 
.A(n_4723),
.B(n_4613),
.Y(n_4824)
);

BUFx2_ASAP7_75t_L g4825 ( 
.A(n_4723),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4742),
.Y(n_4826)
);

AND2x2_ASAP7_75t_L g4827 ( 
.A(n_4766),
.B(n_4622),
.Y(n_4827)
);

OR2x2_ASAP7_75t_L g4828 ( 
.A(n_4736),
.B(n_4774),
.Y(n_4828)
);

INVx2_ASAP7_75t_L g4829 ( 
.A(n_4783),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4742),
.Y(n_4830)
);

OAI21xp5_ASAP7_75t_SL g4831 ( 
.A1(n_4756),
.A2(n_4670),
.B(n_4667),
.Y(n_4831)
);

NAND3xp33_ASAP7_75t_L g4832 ( 
.A(n_4785),
.B(n_4620),
.C(n_4762),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4785),
.Y(n_4833)
);

NOR2xp33_ASAP7_75t_L g4834 ( 
.A(n_4785),
.B(n_4537),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4785),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4736),
.B(n_4714),
.Y(n_4836)
);

INVxp67_ASAP7_75t_SL g4837 ( 
.A(n_4733),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4766),
.B(n_4629),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4742),
.Y(n_4839)
);

BUFx2_ASAP7_75t_L g4840 ( 
.A(n_4776),
.Y(n_4840)
);

AOI22xp5_ASAP7_75t_L g4841 ( 
.A1(n_4754),
.A2(n_4620),
.B1(n_4621),
.B2(n_4637),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4733),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4790),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4813),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4793),
.B(n_4776),
.Y(n_4845)
);

AND2x4_ASAP7_75t_SL g4846 ( 
.A(n_4813),
.B(n_4756),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4792),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4793),
.B(n_4770),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4817),
.B(n_4776),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4813),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4817),
.B(n_4733),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4820),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4834),
.B(n_4774),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4806),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_4798),
.B(n_4770),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4834),
.B(n_4774),
.Y(n_4856)
);

AND2x2_ASAP7_75t_L g4857 ( 
.A(n_4798),
.B(n_4763),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4827),
.B(n_4763),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4820),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4841),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4827),
.B(n_4740),
.Y(n_4861)
);

BUFx3_ASAP7_75t_L g4862 ( 
.A(n_4840),
.Y(n_4862)
);

INVx1_ASAP7_75t_SL g4863 ( 
.A(n_4824),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4812),
.Y(n_4864)
);

AND2x2_ASAP7_75t_L g4865 ( 
.A(n_4824),
.B(n_4740),
.Y(n_4865)
);

OR2x2_ASAP7_75t_L g4866 ( 
.A(n_4794),
.B(n_4734),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4823),
.Y(n_4867)
);

AND2x4_ASAP7_75t_SL g4868 ( 
.A(n_4789),
.B(n_4721),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4825),
.B(n_4721),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4828),
.Y(n_4870)
);

AND2x2_ASAP7_75t_L g4871 ( 
.A(n_4789),
.B(n_4748),
.Y(n_4871)
);

AND2x2_ASAP7_75t_L g4872 ( 
.A(n_4838),
.B(n_4748),
.Y(n_4872)
);

OR2x2_ASAP7_75t_L g4873 ( 
.A(n_4794),
.B(n_4734),
.Y(n_4873)
);

OR2x2_ASAP7_75t_L g4874 ( 
.A(n_4797),
.B(n_4741),
.Y(n_4874)
);

HB1xp67_ASAP7_75t_L g4875 ( 
.A(n_4801),
.Y(n_4875)
);

AND2x4_ASAP7_75t_L g4876 ( 
.A(n_4795),
.B(n_4721),
.Y(n_4876)
);

NOR2x1_ASAP7_75t_L g4877 ( 
.A(n_4832),
.B(n_4755),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4837),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4838),
.B(n_4754),
.Y(n_4879)
);

INVxp67_ASAP7_75t_SL g4880 ( 
.A(n_4799),
.Y(n_4880)
);

INVx2_ASAP7_75t_L g4881 ( 
.A(n_4796),
.Y(n_4881)
);

OR2x2_ASAP7_75t_L g4882 ( 
.A(n_4797),
.B(n_4741),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4807),
.Y(n_4883)
);

BUFx3_ASAP7_75t_L g4884 ( 
.A(n_4788),
.Y(n_4884)
);

AND2x2_ASAP7_75t_L g4885 ( 
.A(n_4802),
.B(n_4748),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4807),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4803),
.B(n_4754),
.Y(n_4887)
);

HB1xp67_ASAP7_75t_L g4888 ( 
.A(n_4822),
.Y(n_4888)
);

AND2x2_ASAP7_75t_L g4889 ( 
.A(n_4802),
.B(n_4752),
.Y(n_4889)
);

OR2x2_ASAP7_75t_L g4890 ( 
.A(n_4815),
.B(n_4758),
.Y(n_4890)
);

BUFx3_ASAP7_75t_L g4891 ( 
.A(n_4788),
.Y(n_4891)
);

INVx2_ASAP7_75t_L g4892 ( 
.A(n_4796),
.Y(n_4892)
);

INVx2_ASAP7_75t_SL g4893 ( 
.A(n_4842),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4786),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4787),
.B(n_4747),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4861),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4861),
.B(n_4752),
.Y(n_4897)
);

OR2x2_ASAP7_75t_L g4898 ( 
.A(n_4879),
.B(n_4811),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4855),
.B(n_4752),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4855),
.B(n_4775),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4862),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4862),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4872),
.B(n_4848),
.Y(n_4903)
);

INVx3_ASAP7_75t_L g4904 ( 
.A(n_4883),
.Y(n_4904)
);

INVx2_ASAP7_75t_SL g4905 ( 
.A(n_4846),
.Y(n_4905)
);

AND2x4_ASAP7_75t_L g4906 ( 
.A(n_4865),
.B(n_4842),
.Y(n_4906)
);

INVx2_ASAP7_75t_SL g4907 ( 
.A(n_4846),
.Y(n_4907)
);

NOR2x1p5_ASAP7_75t_L g4908 ( 
.A(n_4849),
.B(n_4836),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4848),
.B(n_4745),
.Y(n_4909)
);

HB1xp67_ASAP7_75t_L g4910 ( 
.A(n_4883),
.Y(n_4910)
);

INVxp67_ASAP7_75t_SL g4911 ( 
.A(n_4886),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4872),
.Y(n_4912)
);

INVx2_ASAP7_75t_L g4913 ( 
.A(n_4886),
.Y(n_4913)
);

AOI32xp33_ASAP7_75t_L g4914 ( 
.A1(n_4843),
.A2(n_4775),
.A3(n_4784),
.B1(n_4718),
.B2(n_4726),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4866),
.Y(n_4915)
);

OR2x2_ASAP7_75t_L g4916 ( 
.A(n_4866),
.B(n_4821),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4873),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4873),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4871),
.B(n_4775),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4858),
.B(n_4745),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4874),
.Y(n_4921)
);

INVx3_ASAP7_75t_L g4922 ( 
.A(n_4884),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4874),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4882),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4858),
.B(n_4745),
.Y(n_4925)
);

OR2x2_ASAP7_75t_L g4926 ( 
.A(n_4882),
.B(n_4818),
.Y(n_4926)
);

AND2x4_ASAP7_75t_L g4927 ( 
.A(n_4865),
.B(n_4749),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4871),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4857),
.B(n_4749),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4887),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4857),
.B(n_4718),
.Y(n_4931)
);

AND2x2_ASAP7_75t_L g4932 ( 
.A(n_4885),
.B(n_4718),
.Y(n_4932)
);

AND2x2_ASAP7_75t_L g4933 ( 
.A(n_4885),
.B(n_4749),
.Y(n_4933)
);

AOI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4843),
.A2(n_4810),
.B1(n_4621),
.B2(n_4637),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4884),
.Y(n_4935)
);

OR2x2_ASAP7_75t_L g4936 ( 
.A(n_4909),
.B(n_4853),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4900),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4920),
.B(n_4856),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4903),
.Y(n_4939)
);

OAI21xp5_ASAP7_75t_L g4940 ( 
.A1(n_4934),
.A2(n_4831),
.B(n_4877),
.Y(n_4940)
);

OR2x2_ASAP7_75t_L g4941 ( 
.A(n_4925),
.B(n_4931),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4903),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4919),
.Y(n_4943)
);

NOR3xp33_ASAP7_75t_L g4944 ( 
.A(n_4915),
.B(n_4880),
.C(n_4895),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4932),
.B(n_4889),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_L g4946 ( 
.A(n_4911),
.B(n_4852),
.Y(n_4946)
);

OAI21xp5_ASAP7_75t_L g4947 ( 
.A1(n_4911),
.A2(n_4875),
.B(n_4860),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4897),
.B(n_4889),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4922),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4933),
.B(n_4863),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_4922),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4922),
.Y(n_4952)
);

OR2x2_ASAP7_75t_L g4953 ( 
.A(n_4916),
.B(n_4852),
.Y(n_4953)
);

NAND2x1p5_ASAP7_75t_L g4954 ( 
.A(n_4935),
.B(n_4859),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4910),
.B(n_4859),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_L g4956 ( 
.A(n_4910),
.B(n_4791),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4933),
.B(n_4929),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_4914),
.B(n_4800),
.Y(n_4958)
);

AND2x2_ASAP7_75t_L g4959 ( 
.A(n_4929),
.B(n_4891),
.Y(n_4959)
);

INVx4_ASAP7_75t_L g4960 ( 
.A(n_4935),
.Y(n_4960)
);

NAND2x1_ASAP7_75t_L g4961 ( 
.A(n_4927),
.B(n_4749),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4928),
.B(n_4800),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4928),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4896),
.B(n_4891),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4912),
.B(n_4726),
.Y(n_4965)
);

INVx2_ASAP7_75t_L g4966 ( 
.A(n_4927),
.Y(n_4966)
);

A2O1A1Ixp33_ASAP7_75t_L g4967 ( 
.A1(n_4913),
.A2(n_4758),
.B(n_4860),
.C(n_4768),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_4927),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4917),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_4959),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4948),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4945),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4965),
.Y(n_4973)
);

NAND2x1p5_ASAP7_75t_L g4974 ( 
.A(n_4953),
.B(n_4901),
.Y(n_4974)
);

INVx1_ASAP7_75t_SL g4975 ( 
.A(n_4957),
.Y(n_4975)
);

NOR2x1p5_ASAP7_75t_L g4976 ( 
.A(n_4961),
.B(n_4845),
.Y(n_4976)
);

OR2x6_ASAP7_75t_L g4977 ( 
.A(n_4966),
.B(n_4905),
.Y(n_4977)
);

OAI21xp33_ASAP7_75t_L g4978 ( 
.A1(n_4950),
.A2(n_4899),
.B(n_4726),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4954),
.Y(n_4979)
);

OR2x2_ASAP7_75t_L g4980 ( 
.A(n_4939),
.B(n_4918),
.Y(n_4980)
);

AND2x2_ASAP7_75t_L g4981 ( 
.A(n_4942),
.B(n_4921),
.Y(n_4981)
);

OR2x2_ASAP7_75t_L g4982 ( 
.A(n_4954),
.B(n_4923),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4964),
.B(n_4905),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4946),
.Y(n_4984)
);

NOR2xp33_ASAP7_75t_L g4985 ( 
.A(n_4960),
.B(n_4816),
.Y(n_4985)
);

INVx1_ASAP7_75t_SL g4986 ( 
.A(n_4941),
.Y(n_4986)
);

OR2x6_ASAP7_75t_L g4987 ( 
.A(n_4968),
.B(n_4907),
.Y(n_4987)
);

NAND2x1p5_ASAP7_75t_L g4988 ( 
.A(n_4960),
.B(n_4902),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4937),
.B(n_4924),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4946),
.Y(n_4990)
);

AND2x2_ASAP7_75t_L g4991 ( 
.A(n_4943),
.B(n_4907),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4955),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4951),
.B(n_4868),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4955),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4947),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4963),
.B(n_4868),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4944),
.B(n_4908),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4982),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4974),
.Y(n_4999)
);

NOR3xp33_ASAP7_75t_L g5000 ( 
.A(n_4995),
.B(n_4947),
.C(n_4940),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4975),
.B(n_4870),
.Y(n_5001)
);

AOI32xp33_ASAP7_75t_L g5002 ( 
.A1(n_4995),
.A2(n_4904),
.A3(n_4913),
.B1(n_4997),
.B2(n_4796),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4976),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4986),
.B(n_4906),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4988),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4979),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4971),
.B(n_4888),
.Y(n_5007)
);

INVx2_ASAP7_75t_L g5008 ( 
.A(n_4977),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4978),
.B(n_4904),
.Y(n_5009)
);

INVx2_ASAP7_75t_L g5010 ( 
.A(n_4977),
.Y(n_5010)
);

INVxp67_ASAP7_75t_L g5011 ( 
.A(n_4985),
.Y(n_5011)
);

OAI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4992),
.A2(n_4940),
.B(n_4967),
.Y(n_5012)
);

NOR2xp67_ASAP7_75t_SL g5013 ( 
.A(n_4970),
.B(n_4949),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4979),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4987),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4972),
.B(n_4906),
.Y(n_5016)
);

NOR2xp33_ASAP7_75t_L g5017 ( 
.A(n_4994),
.B(n_4851),
.Y(n_5017)
);

NAND2x1p5_ASAP7_75t_L g5018 ( 
.A(n_4991),
.B(n_4952),
.Y(n_5018)
);

OR2x2_ASAP7_75t_L g5019 ( 
.A(n_4987),
.B(n_4926),
.Y(n_5019)
);

AO21x1_ASAP7_75t_L g5020 ( 
.A1(n_5000),
.A2(n_4956),
.B(n_4962),
.Y(n_5020)
);

AOI21xp33_ASAP7_75t_SL g5021 ( 
.A1(n_5019),
.A2(n_4956),
.B(n_4962),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_L g5022 ( 
.A(n_5001),
.B(n_4906),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_5004),
.Y(n_5023)
);

INVx2_ASAP7_75t_L g5024 ( 
.A(n_5018),
.Y(n_5024)
);

OAI22xp5_ASAP7_75t_L g5025 ( 
.A1(n_5016),
.A2(n_4980),
.B1(n_4890),
.B2(n_4969),
.Y(n_5025)
);

AND2x2_ASAP7_75t_L g5026 ( 
.A(n_5007),
.B(n_4981),
.Y(n_5026)
);

AOI22xp5_ASAP7_75t_L g5027 ( 
.A1(n_5015),
.A2(n_4747),
.B1(n_4893),
.B2(n_4808),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_5008),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_5012),
.Y(n_5029)
);

OAI22xp5_ASAP7_75t_L g5030 ( 
.A1(n_4998),
.A2(n_4890),
.B1(n_4973),
.B2(n_4958),
.Y(n_5030)
);

OR2x2_ASAP7_75t_L g5031 ( 
.A(n_5010),
.B(n_4898),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_5013),
.Y(n_5032)
);

OR2x2_ASAP7_75t_L g5033 ( 
.A(n_4999),
.B(n_4844),
.Y(n_5033)
);

OR2x2_ASAP7_75t_L g5034 ( 
.A(n_5009),
.B(n_4844),
.Y(n_5034)
);

INVxp67_ASAP7_75t_SL g5035 ( 
.A(n_5009),
.Y(n_5035)
);

AOI21xp33_ASAP7_75t_L g5036 ( 
.A1(n_5012),
.A2(n_4743),
.B(n_4738),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_5003),
.B(n_4989),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_5029),
.B(n_4850),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_5026),
.B(n_4973),
.Y(n_5039)
);

NOR2x1_ASAP7_75t_L g5040 ( 
.A(n_5022),
.B(n_4983),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_5037),
.B(n_4850),
.Y(n_5041)
);

AOI22xp5_ASAP7_75t_L g5042 ( 
.A1(n_5032),
.A2(n_5017),
.B1(n_4893),
.B2(n_4804),
.Y(n_5042)
);

INVx2_ASAP7_75t_SL g5043 ( 
.A(n_5031),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_5020),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_5024),
.B(n_4867),
.Y(n_5045)
);

OAI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_5029),
.A2(n_4958),
.B(n_4992),
.Y(n_5046)
);

OAI21xp5_ASAP7_75t_SL g5047 ( 
.A1(n_5027),
.A2(n_5002),
.B(n_5011),
.Y(n_5047)
);

A2O1A1Ixp33_ASAP7_75t_L g5048 ( 
.A1(n_5036),
.A2(n_5002),
.B(n_4990),
.C(n_4984),
.Y(n_5048)
);

OAI221xp5_ASAP7_75t_L g5049 ( 
.A1(n_5035),
.A2(n_4835),
.B1(n_4833),
.B2(n_4829),
.C(n_4808),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_5021),
.B(n_4804),
.Y(n_5050)
);

AOI21xp5_ASAP7_75t_L g5051 ( 
.A1(n_5030),
.A2(n_4869),
.B(n_4996),
.Y(n_5051)
);

AOI32xp33_ASAP7_75t_L g5052 ( 
.A1(n_5025),
.A2(n_4904),
.A3(n_4878),
.B1(n_4990),
.B2(n_4984),
.Y(n_5052)
);

AOI221xp5_ASAP7_75t_SL g5053 ( 
.A1(n_5023),
.A2(n_4805),
.B1(n_4809),
.B2(n_4864),
.C(n_4781),
.Y(n_5053)
);

AND2x2_ASAP7_75t_L g5054 ( 
.A(n_5033),
.B(n_4847),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_5034),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_5028),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_5026),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_5026),
.Y(n_5058)
);

OAI211xp5_ASAP7_75t_L g5059 ( 
.A1(n_5052),
.A2(n_4993),
.B(n_5005),
.C(n_5006),
.Y(n_5059)
);

INVx2_ASAP7_75t_SL g5060 ( 
.A(n_5041),
.Y(n_5060)
);

AOI22xp5_ASAP7_75t_L g5061 ( 
.A1(n_5055),
.A2(n_4833),
.B1(n_4835),
.B2(n_4829),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5043),
.B(n_4876),
.Y(n_5062)
);

AOI322xp5_ASAP7_75t_L g5063 ( 
.A1(n_5044),
.A2(n_4768),
.A3(n_4762),
.B1(n_4743),
.B2(n_4744),
.C1(n_4759),
.C2(n_4738),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_5039),
.Y(n_5064)
);

AND2x2_ASAP7_75t_L g5065 ( 
.A(n_5040),
.B(n_4854),
.Y(n_5065)
);

O2A1O1Ixp33_ASAP7_75t_L g5066 ( 
.A1(n_5044),
.A2(n_5014),
.B(n_4892),
.C(n_4881),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_5054),
.B(n_4781),
.Y(n_5067)
);

O2A1O1Ixp5_ASAP7_75t_L g5068 ( 
.A1(n_5046),
.A2(n_4892),
.B(n_4881),
.C(n_4876),
.Y(n_5068)
);

INVx1_ASAP7_75t_SL g5069 ( 
.A(n_5038),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_5057),
.Y(n_5070)
);

NOR3xp33_ASAP7_75t_L g5071 ( 
.A(n_5047),
.B(n_4930),
.C(n_4936),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_5058),
.Y(n_5072)
);

OAI21xp33_ASAP7_75t_L g5073 ( 
.A1(n_5045),
.A2(n_4938),
.B(n_4894),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_5056),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_5042),
.B(n_4876),
.Y(n_5075)
);

AOI22xp5_ASAP7_75t_L g5076 ( 
.A1(n_5050),
.A2(n_4738),
.B1(n_4744),
.B2(n_4743),
.Y(n_5076)
);

INVx3_ASAP7_75t_L g5077 ( 
.A(n_5053),
.Y(n_5077)
);

OAI22xp33_ASAP7_75t_L g5078 ( 
.A1(n_5049),
.A2(n_4759),
.B1(n_4744),
.B2(n_4636),
.Y(n_5078)
);

AOI32xp33_ASAP7_75t_L g5079 ( 
.A1(n_5048),
.A2(n_4814),
.A3(n_4819),
.B1(n_4722),
.B2(n_4826),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_L g5080 ( 
.A1(n_5051),
.A2(n_4759),
.B1(n_4771),
.B2(n_4760),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_5043),
.B(n_4746),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_5041),
.Y(n_5082)
);

OR2x2_ASAP7_75t_L g5083 ( 
.A(n_5038),
.B(n_4746),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5041),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_5043),
.B(n_4769),
.Y(n_5085)
);

OAI322xp33_ASAP7_75t_L g5086 ( 
.A1(n_5044),
.A2(n_4722),
.A3(n_4839),
.B1(n_4830),
.B2(n_4719),
.C1(n_4779),
.C2(n_4767),
.Y(n_5086)
);

AOI211xp5_ASAP7_75t_L g5087 ( 
.A1(n_5078),
.A2(n_4719),
.B(n_4772),
.C(n_4767),
.Y(n_5087)
);

AOI22xp5_ASAP7_75t_L g5088 ( 
.A1(n_5060),
.A2(n_4780),
.B1(n_4760),
.B2(n_4778),
.Y(n_5088)
);

AOI221xp5_ASAP7_75t_L g5089 ( 
.A1(n_5066),
.A2(n_4777),
.B1(n_4772),
.B2(n_4779),
.C(n_4778),
.Y(n_5089)
);

AOI21xp5_ASAP7_75t_L g5090 ( 
.A1(n_5081),
.A2(n_4771),
.B(n_4760),
.Y(n_5090)
);

AOI22xp33_ASAP7_75t_L g5091 ( 
.A1(n_5069),
.A2(n_4771),
.B1(n_4780),
.B2(n_4778),
.Y(n_5091)
);

AOI221xp5_ASAP7_75t_L g5092 ( 
.A1(n_5080),
.A2(n_4777),
.B1(n_4780),
.B2(n_4742),
.C(n_4750),
.Y(n_5092)
);

OAI22xp5_ASAP7_75t_L g5093 ( 
.A1(n_5064),
.A2(n_4607),
.B1(n_4769),
.B2(n_4702),
.Y(n_5093)
);

AOI211xp5_ASAP7_75t_L g5094 ( 
.A1(n_5065),
.A2(n_4769),
.B(n_4700),
.C(n_4704),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_5083),
.Y(n_5095)
);

INVxp67_ASAP7_75t_L g5096 ( 
.A(n_5085),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5062),
.Y(n_5097)
);

NOR2xp33_ASAP7_75t_L g5098 ( 
.A(n_5082),
.B(n_4569),
.Y(n_5098)
);

NAND2x1_ASAP7_75t_L g5099 ( 
.A(n_5067),
.B(n_4755),
.Y(n_5099)
);

INVxp67_ASAP7_75t_L g5100 ( 
.A(n_5075),
.Y(n_5100)
);

NOR2xp33_ASAP7_75t_L g5101 ( 
.A(n_5084),
.B(n_4755),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5068),
.Y(n_5102)
);

OAI211xp5_ASAP7_75t_L g5103 ( 
.A1(n_5073),
.A2(n_4755),
.B(n_4782),
.C(n_4632),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5061),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5070),
.Y(n_5105)
);

XNOR2xp5_ASAP7_75t_L g5106 ( 
.A(n_5072),
.B(n_4537),
.Y(n_5106)
);

OAI22xp33_ASAP7_75t_L g5107 ( 
.A1(n_5076),
.A2(n_4636),
.B1(n_4782),
.B2(n_4750),
.Y(n_5107)
);

AOI221xp5_ASAP7_75t_L g5108 ( 
.A1(n_5074),
.A2(n_4737),
.B1(n_4732),
.B2(n_4725),
.C(n_4769),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_5071),
.Y(n_5109)
);

AND2x2_ASAP7_75t_L g5110 ( 
.A(n_5077),
.B(n_4652),
.Y(n_5110)
);

OAI22xp5_ASAP7_75t_L g5111 ( 
.A1(n_5077),
.A2(n_4782),
.B1(n_4699),
.B2(n_4628),
.Y(n_5111)
);

AOI221xp5_ASAP7_75t_L g5112 ( 
.A1(n_5086),
.A2(n_4737),
.B1(n_4732),
.B2(n_4725),
.C(n_4730),
.Y(n_5112)
);

O2A1O1Ixp33_ASAP7_75t_L g5113 ( 
.A1(n_5059),
.A2(n_4576),
.B(n_4681),
.C(n_4690),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_5063),
.Y(n_5114)
);

OAI221xp5_ASAP7_75t_L g5115 ( 
.A1(n_5079),
.A2(n_4782),
.B1(n_4730),
.B2(n_4724),
.C(n_4639),
.Y(n_5115)
);

OR2x2_ASAP7_75t_L g5116 ( 
.A(n_5083),
.B(n_4694),
.Y(n_5116)
);

NOR3xp33_ASAP7_75t_L g5117 ( 
.A(n_5062),
.B(n_4681),
.C(n_4673),
.Y(n_5117)
);

AOI22xp33_ASAP7_75t_L g5118 ( 
.A1(n_5069),
.A2(n_4730),
.B1(n_4724),
.B2(n_4690),
.Y(n_5118)
);

OAI221xp5_ASAP7_75t_L g5119 ( 
.A1(n_5081),
.A2(n_4782),
.B1(n_4730),
.B2(n_4724),
.C(n_4686),
.Y(n_5119)
);

XOR2x2_ASAP7_75t_L g5120 ( 
.A(n_5081),
.B(n_4612),
.Y(n_5120)
);

INVxp67_ASAP7_75t_SL g5121 ( 
.A(n_5100),
.Y(n_5121)
);

AOI221xp5_ASAP7_75t_L g5122 ( 
.A1(n_5113),
.A2(n_4724),
.B1(n_4782),
.B2(n_4617),
.C(n_4619),
.Y(n_5122)
);

AOI221xp5_ASAP7_75t_L g5123 ( 
.A1(n_5117),
.A2(n_4782),
.B1(n_4608),
.B2(n_4609),
.C(n_4698),
.Y(n_5123)
);

NOR2xp33_ASAP7_75t_L g5124 ( 
.A(n_5106),
.B(n_4642),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_SL g5125 ( 
.A(n_5102),
.B(n_4686),
.Y(n_5125)
);

NOR2x1_ASAP7_75t_L g5126 ( 
.A(n_5105),
.B(n_4669),
.Y(n_5126)
);

AOI21xp5_ASAP7_75t_L g5127 ( 
.A1(n_5110),
.A2(n_4676),
.B(n_4621),
.Y(n_5127)
);

AOI322xp5_ASAP7_75t_L g5128 ( 
.A1(n_5114),
.A2(n_4673),
.A3(n_4697),
.B1(n_4706),
.B2(n_4696),
.C1(n_4684),
.C2(n_4707),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_L g5129 ( 
.A(n_5118),
.B(n_4679),
.Y(n_5129)
);

AOI21xp5_ASAP7_75t_L g5130 ( 
.A1(n_5109),
.A2(n_4631),
.B(n_4642),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_L g5131 ( 
.A(n_5120),
.B(n_4679),
.Y(n_5131)
);

AOI211xp5_ASAP7_75t_L g5132 ( 
.A1(n_5111),
.A2(n_4554),
.B(n_4638),
.C(n_4692),
.Y(n_5132)
);

OAI21xp33_ASAP7_75t_SL g5133 ( 
.A1(n_5101),
.A2(n_4675),
.B(n_4671),
.Y(n_5133)
);

NAND2xp5_ASAP7_75t_L g5134 ( 
.A(n_5091),
.B(n_4679),
.Y(n_5134)
);

AOI221xp5_ASAP7_75t_L g5135 ( 
.A1(n_5107),
.A2(n_4706),
.B1(n_4697),
.B2(n_4696),
.C(n_4568),
.Y(n_5135)
);

OAI21xp5_ASAP7_75t_L g5136 ( 
.A1(n_5096),
.A2(n_4648),
.B(n_4618),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_SL g5137 ( 
.A(n_5095),
.B(n_4579),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_5088),
.Y(n_5138)
);

OAI31xp33_ASAP7_75t_L g5139 ( 
.A1(n_5104),
.A2(n_4638),
.A3(n_4618),
.B(n_4568),
.Y(n_5139)
);

AOI211xp5_ASAP7_75t_L g5140 ( 
.A1(n_5097),
.A2(n_4687),
.B(n_4542),
.C(n_4543),
.Y(n_5140)
);

NAND3xp33_ASAP7_75t_L g5141 ( 
.A(n_5098),
.B(n_4651),
.C(n_4650),
.Y(n_5141)
);

NAND4xp25_ASAP7_75t_L g5142 ( 
.A(n_5090),
.B(n_4668),
.C(n_4650),
.D(n_4651),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_L g5143 ( 
.A(n_5094),
.B(n_4668),
.Y(n_5143)
);

AOI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_5092),
.A2(n_4637),
.B1(n_4648),
.B2(n_4645),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_5087),
.B(n_4665),
.Y(n_5145)
);

OAI21xp33_ASAP7_75t_SL g5146 ( 
.A1(n_5112),
.A2(n_4649),
.B(n_4643),
.Y(n_5146)
);

NAND4xp25_ASAP7_75t_L g5147 ( 
.A(n_5089),
.B(n_4543),
.C(n_4623),
.D(n_4688),
.Y(n_5147)
);

AOI211xp5_ASAP7_75t_L g5148 ( 
.A1(n_5115),
.A2(n_4660),
.B(n_4654),
.C(n_4666),
.Y(n_5148)
);

OAI22xp5_ASAP7_75t_L g5149 ( 
.A1(n_5119),
.A2(n_4659),
.B1(n_4568),
.B2(n_4547),
.Y(n_5149)
);

NOR3x1_ASAP7_75t_L g5150 ( 
.A(n_5121),
.B(n_5099),
.C(n_5103),
.Y(n_5150)
);

AO21x1_ASAP7_75t_L g5151 ( 
.A1(n_5137),
.A2(n_5093),
.B(n_5116),
.Y(n_5151)
);

OAI21xp33_ASAP7_75t_SL g5152 ( 
.A1(n_5126),
.A2(n_5108),
.B(n_4507),
.Y(n_5152)
);

AND3x4_ASAP7_75t_L g5153 ( 
.A(n_5125),
.B(n_4487),
.C(n_4489),
.Y(n_5153)
);

NAND3xp33_ASAP7_75t_L g5154 ( 
.A(n_5138),
.B(n_5124),
.C(n_5130),
.Y(n_5154)
);

AOI21xp5_ASAP7_75t_SL g5155 ( 
.A1(n_5145),
.A2(n_4489),
.B(n_4475),
.Y(n_5155)
);

AND2x2_ASAP7_75t_SL g5156 ( 
.A(n_5143),
.B(n_5131),
.Y(n_5156)
);

OAI211xp5_ASAP7_75t_L g5157 ( 
.A1(n_5122),
.A2(n_4547),
.B(n_4623),
.C(n_4487),
.Y(n_5157)
);

NOR2xp33_ASAP7_75t_L g5158 ( 
.A(n_5142),
.B(n_4579),
.Y(n_5158)
);

INVx2_ASAP7_75t_L g5159 ( 
.A(n_5134),
.Y(n_5159)
);

AOI221xp5_ASAP7_75t_L g5160 ( 
.A1(n_5129),
.A2(n_4547),
.B1(n_4645),
.B2(n_4665),
.C(n_4579),
.Y(n_5160)
);

AOI21xp33_ASAP7_75t_L g5161 ( 
.A1(n_5141),
.A2(n_4612),
.B(n_4561),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_5136),
.Y(n_5162)
);

NOR4xp25_ASAP7_75t_L g5163 ( 
.A(n_5146),
.B(n_4615),
.C(n_4571),
.D(n_4564),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_5127),
.B(n_4579),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_5144),
.B(n_4579),
.Y(n_5165)
);

AOI321xp33_ASAP7_75t_L g5166 ( 
.A1(n_5123),
.A2(n_5132),
.A3(n_5135),
.B1(n_5148),
.B2(n_5149),
.C(n_5140),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_SL g5167 ( 
.A(n_5139),
.B(n_4615),
.Y(n_5167)
);

AOI21xp33_ASAP7_75t_SL g5168 ( 
.A1(n_5133),
.A2(n_4561),
.B(n_4588),
.Y(n_5168)
);

OAI22xp5_ASAP7_75t_L g5169 ( 
.A1(n_5147),
.A2(n_4519),
.B1(n_4588),
.B2(n_4602),
.Y(n_5169)
);

OAI322xp33_ASAP7_75t_L g5170 ( 
.A1(n_5167),
.A2(n_5128),
.A3(n_4644),
.B1(n_4585),
.B2(n_4519),
.C1(n_4557),
.C2(n_4582),
.Y(n_5170)
);

OAI221xp5_ASAP7_75t_L g5171 ( 
.A1(n_5163),
.A2(n_4482),
.B1(n_4492),
.B2(n_4703),
.C(n_4710),
.Y(n_5171)
);

NOR3xp33_ASAP7_75t_L g5172 ( 
.A(n_5154),
.B(n_5162),
.C(n_5159),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_5164),
.Y(n_5173)
);

OAI211xp5_ASAP7_75t_L g5174 ( 
.A1(n_5166),
.A2(n_4674),
.B(n_4472),
.C(n_4553),
.Y(n_5174)
);

AOI21xp5_ASAP7_75t_L g5175 ( 
.A1(n_5165),
.A2(n_4555),
.B(n_4553),
.Y(n_5175)
);

AND3x2_ASAP7_75t_L g5176 ( 
.A(n_5158),
.B(n_4555),
.C(n_4594),
.Y(n_5176)
);

AND2x2_ASAP7_75t_L g5177 ( 
.A(n_5160),
.B(n_4504),
.Y(n_5177)
);

NOR3xp33_ASAP7_75t_L g5178 ( 
.A(n_5152),
.B(n_4472),
.C(n_4578),
.Y(n_5178)
);

AOI22x1_ASAP7_75t_SL g5179 ( 
.A1(n_5150),
.A2(n_4594),
.B1(n_4574),
.B2(n_4524),
.Y(n_5179)
);

NOR2xp67_ASAP7_75t_L g5180 ( 
.A(n_5157),
.B(n_639),
.Y(n_5180)
);

AND2x2_ASAP7_75t_L g5181 ( 
.A(n_5168),
.B(n_4504),
.Y(n_5181)
);

NOR4xp25_ASAP7_75t_SL g5182 ( 
.A(n_5151),
.B(n_4562),
.C(n_4491),
.D(n_4550),
.Y(n_5182)
);

NAND3xp33_ASAP7_75t_SL g5183 ( 
.A(n_5153),
.B(n_4540),
.C(n_4524),
.Y(n_5183)
);

OAI21xp5_ASAP7_75t_SL g5184 ( 
.A1(n_5161),
.A2(n_4540),
.B(n_4531),
.Y(n_5184)
);

NOR2xp33_ASAP7_75t_L g5185 ( 
.A(n_5155),
.B(n_4522),
.Y(n_5185)
);

NAND3xp33_ASAP7_75t_SL g5186 ( 
.A(n_5156),
.B(n_4522),
.C(n_4600),
.Y(n_5186)
);

NOR2xp33_ASAP7_75t_L g5187 ( 
.A(n_5169),
.B(n_4539),
.Y(n_5187)
);

NOR2x1_ASAP7_75t_L g5188 ( 
.A(n_5173),
.B(n_4550),
.Y(n_5188)
);

NOR2xp33_ASAP7_75t_L g5189 ( 
.A(n_5181),
.B(n_4539),
.Y(n_5189)
);

AOI22xp5_ASAP7_75t_L g5190 ( 
.A1(n_5172),
.A2(n_4504),
.B1(n_4510),
.B2(n_4550),
.Y(n_5190)
);

NOR3xp33_ASAP7_75t_L g5191 ( 
.A(n_5180),
.B(n_4531),
.C(n_4541),
.Y(n_5191)
);

OAI211xp5_ASAP7_75t_SL g5192 ( 
.A1(n_5185),
.A2(n_640),
.B(n_641),
.C(n_642),
.Y(n_5192)
);

AOI21xp5_ASAP7_75t_L g5193 ( 
.A1(n_5177),
.A2(n_4482),
.B(n_4510),
.Y(n_5193)
);

NOR3xp33_ASAP7_75t_L g5194 ( 
.A(n_5186),
.B(n_4531),
.C(n_4541),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_5178),
.B(n_4541),
.Y(n_5195)
);

NOR2x1_ASAP7_75t_L g5196 ( 
.A(n_5183),
.B(n_4482),
.Y(n_5196)
);

AND2x2_ASAP7_75t_L g5197 ( 
.A(n_5184),
.B(n_4530),
.Y(n_5197)
);

NOR4xp75_ASAP7_75t_L g5198 ( 
.A(n_5170),
.B(n_4605),
.C(n_642),
.D(n_643),
.Y(n_5198)
);

INVx1_ASAP7_75t_SL g5199 ( 
.A(n_5187),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_5175),
.B(n_4510),
.Y(n_5200)
);

NOR2x1_ASAP7_75t_L g5201 ( 
.A(n_5174),
.B(n_4499),
.Y(n_5201)
);

NOR3x1_ASAP7_75t_L g5202 ( 
.A(n_5171),
.B(n_4605),
.C(n_643),
.Y(n_5202)
);

OAI211xp5_ASAP7_75t_SL g5203 ( 
.A1(n_5179),
.A2(n_641),
.B(n_644),
.C(n_645),
.Y(n_5203)
);

NOR2x1_ASAP7_75t_L g5204 ( 
.A(n_5176),
.B(n_4499),
.Y(n_5204)
);

NOR3xp33_ASAP7_75t_L g5205 ( 
.A(n_5182),
.B(n_4572),
.C(n_4570),
.Y(n_5205)
);

AND2x4_ASAP7_75t_L g5206 ( 
.A(n_5172),
.B(n_4559),
.Y(n_5206)
);

NOR2x1_ASAP7_75t_L g5207 ( 
.A(n_5203),
.B(n_4499),
.Y(n_5207)
);

A2O1A1Ixp33_ASAP7_75t_L g5208 ( 
.A1(n_5196),
.A2(n_4572),
.B(n_4570),
.C(n_4563),
.Y(n_5208)
);

INVxp67_ASAP7_75t_L g5209 ( 
.A(n_5206),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_5200),
.Y(n_5210)
);

O2A1O1Ixp33_ASAP7_75t_L g5211 ( 
.A1(n_5199),
.A2(n_4562),
.B(n_4492),
.C(n_4559),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5195),
.Y(n_5212)
);

OA22x2_ASAP7_75t_L g5213 ( 
.A1(n_5197),
.A2(n_4492),
.B1(n_4563),
.B2(n_4530),
.Y(n_5213)
);

AO22x2_ASAP7_75t_L g5214 ( 
.A1(n_5205),
.A2(n_4562),
.B1(n_4492),
.B2(n_647),
.Y(n_5214)
);

NOR2x1_ASAP7_75t_L g5215 ( 
.A(n_5192),
.B(n_4566),
.Y(n_5215)
);

AND2x2_ASAP7_75t_L g5216 ( 
.A(n_5191),
.B(n_4583),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_5189),
.B(n_4606),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_5202),
.Y(n_5218)
);

AO22x2_ASAP7_75t_L g5219 ( 
.A1(n_5193),
.A2(n_645),
.B1(n_646),
.B2(n_647),
.Y(n_5219)
);

INVxp67_ASAP7_75t_L g5220 ( 
.A(n_5201),
.Y(n_5220)
);

AO22x2_ASAP7_75t_L g5221 ( 
.A1(n_5194),
.A2(n_646),
.B1(n_648),
.B2(n_649),
.Y(n_5221)
);

NOR2xp67_ASAP7_75t_L g5222 ( 
.A(n_5190),
.B(n_648),
.Y(n_5222)
);

AOI22xp5_ASAP7_75t_L g5223 ( 
.A1(n_5204),
.A2(n_4566),
.B1(n_4583),
.B2(n_4606),
.Y(n_5223)
);

NOR2x1_ASAP7_75t_L g5224 ( 
.A(n_5188),
.B(n_4566),
.Y(n_5224)
);

OR2x2_ASAP7_75t_L g5225 ( 
.A(n_5217),
.B(n_5198),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_5219),
.Y(n_5226)
);

NAND4xp25_ASAP7_75t_L g5227 ( 
.A(n_5218),
.B(n_4604),
.C(n_650),
.D(n_651),
.Y(n_5227)
);

NAND5xp2_ASAP7_75t_L g5228 ( 
.A(n_5210),
.B(n_649),
.C(n_650),
.D(n_652),
.E(n_653),
.Y(n_5228)
);

NAND3xp33_ASAP7_75t_L g5229 ( 
.A(n_5220),
.B(n_4591),
.C(n_654),
.Y(n_5229)
);

NAND4xp75_ASAP7_75t_L g5230 ( 
.A(n_5212),
.B(n_4591),
.C(n_654),
.D(n_655),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5209),
.B(n_4606),
.Y(n_5231)
);

OR2x2_ASAP7_75t_L g5232 ( 
.A(n_5216),
.B(n_4583),
.Y(n_5232)
);

INVx2_ASAP7_75t_L g5233 ( 
.A(n_5221),
.Y(n_5233)
);

NAND3xp33_ASAP7_75t_L g5234 ( 
.A(n_5222),
.B(n_4591),
.C(n_656),
.Y(n_5234)
);

NOR3xp33_ASAP7_75t_L g5235 ( 
.A(n_5215),
.B(n_653),
.C(n_656),
.Y(n_5235)
);

NAND4xp75_ASAP7_75t_L g5236 ( 
.A(n_5207),
.B(n_657),
.C(n_658),
.D(n_659),
.Y(n_5236)
);

NOR2xp33_ASAP7_75t_L g5237 ( 
.A(n_5226),
.B(n_5208),
.Y(n_5237)
);

AND2x2_ASAP7_75t_L g5238 ( 
.A(n_5233),
.B(n_5213),
.Y(n_5238)
);

NOR2x1_ASAP7_75t_L g5239 ( 
.A(n_5236),
.B(n_5224),
.Y(n_5239)
);

NOR2x1_ASAP7_75t_L g5240 ( 
.A(n_5225),
.B(n_5211),
.Y(n_5240)
);

INVx2_ASAP7_75t_SL g5241 ( 
.A(n_5234),
.Y(n_5241)
);

AND2x4_ASAP7_75t_L g5242 ( 
.A(n_5235),
.B(n_5223),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5228),
.Y(n_5243)
);

AND2x4_ASAP7_75t_L g5244 ( 
.A(n_5238),
.B(n_5229),
.Y(n_5244)
);

XNOR2x1_ASAP7_75t_SL g5245 ( 
.A(n_5241),
.B(n_5214),
.Y(n_5245)
);

AND2x4_ASAP7_75t_L g5246 ( 
.A(n_5243),
.B(n_5232),
.Y(n_5246)
);

BUFx2_ASAP7_75t_L g5247 ( 
.A(n_5240),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5247),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5245),
.Y(n_5249)
);

AO22x2_ASAP7_75t_L g5250 ( 
.A1(n_5248),
.A2(n_5246),
.B1(n_5244),
.B2(n_5242),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_5250),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5251),
.Y(n_5252)
);

AOI21xp5_ASAP7_75t_L g5253 ( 
.A1(n_5252),
.A2(n_5249),
.B(n_5237),
.Y(n_5253)
);

OAI22xp5_ASAP7_75t_L g5254 ( 
.A1(n_5253),
.A2(n_5239),
.B1(n_5230),
.B2(n_5231),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5254),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_5255),
.Y(n_5256)
);

AOI22xp5_ASAP7_75t_L g5257 ( 
.A1(n_5256),
.A2(n_5227),
.B1(n_662),
.B2(n_663),
.Y(n_5257)
);

AOI22x1_ASAP7_75t_L g5258 ( 
.A1(n_5257),
.A2(n_661),
.B1(n_662),
.B2(n_664),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_5258),
.Y(n_5259)
);

OA21x2_ASAP7_75t_L g5260 ( 
.A1(n_5259),
.A2(n_661),
.B(n_664),
.Y(n_5260)
);

AOI22xp33_ASAP7_75t_L g5261 ( 
.A1(n_5260),
.A2(n_668),
.B1(n_669),
.B2(n_670),
.Y(n_5261)
);

AOI22xp5_ASAP7_75t_L g5262 ( 
.A1(n_5261),
.A2(n_673),
.B1(n_674),
.B2(n_675),
.Y(n_5262)
);

AOI211xp5_ASAP7_75t_L g5263 ( 
.A1(n_5262),
.A2(n_673),
.B(n_674),
.C(n_675),
.Y(n_5263)
);


endmodule