module fake_jpeg_13645_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_19),
.B1(n_29),
.B2(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_56),
.B1(n_32),
.B2(n_18),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_19),
.B1(n_29),
.B2(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_93),
.B1(n_96),
.B2(n_58),
.Y(n_102)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_86),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_52),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_60),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_0),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_46),
.B1(n_45),
.B2(n_15),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_62),
.B1(n_65),
.B2(n_18),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_71),
.B(n_65),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_107),
.B(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_10),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_52),
.B(n_31),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_111),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_0),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_52),
.B(n_39),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_86),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_89),
.C(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.C(n_101),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_91),
.C(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_10),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_78),
.B1(n_93),
.B2(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_130),
.B1(n_109),
.B2(n_102),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_130),
.B1(n_108),
.B2(n_128),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_142),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_107),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_144),
.B(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.Y(n_157)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_119),
.C(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_151),
.C(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_129),
.C(n_112),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_101),
.C(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_160),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_125),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_140),
.C(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_165),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_152),
.B(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_159),
.C(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_125),
.Y(n_165)
);

NAND4xp25_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_105),
.C(n_14),
.D(n_11),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_106),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_134),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_112),
.B(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_114),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_173),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_105),
.Y(n_177)
);


endmodule