module fake_jpeg_10596_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_29),
.Y(n_36)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_22),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_15),
.B1(n_20),
.B2(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_19),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_45),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_19),
.B1(n_23),
.B2(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_48),
.B1(n_31),
.B2(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_39),
.C(n_27),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_60),
.C(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_47),
.B1(n_46),
.B2(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_55),
.B1(n_33),
.B2(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_15),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_51),
.B1(n_61),
.B2(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_85),
.B1(n_46),
.B2(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_75),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_69),
.C(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_64),
.C(n_37),
.Y(n_101)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_72),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_82),
.Y(n_95)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_3),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_63),
.B(n_73),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_85),
.B1(n_30),
.B2(n_76),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_89),
.B1(n_88),
.B2(n_33),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_105),
.C(n_98),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_82),
.C(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_3),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_3),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_115),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_101),
.C(n_102),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_96),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_114),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_96),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_103),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_99),
.C(n_13),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_99),
.Y(n_125)
);

NAND2x1_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_109),
.B1(n_104),
.B2(n_110),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_106),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_127),
.A3(n_12),
.B1(n_24),
.B2(n_121),
.C1(n_10),
.C2(n_9),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_13),
.B1(n_21),
.B2(n_17),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_126),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_4),
.A3(n_7),
.B1(n_33),
.B2(n_122),
.C1(n_121),
.C2(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_7),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_131),
.A2(n_132),
.B(n_128),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_122),
.Y(n_134)
);


endmodule