module fake_jpeg_22196_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_32),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_56),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_27),
.B1(n_17),
.B2(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_27),
.B1(n_17),
.B2(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_77),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_76),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_39),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_40),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_40),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

BUFx12f_ASAP7_75t_SL g90 ( 
.A(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_92),
.B1(n_41),
.B2(n_65),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_90),
.B1(n_83),
.B2(n_88),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_27),
.B1(n_54),
.B2(n_67),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_48),
.B1(n_27),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_35),
.B1(n_41),
.B2(n_33),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_109),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_21),
.B1(n_31),
.B2(n_16),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_113),
.B1(n_25),
.B2(n_23),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_33),
.C(n_38),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_73),
.C(n_77),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_31),
.B1(n_16),
.B2(n_41),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_34),
.Y(n_136)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_35),
.B1(n_33),
.B2(n_38),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_129),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_143),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_104),
.C(n_115),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_130),
.Y(n_157)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_85),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_137),
.B(n_34),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_86),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_72),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_146),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_144),
.B(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_96),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_101),
.B1(n_25),
.B2(n_23),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_39),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_104),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_163),
.B(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_117),
.B1(n_107),
.B2(n_112),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_168),
.B1(n_125),
.B2(n_122),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_124),
.Y(n_154)
);

AO21x2_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_75),
.B(n_76),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_161),
.B1(n_167),
.B2(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_148),
.C(n_126),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_104),
.B1(n_72),
.B2(n_80),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_116),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_75),
.B1(n_82),
.B2(n_94),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_76),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_82),
.B1(n_76),
.B2(n_94),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_127),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_123),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_128),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_176),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_157),
.B(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_186),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_197),
.C(n_169),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_142),
.C(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_91),
.C(n_70),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_196),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_133),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_193),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_137),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_91),
.B1(n_167),
.B2(n_121),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_196),
.A2(n_158),
.B(n_149),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_209),
.B(n_218),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_161),
.B1(n_172),
.B2(n_158),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_219),
.B1(n_63),
.B2(n_110),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_212),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_158),
.B(n_153),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_197),
.B(n_137),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_175),
.B(n_25),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_169),
.C(n_152),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_185),
.A2(n_125),
.B1(n_150),
.B2(n_171),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_226),
.B1(n_224),
.B2(n_223),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_181),
.B1(n_180),
.B2(n_182),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_201),
.A2(n_139),
.B(n_132),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_123),
.B1(n_134),
.B2(n_101),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_42),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_184),
.A2(n_185),
.B(n_178),
.C(n_194),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_199),
.B(n_190),
.C(n_198),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_96),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_39),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_186),
.A2(n_91),
.B1(n_70),
.B2(n_38),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_1),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_235),
.B1(n_240),
.B2(n_221),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_221),
.A2(n_199),
.B1(n_192),
.B2(n_187),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_229),
.A2(n_247),
.B(n_228),
.C(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_238),
.B1(n_245),
.B2(n_24),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_233),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_30),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_0),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_218),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_248),
.B(n_249),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_214),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_223),
.B1(n_215),
.B2(n_208),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_202),
.B(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_246),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_203),
.A2(n_209),
.B1(n_204),
.B2(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_213),
.B(n_19),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_29),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_165),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_165),
.B(n_131),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_212),
.C(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_255),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_207),
.C(n_227),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_211),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_216),
.C(n_131),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_268),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_28),
.CI(n_39),
.CON(n_262),
.SN(n_262)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_235),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_233),
.B(n_240),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_235),
.B(n_89),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_23),
.B1(n_110),
.B2(n_22),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_269),
.B1(n_24),
.B2(n_18),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_267)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_89),
.C(n_36),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_36),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_238),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_280),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_251),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_286),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_262),
.B(n_264),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_28),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_283),
.C(n_287),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_11),
.B(n_15),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_258),
.B(n_11),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_289),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_295),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_281),
.A2(n_264),
.B(n_262),
.C(n_256),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_280),
.B(n_274),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_254),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_302),
.B(n_8),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_252),
.C(n_255),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.C(n_2),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_268),
.C(n_253),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_310),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_271),
.B1(n_266),
.B2(n_270),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_304),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_42),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_9),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.C(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_28),
.C(n_18),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_18),
.C(n_24),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_9),
.B(n_13),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_8),
.C(n_13),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_313),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_10),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_296),
.B(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_293),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_291),
.C(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_323),
.C(n_313),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_327),
.C(n_328),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_303),
.Y(n_325)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_315),
.C(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_24),
.C(n_18),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_6),
.C(n_12),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_5),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_326),
.B(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_333),
.C(n_39),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_2),
.C(n_3),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_39),
.B(n_4),
.C(n_6),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_4),
.C(n_5),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_6),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_7),
.C(n_39),
.Y(n_341)
);


endmodule