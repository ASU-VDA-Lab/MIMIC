module fake_jpeg_11468_n_40 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_0),
.C(n_4),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_11),
.B(n_1),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_23),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_24),
.Y(n_25)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_18),
.B1(n_13),
.B2(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_23),
.C(n_7),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.C(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_28),
.C(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_6),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_23),
.B1(n_7),
.B2(n_8),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_37),
.B1(n_35),
.B2(n_9),
.Y(n_40)
);


endmodule