module fake_jpeg_18354_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_8),
.CON(n_40),
.SN(n_40)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_40),
.B(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_47),
.Y(n_82)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_9),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_0),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_74),
.Y(n_85)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_6),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_6),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_28),
.B(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_70),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_64),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_32),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_29),
.Y(n_98)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_32),
.B1(n_27),
.B2(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_99),
.B1(n_109),
.B2(n_62),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_30),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_21),
.B1(n_29),
.B2(n_23),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_102),
.B1(n_107),
.B2(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_14),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_72),
.B1(n_55),
.B2(n_52),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_21),
.B1(n_31),
.B2(n_16),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_70),
.B1(n_43),
.B2(n_68),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_21),
.B1(n_31),
.B2(n_16),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_37),
.B1(n_18),
.B2(n_35),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_46),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_39),
.B(n_37),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_35),
.B1(n_22),
.B2(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_39),
.B(n_22),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_44),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_24),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_118),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_117),
.A2(n_152),
.B1(n_88),
.B2(n_76),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_120),
.Y(n_164)
);

OA22x2_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_48),
.B1(n_69),
.B2(n_70),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_45),
.B1(n_48),
.B2(n_69),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_69),
.B1(n_22),
.B2(n_66),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_123),
.A2(n_151),
.B(n_86),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_44),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_124),
.B(n_155),
.CI(n_12),
.CON(n_191),
.SN(n_191)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_87),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_137),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_44),
.Y(n_137)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_88),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_41),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_153),
.C(n_49),
.Y(n_181)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_146),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_91),
.B1(n_81),
.B2(n_83),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_144),
.B1(n_150),
.B2(n_112),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_60),
.B1(n_56),
.B2(n_50),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_63),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_97),
.B(n_63),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_82),
.B(n_12),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_75),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_177),
.C(n_116),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_105),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_176),
.B(n_180),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_95),
.B1(n_110),
.B2(n_112),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_163),
.A2(n_174),
.B1(n_179),
.B2(n_192),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_183),
.B1(n_131),
.B2(n_154),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_110),
.B1(n_76),
.B2(n_78),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_105),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_108),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_178),
.A2(n_146),
.B1(n_148),
.B2(n_142),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_119),
.A2(n_78),
.B1(n_101),
.B2(n_86),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_101),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_190),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_93),
.B1(n_86),
.B2(n_103),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_120),
.A2(n_103),
.B(n_93),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_153),
.B(n_139),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_155),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_125),
.A2(n_60),
.B1(n_56),
.B2(n_50),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_193),
.B(n_201),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_120),
.B(n_143),
.C(n_123),
.D(n_124),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_194),
.A2(n_206),
.B(n_212),
.Y(n_252)
);

XNOR2x2_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_157),
.B(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_118),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_124),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_161),
.B(n_136),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_214),
.Y(n_230)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

AND2x4_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_120),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

NAND2x1_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_132),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_213),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_162),
.B(n_128),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_141),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_224),
.B1(n_227),
.B2(n_168),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_228),
.B1(n_179),
.B2(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_127),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_220),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_189),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_126),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_153),
.B1(n_147),
.B2(n_49),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_153),
.B1(n_84),
.B2(n_145),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_145),
.B1(n_130),
.B2(n_2),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_229),
.A2(n_234),
.B1(n_228),
.B2(n_209),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_231),
.B(n_235),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_211),
.B1(n_227),
.B2(n_224),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_183),
.B1(n_164),
.B2(n_168),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_162),
.Y(n_235)
);

NAND2x1_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_176),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_240),
.B(n_247),
.Y(n_267)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_164),
.A3(n_176),
.B1(n_160),
.B2(n_181),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_238),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_160),
.B1(n_174),
.B2(n_187),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_191),
.C(n_187),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_173),
.B(n_158),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_167),
.C(n_173),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_167),
.C(n_130),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_215),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_260),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_198),
.A2(n_158),
.B(n_159),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_212),
.B(n_206),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_213),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_130),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_198),
.B(n_220),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_265),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_260),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_277),
.B1(n_287),
.B2(n_240),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_236),
.B(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_229),
.B(n_234),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_232),
.A2(n_211),
.B1(n_199),
.B2(n_218),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_206),
.Y(n_278)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_222),
.B(n_194),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_285),
.B1(n_289),
.B2(n_230),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_251),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_280),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_258),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_193),
.B1(n_208),
.B2(n_216),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_284),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_210),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_195),
.B1(n_197),
.B2(n_172),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_237),
.A2(n_197),
.B1(n_172),
.B2(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_254),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_302),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_294),
.A2(n_255),
.B1(n_259),
.B2(n_256),
.Y(n_334)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_233),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_298),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_233),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_301),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_276),
.B1(n_274),
.B2(n_279),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_248),
.C(n_246),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_238),
.C(n_242),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_266),
.C(n_262),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_242),
.C(n_247),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_316),
.C(n_286),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_233),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_315),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_244),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_239),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_278),
.B(n_285),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_324),
.B(n_314),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_230),
.B1(n_270),
.B2(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_294),
.A2(n_290),
.B1(n_268),
.B2(n_235),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_305),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_278),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_278),
.C(n_289),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_326),
.C(n_329),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_288),
.C(n_272),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_275),
.C(n_277),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_280),
.C(n_283),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_308),
.C(n_316),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_304),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_333),
.Y(n_348)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_336),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_305),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_337),
.B(n_338),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_256),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_347),
.C(n_355),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_299),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_345),
.Y(n_361)
);

AO22x1_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_299),
.B1(n_313),
.B2(n_301),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_344),
.Y(n_366)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

AOI322xp5_ASAP7_75t_SL g344 ( 
.A1(n_328),
.A2(n_297),
.A3(n_298),
.B1(n_312),
.B2(n_315),
.C1(n_300),
.C2(n_302),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_309),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_323),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_241),
.C(n_259),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_327),
.A2(n_241),
.B1(n_221),
.B2(n_203),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_337),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_334),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_0),
.C(n_3),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_332),
.B(n_324),
.Y(n_357)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_328),
.Y(n_359)
);

AOI31xp33_ASAP7_75t_L g372 ( 
.A1(n_359),
.A2(n_360),
.A3(n_368),
.B(n_339),
.Y(n_372)
);

OAI221xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_318),
.B1(n_317),
.B2(n_325),
.C(n_319),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_363),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_354),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_329),
.C(n_323),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_339),
.C(n_346),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_369),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_367),
.B(n_330),
.Y(n_376)
);

XOR2x1_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_324),
.Y(n_368)
);

NOR2x1_ASAP7_75t_SL g378 ( 
.A(n_368),
.B(n_352),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_374),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_372),
.A2(n_4),
.B(n_5),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_345),
.C(n_341),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_377),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_355),
.C(n_330),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_362),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_366),
.B(n_348),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_381),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_352),
.B(n_351),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_380),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_3),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_385),
.Y(n_393)
);

AO21x1_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_359),
.B(n_364),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_4),
.B(n_10),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_370),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_361),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_389),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_15),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_11),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_SL g398 ( 
.A(n_391),
.B(n_11),
.C(n_13),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_373),
.B(n_377),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_394),
.B(n_396),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_374),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_4),
.B(n_11),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_382),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_398),
.B(n_399),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_400),
.B(n_402),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_390),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_395),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_384),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_405),
.Y(n_408)
);

AOI321xp33_ASAP7_75t_SL g407 ( 
.A1(n_404),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_401),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_406),
.C(n_407),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_14),
.C(n_15),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_15),
.Y(n_411)
);


endmodule