module fake_jpeg_550_n_192 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_22),
.B(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_13),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_56),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_72),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_58),
.B1(n_66),
.B2(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_59),
.B1(n_47),
.B2(n_63),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_89),
.Y(n_93)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_78),
.Y(n_104)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_50),
.B1(n_63),
.B2(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_58),
.B1(n_61),
.B2(n_51),
.Y(n_90)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_97),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_52),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_49),
.Y(n_120)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_60),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_61),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_67),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_0),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_88),
.B1(n_85),
.B2(n_84),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_107),
.B1(n_98),
.B2(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_101),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_80),
.B(n_47),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_49),
.B(n_4),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_64),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_3),
.C(n_4),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_124),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_49),
.B1(n_48),
.B2(n_57),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_1),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_2),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_2),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_49),
.B1(n_48),
.B2(n_57),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_147),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_143),
.Y(n_164)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR4xp25_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_44),
.C(n_43),
.D(n_42),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_3),
.B(n_5),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_40),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_120),
.B(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_150),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_154),
.B1(n_162),
.B2(n_166),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_39),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_38),
.B(n_33),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_165),
.B(n_134),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx4f_ASAP7_75t_SL g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_133),
.C(n_149),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_169),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_140),
.C(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_174),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_144),
.CI(n_138),
.CON(n_173),
.SN(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_18),
.C(n_32),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_161),
.B1(n_175),
.B2(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_153),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_158),
.B1(n_171),
.B2(n_163),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_187),
.A3(n_188),
.B1(n_157),
.B2(n_183),
.C1(n_185),
.C2(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_176),
.C(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_173),
.B1(n_166),
.B2(n_154),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_187),
.C(n_151),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_164),
.C(n_137),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.C(n_16),
.Y(n_192)
);


endmodule