module fake_ariane_2403_n_1655 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1655);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1655;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_10),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_13),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_77),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_67),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_44),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_33),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_44),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_107),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_81),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_38),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_1),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_54),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_38),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_50),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_2),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_108),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_92),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_79),
.Y(n_192)
);

BUFx8_ASAP7_75t_SL g193 ( 
.A(n_147),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_66),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_21),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_31),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_27),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_6),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_99),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_4),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_19),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_89),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_58),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_138),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_98),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_63),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_5),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_72),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_14),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_51),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_110),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_83),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_74),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_94),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_93),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_35),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_103),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_8),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_29),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_114),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_60),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_82),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_23),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_30),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_80),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_104),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_21),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_144),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_64),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_40),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_23),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_90),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_32),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_140),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_121),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_115),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_111),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_25),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_117),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_15),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_86),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_16),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_49),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_4),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_97),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_55),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_8),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_13),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_31),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_146),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_43),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_113),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_96),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_109),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_28),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_142),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_30),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_46),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_78),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_36),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_70),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_39),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_85),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_26),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_52),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_126),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_47),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_61),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_152),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_250),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_193),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_200),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_235),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_204),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_157),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_157),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_159),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_159),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_290),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_249),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_181),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_173),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_169),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_153),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_189),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_166),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_186),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_153),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_195),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_167),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_169),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_261),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_163),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_167),
.Y(n_338)
);

BUFx2_ASAP7_75t_SL g339 ( 
.A(n_163),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_172),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_177),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_215),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_215),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_196),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_222),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_222),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_244),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_198),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_244),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_183),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_199),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_187),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_191),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_272),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_202),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_249),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_281),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_212),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_224),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_203),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_259),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_266),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_279),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_284),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_163),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_264),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_277),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_210),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_300),
.A2(n_263),
.B1(n_245),
.B2(n_216),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_353),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_170),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_314),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_258),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_R g399 ( 
.A(n_304),
.B(n_180),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_313),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_324),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_303),
.A2(n_297),
.B1(n_220),
.B2(n_294),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_331),
.B(n_296),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_307),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_346),
.B(n_151),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_303),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_182),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_322),
.B(n_230),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_356),
.B(n_264),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_343),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_345),
.B(n_182),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_348),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_317),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_356),
.B(n_264),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_350),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_158),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_358),
.B(n_292),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_336),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_358),
.B(n_292),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_315),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_315),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_361),
.B(n_364),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_316),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_361),
.B(n_292),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_318),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_318),
.A2(n_162),
.B(n_161),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_355),
.B(n_175),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_357),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_405),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_379),
.B(n_312),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_405),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_379),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_411),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_379),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_405),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_418),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_339),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_418),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_L g461 ( 
.A1(n_376),
.A2(n_310),
.B1(n_321),
.B2(n_359),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_404),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_L g465 ( 
.A1(n_376),
.A2(n_403),
.B1(n_407),
.B2(n_411),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_399),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_392),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_374),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_425),
.B(n_330),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_425),
.B(n_362),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_413),
.B(n_338),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_425),
.A2(n_265),
.B1(n_268),
.B2(n_177),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_431),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_339),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_431),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_L g484 ( 
.A(n_399),
.B(n_333),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_443),
.A2(n_334),
.B1(n_341),
.B2(n_366),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_412),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_383),
.B(n_344),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_431),
.B(n_347),
.Y(n_493)
);

NAND2x1p5_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_402),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_434),
.B(n_351),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_385),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_386),
.Y(n_497)
);

INVx8_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_434),
.B(n_354),
.Y(n_499)
);

AND3x2_ASAP7_75t_L g500 ( 
.A(n_409),
.B(n_371),
.C(n_367),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_388),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_364),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_440),
.B(n_363),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_388),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g511 ( 
.A(n_407),
.B(n_373),
.C(n_265),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_440),
.B(n_367),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_368),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_443),
.A2(n_370),
.B1(n_369),
.B2(n_340),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_383),
.B(n_320),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_390),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_390),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_391),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_391),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_383),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_409),
.B(n_302),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_389),
.Y(n_526)
);

AND3x2_ASAP7_75t_L g527 ( 
.A(n_409),
.B(n_368),
.C(n_329),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_393),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_393),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_424),
.B(n_365),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_396),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_389),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_437),
.B(n_299),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_383),
.B(n_160),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_443),
.A2(n_421),
.B1(n_416),
.B2(n_394),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_389),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_394),
.B(n_154),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_384),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_402),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_437),
.B(n_319),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

CKINVDCx11_ASAP7_75t_R g549 ( 
.A(n_404),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_419),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_394),
.B(n_154),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_394),
.B(n_305),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_428),
.B(n_168),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_394),
.B(n_155),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_442),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_443),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_443),
.B(n_319),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_416),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_384),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_423),
.B(n_178),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_403),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_384),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_416),
.B(n_323),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_435),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_435),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_442),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_375),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_442),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_416),
.B(n_175),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_421),
.B(n_176),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_401),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_421),
.B(n_208),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_421),
.B(n_248),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_413),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_415),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_420),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_437),
.B(n_155),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_459),
.B(n_421),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_459),
.A2(n_417),
.B1(n_430),
.B2(n_429),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_524),
.B(n_429),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_471),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_524),
.B(n_156),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_566),
.A2(n_430),
.B1(n_417),
.B2(n_420),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_524),
.B(n_156),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_474),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_458),
.B(n_408),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_514),
.A2(n_478),
.B1(n_498),
.B2(n_560),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_453),
.B(n_408),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_559),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_476),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_524),
.B(n_164),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_498),
.B(n_458),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_508),
.B(n_164),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_460),
.B(n_410),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_410),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_566),
.A2(n_432),
.B1(n_422),
.B2(n_426),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_479),
.B(n_426),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_469),
.B(n_432),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_482),
.B(n_436),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_541),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_482),
.B(n_436),
.Y(n_615)
);

INVxp33_ASAP7_75t_L g616 ( 
.A(n_549),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_559),
.B(n_439),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_486),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_462),
.A2(n_360),
.B1(n_433),
.B2(n_444),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_490),
.Y(n_621)
);

BUFx6f_ASAP7_75t_SL g622 ( 
.A(n_473),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_467),
.B(n_309),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_567),
.B(n_268),
.C(n_220),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_514),
.A2(n_219),
.B1(n_174),
.B2(n_282),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_490),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_473),
.B(n_439),
.Y(n_627)
);

NAND2x1p5_ASAP7_75t_L g628 ( 
.A(n_561),
.B(n_441),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_473),
.B(n_441),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_498),
.B(n_165),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_508),
.B(n_171),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_473),
.B(n_171),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_567),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_557),
.B(n_174),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_498),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_557),
.B(n_219),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_543),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_496),
.Y(n_638)
);

BUFx5_ASAP7_75t_L g639 ( 
.A(n_573),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_498),
.B(n_262),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_453),
.B(n_223),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_496),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_455),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_480),
.B(n_262),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_456),
.B(n_232),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_561),
.A2(n_243),
.B(n_179),
.C(n_233),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_543),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_502),
.B(n_513),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_469),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_456),
.B(n_236),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_514),
.B(n_240),
.Y(n_652)
);

INVxp33_ASAP7_75t_L g653 ( 
.A(n_463),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_526),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_480),
.B(n_267),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_560),
.Y(n_656)
);

AND2x2_ASAP7_75t_SL g657 ( 
.A(n_540),
.B(n_185),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_497),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_557),
.B(n_274),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_502),
.B(n_274),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_513),
.B(n_278),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_537),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_492),
.B(n_278),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_526),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_526),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_526),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_526),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_480),
.B(n_293),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_481),
.A2(n_387),
.B(n_398),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_514),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_514),
.A2(n_294),
.B1(n_288),
.B2(n_271),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_472),
.B(n_242),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_584),
.B(n_323),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_576),
.B(n_211),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_573),
.A2(n_295),
.B1(n_192),
.B2(n_228),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_455),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_465),
.B(n_288),
.C(n_271),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_500),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_576),
.B(n_217),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_493),
.B(n_254),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_535),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_560),
.B(n_325),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_535),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_553),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_495),
.B(n_273),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_481),
.B(n_273),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_560),
.A2(n_218),
.B1(n_221),
.B2(n_225),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_501),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_499),
.B(n_275),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_R g690 ( 
.A(n_525),
.B(n_433),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_467),
.B(n_275),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_535),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_530),
.B(n_280),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_530),
.B(n_280),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_560),
.B(n_325),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_576),
.B(n_226),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_530),
.B(n_285),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_538),
.B(n_285),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_576),
.B(n_229),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_478),
.B(n_444),
.Y(n_700)
);

OAI21xp33_ASAP7_75t_L g701 ( 
.A1(n_555),
.A2(n_297),
.B(n_286),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_477),
.B(n_286),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_535),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_547),
.B(n_184),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_577),
.A2(n_582),
.B1(n_579),
.B2(n_586),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_527),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_547),
.B(n_578),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_477),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_505),
.B(n_246),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_580),
.B(n_188),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_494),
.B(n_252),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_484),
.B(n_192),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_535),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_583),
.B(n_190),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_537),
.B(n_194),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_R g716 ( 
.A(n_532),
.B(n_295),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_542),
.B(n_256),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_579),
.B(n_201),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_569),
.B(n_228),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_451),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_445),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_585),
.B(n_209),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_585),
.B(n_213),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_588),
.A2(n_270),
.B1(n_227),
.B2(n_239),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_569),
.B(n_231),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_569),
.B(n_234),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_517),
.B(n_0),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_569),
.B(n_237),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_518),
.Y(n_729)
);

BUFx8_ASAP7_75t_L g730 ( 
.A(n_577),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_574),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_569),
.B(n_238),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_564),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_494),
.B(n_230),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_551),
.B(n_0),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_577),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_494),
.B(n_230),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_577),
.A2(n_255),
.B1(n_257),
.B2(n_260),
.Y(n_738)
);

BUFx6f_ASAP7_75t_SL g739 ( 
.A(n_577),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_489),
.B(n_295),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_656),
.B(n_556),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_721),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_676),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_635),
.B(n_536),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_601),
.B(n_488),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_736),
.Y(n_746)
);

OR2x2_ASAP7_75t_SL g747 ( 
.A(n_727),
.B(n_511),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_601),
.B(n_707),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_656),
.B(n_564),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_635),
.B(n_536),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_598),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_591),
.A2(n_529),
.B(n_501),
.C(n_506),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_736),
.B(n_564),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_662),
.B(n_577),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_708),
.B(n_461),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_736),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_603),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_612),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_734),
.A2(n_503),
.B(n_491),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_643),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_618),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_639),
.B(n_544),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_702),
.B(n_534),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_633),
.B(n_534),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_639),
.B(n_600),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_622),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_599),
.B(n_577),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_607),
.B(n_489),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_674),
.A2(n_544),
.B(n_546),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_620),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_650),
.B(n_555),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_730),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_621),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_684),
.B(n_539),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_639),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_626),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_638),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_639),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_642),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_658),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_639),
.Y(n_782)
);

XNOR2xp5_ASAP7_75t_L g783 ( 
.A(n_619),
.B(n_565),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_608),
.B(n_489),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_589),
.B(n_491),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_622),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_690),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_739),
.B(n_548),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_690),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_R g790 ( 
.A(n_623),
.B(n_503),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_657),
.A2(n_550),
.B1(n_554),
.B2(n_562),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_600),
.B(n_705),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_730),
.Y(n_793)
);

INVx5_ASAP7_75t_L g794 ( 
.A(n_682),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_688),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_649),
.B(n_548),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_657),
.B(n_552),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_628),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_653),
.B(n_550),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_629),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_731),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_660),
.B(n_565),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_677),
.A2(n_506),
.B1(n_519),
.B2(n_520),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_627),
.B(n_558),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_590),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_661),
.B(n_558),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_682),
.B(n_519),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_695),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_695),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_719),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_720),
.B(n_520),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_712),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_L g813 ( 
.A(n_733),
.B(n_523),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_641),
.B(n_554),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_735),
.A2(n_675),
.B1(n_717),
.B2(n_652),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_592),
.Y(n_816)
);

HB1xp67_ASAP7_75t_SL g817 ( 
.A(n_678),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_610),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_641),
.B(n_562),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_719),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_628),
.B(n_507),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_613),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_729),
.B(n_523),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_615),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_617),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_693),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_737),
.A2(n_448),
.B(n_449),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_SL g828 ( 
.A(n_624),
.B(n_529),
.C(n_531),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_614),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_637),
.B(n_531),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_646),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_596),
.B(n_507),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_648),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_593),
.B(n_522),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_645),
.B(n_509),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_611),
.B(n_522),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_694),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_L g838 ( 
.A(n_715),
.B(n_574),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_739),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_652),
.A2(n_528),
.B1(n_533),
.B2(n_575),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_645),
.B(n_509),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_735),
.A2(n_528),
.B1(n_533),
.B2(n_575),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_654),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_673),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_669),
.A2(n_470),
.B(n_448),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_593),
.B(n_510),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_664),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_665),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_675),
.A2(n_587),
.B1(n_581),
.B2(n_510),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_651),
.B(n_512),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_717),
.A2(n_587),
.B1(n_581),
.B2(n_512),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_709),
.A2(n_515),
.B1(n_572),
.B2(n_571),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_SL g853 ( 
.A(n_663),
.B(n_515),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_716),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_716),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_651),
.B(n_516),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_667),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_704),
.B(n_516),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_681),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_632),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_602),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_691),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_697),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_706),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_683),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_596),
.B(n_521),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_686),
.B(n_521),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_709),
.B(n_570),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_692),
.B(n_574),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_671),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_663),
.B(n_570),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_703),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_698),
.B(n_685),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_725),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_726),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_728),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_713),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_732),
.B(n_572),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_625),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_710),
.B(n_714),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_670),
.B(n_446),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_674),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_609),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_679),
.Y(n_885)
);

AO22x1_ASAP7_75t_L g886 ( 
.A1(n_616),
.A2(n_447),
.B1(n_454),
.B2(n_449),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_740),
.Y(n_887)
);

BUFx8_ASAP7_75t_L g888 ( 
.A(n_685),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_605),
.B(n_630),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_718),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_689),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_679),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_689),
.A2(n_450),
.B1(n_452),
.B2(n_454),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_701),
.B(n_450),
.Y(n_894)
);

BUFx12f_ASAP7_75t_L g895 ( 
.A(n_672),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_672),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_687),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_680),
.B(n_452),
.Y(n_898)
);

AO22x1_ASAP7_75t_L g899 ( 
.A1(n_680),
.A2(n_464),
.B1(n_457),
.B2(n_466),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_696),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_SL g901 ( 
.A1(n_724),
.A2(n_269),
.B1(n_214),
.B2(n_189),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_696),
.A2(n_468),
.B1(n_457),
.B2(n_464),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_595),
.B(n_466),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_699),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_699),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_711),
.B(n_470),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_722),
.B(n_475),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_595),
.B(n_475),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_723),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_895),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_748),
.B(n_597),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_794),
.B(n_896),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_891),
.A2(n_647),
.B(n_631),
.C(n_634),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_743),
.B(n_604),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_790),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_745),
.B(n_604),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_761),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_815),
.A2(n_631),
.B1(n_606),
.B2(n_659),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_SL g919 ( 
.A(n_794),
.B(n_640),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_SL g920 ( 
.A1(n_770),
.A2(n_644),
.B(n_655),
.C(n_668),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_874),
.B(n_606),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_790),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_845),
.A2(n_737),
.B(n_483),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_750),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_792),
.A2(n_636),
.B(n_659),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_754),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_820),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_854),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_752),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_890),
.A2(n_504),
.B(n_487),
.C(n_485),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_SL g931 ( 
.A1(n_823),
.A2(n_485),
.B(n_487),
.C(n_504),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_SL g932 ( 
.A1(n_880),
.A2(n_738),
.B1(n_269),
.B2(n_214),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_794),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_897),
.B(n_545),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_897),
.B(n_545),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_794),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_R g937 ( 
.A(n_855),
.B(n_789),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_810),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_823),
.A2(n_563),
.B(n_545),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_L g940 ( 
.A1(n_815),
.A2(n_563),
.B(n_545),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_746),
.B(n_189),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_755),
.B(n_563),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_827),
.A2(n_381),
.B(n_398),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_871),
.A2(n_563),
.B1(n_230),
.B2(n_375),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_767),
.B(n_563),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_792),
.A2(n_189),
.B1(n_214),
.B2(n_269),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_810),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_769),
.A2(n_568),
.B(n_398),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_754),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_742),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_758),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_808),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_784),
.A2(n_568),
.B(n_382),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_763),
.A2(n_568),
.B(n_382),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_759),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_783),
.A2(n_230),
.B1(n_375),
.B2(n_568),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_811),
.A2(n_377),
.B(n_378),
.C(n_387),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_766),
.A2(n_214),
.B1(n_269),
.B2(n_375),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_818),
.B(n_9),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_755),
.B(n_378),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_786),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_822),
.B(n_11),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_807),
.A2(n_825),
.B1(n_824),
.B2(n_803),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_773),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_756),
.B(n_12),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_811),
.B(n_14),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_775),
.B(n_15),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_809),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_766),
.A2(n_214),
.B1(n_269),
.B2(n_375),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_762),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_875),
.B(n_16),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_861),
.B(n_17),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_754),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_861),
.B(n_17),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_771),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_876),
.B(n_18),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_773),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_834),
.A2(n_753),
.B(n_828),
.C(n_909),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_834),
.A2(n_377),
.B(n_387),
.C(n_381),
.Y(n_979)
);

OAI22x1_ASAP7_75t_L g980 ( 
.A1(n_877),
.A2(n_377),
.B1(n_20),
.B2(n_22),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_799),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_787),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_802),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_SL g984 ( 
.A1(n_753),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_813),
.A2(n_837),
.B(n_864),
.C(n_826),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_793),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_828),
.A2(n_397),
.B(n_395),
.C(n_384),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_817),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_888),
.A2(n_230),
.B1(n_395),
.B2(n_384),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_764),
.B(n_28),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_763),
.A2(n_397),
.B(n_395),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_909),
.A2(n_397),
.B(n_395),
.C(n_384),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_793),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_774),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_767),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_749),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_777),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_786),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_844),
.A2(n_835),
.B(n_841),
.C(n_850),
.Y(n_999)
);

INVx3_ASAP7_75t_SL g1000 ( 
.A(n_863),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_778),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_856),
.A2(n_397),
.B(n_395),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_801),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_800),
.B(n_29),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_765),
.B(n_32),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_884),
.A2(n_397),
.B1(n_384),
.B2(n_36),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_780),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_888),
.A2(n_397),
.B1(n_35),
.B2(n_37),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_772),
.B(n_34),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_908),
.A2(n_34),
.B(n_41),
.C(n_42),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_797),
.A2(n_862),
.B1(n_804),
.B2(n_842),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_844),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_842),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_801),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_865),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_908),
.A2(n_56),
.B(n_57),
.C(n_59),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_749),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_781),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_901),
.A2(n_76),
.B1(n_95),
.B2(n_101),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_747),
.B(n_118),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_801),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_776),
.A2(n_128),
.B(n_133),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_796),
.A2(n_134),
.B1(n_141),
.B2(n_148),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_746),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_SL g1025 ( 
.A1(n_744),
.A2(n_149),
.B(n_751),
.C(n_785),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_812),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_832),
.A2(n_867),
.B(n_760),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_795),
.B(n_836),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_779),
.A2(n_782),
.B(n_907),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_836),
.B(n_741),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_846),
.A2(n_768),
.B(n_887),
.C(n_819),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_806),
.B(n_741),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_882),
.A2(n_846),
.B1(n_887),
.B2(n_798),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_833),
.B(n_801),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_SL g1035 ( 
.A(n_746),
.B(n_788),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_878),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_878),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_963),
.B(n_798),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_939),
.A2(n_782),
.B(n_779),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_988),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_916),
.B(n_886),
.Y(n_1041)
);

NAND3x1_ASAP7_75t_L g1042 ( 
.A(n_1020),
.B(n_840),
.C(n_839),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_982),
.B(n_833),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_SL g1044 ( 
.A1(n_911),
.A2(n_814),
.B(n_872),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_966),
.A2(n_889),
.B(n_859),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_924),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_923),
.A2(n_943),
.B(n_1002),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_965),
.B(n_882),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_918),
.A2(n_899),
.B(n_906),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_978),
.A2(n_913),
.B(n_751),
.C(n_744),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_921),
.B(n_869),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_918),
.A2(n_898),
.B(n_868),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_938),
.B(n_903),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_996),
.B(n_839),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_999),
.A2(n_853),
.B(n_821),
.Y(n_1055)
);

AO31x2_ASAP7_75t_L g1056 ( 
.A1(n_925),
.A2(n_1031),
.A3(n_958),
.B(n_969),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_940),
.A2(n_852),
.B1(n_791),
.B2(n_851),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_947),
.B(n_873),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1033),
.B(n_934),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_996),
.B(n_746),
.Y(n_1060)
);

OAI22x1_ASAP7_75t_L g1061 ( 
.A1(n_914),
.A2(n_905),
.B1(n_904),
.B2(n_900),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_L g1062 ( 
.A(n_936),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_L g1063 ( 
.A(n_983),
.B(n_838),
.C(n_904),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_935),
.B(n_905),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_922),
.B(n_889),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_922),
.B(n_829),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_910),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_958),
.A2(n_892),
.A3(n_885),
.B(n_883),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_964),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_941),
.A2(n_919),
.B(n_1025),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_941),
.A2(n_892),
.B(n_902),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_969),
.A2(n_894),
.A3(n_860),
.B(n_866),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_929),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_981),
.B(n_1037),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1027),
.A2(n_893),
.B(n_902),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_950),
.Y(n_1076)
);

AO21x1_ASAP7_75t_L g1077 ( 
.A1(n_1011),
.A2(n_830),
.B(n_870),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_951),
.Y(n_1078)
);

OA21x2_ASAP7_75t_L g1079 ( 
.A1(n_1027),
.A2(n_849),
.B(n_866),
.Y(n_1079)
);

AO21x1_ASAP7_75t_L g1080 ( 
.A1(n_985),
.A2(n_870),
.B(n_847),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1000),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_936),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1032),
.B(n_831),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_992),
.A2(n_847),
.A3(n_860),
.B(n_843),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_920),
.A2(n_879),
.B(n_843),
.Y(n_1085)
);

AOI211x1_ASAP7_75t_L g1086 ( 
.A1(n_972),
.A2(n_879),
.B(n_858),
.C(n_873),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_936),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_910),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_987),
.A2(n_879),
.B(n_829),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_971),
.A2(n_858),
.B(n_805),
.C(n_816),
.Y(n_1090)
);

CKINVDCx11_ASAP7_75t_R g1091 ( 
.A(n_1026),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1005),
.B(n_805),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_959),
.A2(n_816),
.B1(n_848),
.B2(n_757),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_955),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_915),
.B(n_857),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_991),
.A2(n_788),
.B(n_857),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1003),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1023),
.A2(n_1016),
.B(n_930),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_SL g1099 ( 
.A1(n_1009),
.A2(n_788),
.B(n_857),
.C(n_1023),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_1028),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_948),
.A2(n_953),
.B(n_954),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1036),
.B(n_982),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_927),
.B(n_1015),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_SL g1104 ( 
.A1(n_1010),
.A2(n_931),
.B(n_962),
.C(n_1004),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_952),
.B(n_968),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1022),
.A2(n_973),
.B(n_1024),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_998),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_979),
.A2(n_957),
.B(n_946),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1035),
.A2(n_942),
.B(n_984),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_917),
.B(n_961),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_990),
.A2(n_967),
.B(n_1006),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1035),
.A2(n_997),
.B(n_975),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_976),
.B(n_1017),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_974),
.B(n_994),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_970),
.A2(n_1007),
.B(n_1018),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1001),
.B(n_1017),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_926),
.A2(n_949),
.B(n_1034),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_926),
.A2(n_949),
.B(n_945),
.Y(n_1118)
);

AOI31xp67_ASAP7_75t_L g1119 ( 
.A1(n_989),
.A2(n_944),
.A3(n_956),
.B(n_912),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1030),
.B(n_928),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_960),
.A2(n_933),
.B(n_932),
.C(n_1019),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_980),
.A2(n_1013),
.A3(n_926),
.B(n_949),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_945),
.A2(n_1021),
.B(n_1012),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1014),
.B(n_1003),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1014),
.B(n_1003),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_945),
.A2(n_1014),
.B(n_1008),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_R g1127 ( 
.A(n_928),
.B(n_964),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_995),
.A2(n_937),
.B(n_977),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_977),
.A2(n_986),
.B(n_993),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_977),
.B(n_986),
.Y(n_1130)
);

NAND3x1_ASAP7_75t_L g1131 ( 
.A(n_993),
.B(n_677),
.C(n_1020),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_R g1132 ( 
.A(n_993),
.B(n_549),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_SL g1133 ( 
.A1(n_966),
.A2(n_911),
.B(n_881),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_925),
.A2(n_918),
.A3(n_1029),
.B(n_1031),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_916),
.B(n_748),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_L g1136 ( 
.A(n_917),
.B(n_650),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1020),
.B(n_896),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_923),
.A2(n_845),
.B(n_943),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_922),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_936),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_924),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_934),
.Y(n_1142)
);

OAI22x1_ASAP7_75t_L g1143 ( 
.A1(n_1020),
.A2(n_896),
.B1(n_783),
.B2(n_727),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_966),
.A2(n_911),
.B(n_881),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_918),
.A2(n_916),
.B(n_978),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_916),
.B(n_748),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_916),
.B(n_748),
.Y(n_1147)
);

INVxp67_ASAP7_75t_SL g1148 ( 
.A(n_934),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_924),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_925),
.A2(n_918),
.A3(n_1029),
.B(n_1031),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_966),
.A2(n_815),
.B1(n_600),
.B2(n_748),
.Y(n_1151)
);

INVx5_ASAP7_75t_L g1152 ( 
.A(n_936),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_932),
.A2(n_700),
.B1(n_815),
.B2(n_619),
.Y(n_1153)
);

AOI221x1_ASAP7_75t_L g1154 ( 
.A1(n_918),
.A2(n_932),
.B1(n_1020),
.B2(n_1010),
.C(n_940),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_916),
.B(n_748),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_925),
.A2(n_918),
.A3(n_1029),
.B(n_1031),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_923),
.A2(n_845),
.B(n_943),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_963),
.A2(n_911),
.B(n_985),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_916),
.B(n_748),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1020),
.B(n_896),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_996),
.B(n_794),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_925),
.A2(n_918),
.B(n_766),
.Y(n_1162)
);

NAND2x1_ASAP7_75t_L g1163 ( 
.A(n_1158),
.B(n_1044),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1069),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1137),
.A2(n_1160),
.B1(n_1143),
.B2(n_1151),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1098),
.A2(n_1145),
.B(n_1070),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1134),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1047),
.A2(n_1157),
.B(n_1138),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1145),
.A2(n_1151),
.B(n_1135),
.C(n_1155),
.Y(n_1169)
);

AOI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1153),
.A2(n_1111),
.B1(n_1159),
.B2(n_1146),
.C(n_1147),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1067),
.B(n_1088),
.Y(n_1171)
);

OAI22x1_ASAP7_75t_L g1172 ( 
.A1(n_1139),
.A2(n_1078),
.B1(n_1073),
.B2(n_1149),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1049),
.A2(n_1055),
.B(n_1085),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1135),
.B(n_1147),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1106),
.A2(n_1096),
.B(n_1039),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_1052),
.A2(n_1080),
.B(n_1075),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1094),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1154),
.A2(n_1093),
.B(n_1109),
.Y(n_1178)
);

AO21x2_ASAP7_75t_L g1179 ( 
.A1(n_1052),
.A2(n_1075),
.B(n_1077),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1111),
.A2(n_1112),
.B(n_1038),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1089),
.A2(n_1071),
.B(n_1045),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1087),
.B(n_1152),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1057),
.A2(n_1093),
.B(n_1064),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1133),
.A2(n_1144),
.B(n_1099),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1155),
.A2(n_1045),
.B(n_1051),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1141),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1079),
.A2(n_1064),
.B(n_1118),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1131),
.A2(n_1107),
.B1(n_1051),
.B2(n_1113),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1079),
.A2(n_1057),
.B(n_1123),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1117),
.A2(n_1108),
.B(n_1126),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1059),
.A2(n_1041),
.B(n_1090),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1081),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1108),
.A2(n_1115),
.B(n_1042),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_SL g1195 ( 
.A(n_1040),
.B(n_1065),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1086),
.B(n_1059),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1103),
.Y(n_1197)
);

INVxp67_ASAP7_75t_SL g1198 ( 
.A(n_1142),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1087),
.B(n_1152),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1130),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1091),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_1148),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1124),
.A2(n_1125),
.B(n_1116),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1124),
.A2(n_1125),
.B(n_1121),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1105),
.Y(n_1205)
);

AO21x2_ASAP7_75t_L g1206 ( 
.A1(n_1063),
.A2(n_1104),
.B(n_1162),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1162),
.A2(n_1092),
.B1(n_1100),
.B2(n_1114),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1050),
.A2(n_1083),
.B(n_1066),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1062),
.A2(n_1060),
.B(n_1095),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1061),
.A2(n_1102),
.B(n_1074),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1072),
.A2(n_1156),
.B(n_1150),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1119),
.A2(n_1043),
.B(n_1110),
.Y(n_1212)
);

AND2x2_ASAP7_75t_SL g1213 ( 
.A(n_1062),
.B(n_1161),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1120),
.A2(n_1139),
.B1(n_1058),
.B2(n_1127),
.C(n_1130),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1128),
.A2(n_1129),
.B(n_1084),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1084),
.A2(n_1150),
.B(n_1156),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1136),
.A2(n_1161),
.B1(n_1054),
.B2(n_1060),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1054),
.A2(n_1140),
.B1(n_1082),
.B2(n_1152),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1097),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1082),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1097),
.A2(n_1140),
.B1(n_1082),
.B2(n_1132),
.C(n_1122),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1140),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1084),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1122),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1122),
.A2(n_1056),
.B1(n_1150),
.B2(n_1156),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1056),
.B(n_1068),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1072),
.A2(n_1056),
.B(n_1068),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1072),
.A2(n_1047),
.B(n_1138),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1068),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1157),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1047),
.A2(n_1157),
.B(n_1138),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_SL g1232 ( 
.A1(n_1145),
.A2(n_1158),
.B(n_1151),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1157),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1118),
.B(n_1117),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1046),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_L g1236 ( 
.A(n_1087),
.B(n_789),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_SL g1237 ( 
.A1(n_1145),
.A2(n_1158),
.B(n_1151),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1047),
.A2(n_1101),
.B(n_1138),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1080),
.A2(n_925),
.A3(n_1077),
.B(n_1154),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1080),
.A2(n_925),
.A3(n_1077),
.B(n_1154),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1137),
.A2(n_1160),
.B1(n_815),
.B2(n_896),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1134),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1046),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1145),
.A2(n_1020),
.B(n_916),
.C(n_1151),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1157),
.Y(n_1245)
);

OR2x6_ASAP7_75t_L g1246 ( 
.A(n_1118),
.B(n_1117),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1046),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1047),
.A2(n_1101),
.B(n_1138),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1157),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1047),
.A2(n_1101),
.B(n_1138),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1046),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1134),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1081),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1134),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1097),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1098),
.A2(n_766),
.B(n_1145),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1081),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1076),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1047),
.A2(n_1101),
.B(n_1138),
.Y(n_1259)
);

AO22x1_ASAP7_75t_L g1260 ( 
.A1(n_1137),
.A2(n_1160),
.B1(n_888),
.B2(n_896),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1153),
.A2(n_815),
.B1(n_1143),
.B2(n_657),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1046),
.Y(n_1262)
);

OAI221xp5_ASAP7_75t_L g1263 ( 
.A1(n_1137),
.A2(n_896),
.B1(n_1160),
.B2(n_891),
.C(n_684),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1046),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1046),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1151),
.A2(n_1145),
.B1(n_600),
.B2(n_1135),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1146),
.B(n_1159),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1146),
.B(n_1159),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1157),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1047),
.A2(n_1138),
.B(n_1157),
.Y(n_1270)
);

AOI22x1_ASAP7_75t_L g1271 ( 
.A1(n_1145),
.A2(n_469),
.B1(n_650),
.B2(n_896),
.Y(n_1271)
);

CKINVDCx12_ASAP7_75t_R g1272 ( 
.A(n_1132),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1137),
.A2(n_1160),
.B(n_891),
.C(n_684),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1171),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1244),
.A2(n_1241),
.B(n_1169),
.C(n_1232),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1165),
.A2(n_1217),
.B1(n_1196),
.B2(n_1212),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1205),
.B(n_1174),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1244),
.A2(n_1261),
.B1(n_1169),
.B2(n_1263),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1272),
.A2(n_1201),
.B1(n_1261),
.B2(n_1189),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1205),
.B(n_1172),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1187),
.B(n_1197),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1256),
.A2(n_1271),
.B1(n_1266),
.B2(n_1170),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1213),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1237),
.A2(n_1266),
.B(n_1273),
.C(n_1166),
.Y(n_1284)
);

OAI31xp33_ASAP7_75t_L g1285 ( 
.A1(n_1267),
.A2(n_1268),
.A3(n_1257),
.B(n_1253),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1198),
.A2(n_1202),
.B1(n_1185),
.B2(n_1193),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1177),
.Y(n_1287)
);

OR2x6_ASAP7_75t_L g1288 ( 
.A(n_1234),
.B(n_1246),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1163),
.A2(n_1208),
.B(n_1206),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1242),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1180),
.A2(n_1179),
.B(n_1176),
.C(n_1254),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1203),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1176),
.A2(n_1242),
.B(n_1254),
.C(n_1252),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1227),
.A2(n_1228),
.B(n_1216),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1186),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1252),
.A2(n_1196),
.B(n_1243),
.C(n_1251),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_L g1297 ( 
.A1(n_1178),
.A2(n_1173),
.B(n_1260),
.C(n_1226),
.Y(n_1297)
);

OR2x6_ASAP7_75t_L g1298 ( 
.A(n_1234),
.B(n_1246),
.Y(n_1298)
);

AOI211xp5_ASAP7_75t_L g1299 ( 
.A1(n_1214),
.A2(n_1195),
.B(n_1221),
.C(n_1224),
.Y(n_1299)
);

AOI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1225),
.A2(n_1235),
.B1(n_1247),
.B2(n_1262),
.C(n_1264),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1196),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1265),
.B(n_1200),
.Y(n_1302)
);

OAI31xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1194),
.A2(n_1184),
.A3(n_1190),
.B(n_1204),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1182),
.A2(n_1199),
.B(n_1192),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1171),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1207),
.B(n_1183),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1238),
.A2(n_1250),
.B(n_1248),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1238),
.A2(n_1248),
.B(n_1259),
.Y(n_1309)
);

INVx3_ASAP7_75t_SL g1310 ( 
.A(n_1201),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1225),
.A2(n_1213),
.B1(n_1207),
.B2(n_1218),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1250),
.A2(n_1259),
.B(n_1190),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1209),
.B(n_1255),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1236),
.A2(n_1181),
.B1(n_1220),
.B2(n_1224),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1194),
.Y(n_1315)
);

INVxp67_ASAP7_75t_SL g1316 ( 
.A(n_1211),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1181),
.A2(n_1199),
.B1(n_1182),
.B2(n_1234),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1168),
.A2(n_1270),
.B(n_1269),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1231),
.A2(n_1245),
.B(n_1230),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1233),
.A2(n_1249),
.B(n_1175),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1191),
.A2(n_1188),
.B(n_1223),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1210),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1246),
.A2(n_1211),
.B1(n_1229),
.B2(n_1258),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1258),
.B(n_1239),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1211),
.A2(n_1231),
.B(n_1239),
.C(n_1240),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_R g1326 ( 
.A(n_1229),
.B(n_1239),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1215),
.B(n_1188),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1240),
.B(n_1187),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1198),
.B(n_1202),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1244),
.A2(n_1151),
.B(n_1154),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1187),
.B(n_1197),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1165),
.A2(n_1160),
.B1(n_1137),
.B2(n_1244),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1205),
.B(n_1174),
.Y(n_1333)
);

NOR2xp67_ASAP7_75t_L g1334 ( 
.A(n_1205),
.B(n_1172),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1166),
.A2(n_1256),
.B(n_1098),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1167),
.Y(n_1336)
);

O2A1O1Ixp5_ASAP7_75t_L g1337 ( 
.A1(n_1244),
.A2(n_1166),
.B(n_1145),
.C(n_1256),
.Y(n_1337)
);

CKINVDCx6p67_ASAP7_75t_R g1338 ( 
.A(n_1272),
.Y(n_1338)
);

O2A1O1Ixp5_ASAP7_75t_L g1339 ( 
.A1(n_1244),
.A2(n_1166),
.B(n_1145),
.C(n_1256),
.Y(n_1339)
);

O2A1O1Ixp5_ASAP7_75t_L g1340 ( 
.A1(n_1244),
.A2(n_1166),
.B(n_1145),
.C(n_1256),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1164),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1187),
.B(n_1197),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1166),
.A2(n_1256),
.B(n_1098),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1277),
.B(n_1333),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1328),
.B(n_1329),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_R g1346 ( 
.A(n_1274),
.B(n_1338),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1295),
.B(n_1290),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1288),
.B(n_1298),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1287),
.Y(n_1349)
);

BUFx2_ASAP7_75t_SL g1350 ( 
.A(n_1280),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1288),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1335),
.A2(n_1343),
.B(n_1275),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1286),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1324),
.Y(n_1354)
);

AOI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1289),
.A2(n_1322),
.B(n_1319),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1290),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1327),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1302),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1292),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1341),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1332),
.A2(n_1337),
.B(n_1339),
.Y(n_1361)
);

AO21x2_ASAP7_75t_L g1362 ( 
.A1(n_1316),
.A2(n_1326),
.B(n_1308),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1310),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1336),
.B(n_1307),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1336),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1308),
.A2(n_1325),
.B(n_1291),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1306),
.B(n_1310),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1281),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1331),
.B(n_1342),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1304),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1315),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1315),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1337),
.B(n_1339),
.Y(n_1373)
);

INVx4_ASAP7_75t_SL g1374 ( 
.A(n_1317),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1294),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1325),
.A2(n_1291),
.B(n_1323),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1340),
.A2(n_1282),
.B(n_1278),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1294),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1301),
.B(n_1343),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1300),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1293),
.Y(n_1381)
);

OR2x6_ASAP7_75t_L g1382 ( 
.A(n_1335),
.B(n_1305),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1293),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1340),
.A2(n_1275),
.B(n_1284),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1353),
.B(n_1334),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1371),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1356),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1375),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1375),
.B(n_1312),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1371),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1373),
.B(n_1296),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1347),
.B(n_1321),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1357),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1378),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1378),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1349),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1345),
.B(n_1309),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1365),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1354),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1361),
.A2(n_1297),
.B(n_1313),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1354),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1370),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1370),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1364),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1347),
.B(n_1321),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1373),
.B(n_1318),
.Y(n_1406)
);

INVx4_ASAP7_75t_L g1407 ( 
.A(n_1382),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1344),
.B(n_1296),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1359),
.Y(n_1409)
);

AO22x1_ASAP7_75t_L g1410 ( 
.A1(n_1377),
.A2(n_1311),
.B1(n_1283),
.B2(n_1314),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1364),
.B(n_1320),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1391),
.A2(n_1384),
.B(n_1352),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1391),
.A2(n_1381),
.B(n_1383),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1388),
.A2(n_1381),
.B(n_1383),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1393),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1410),
.A2(n_1355),
.B(n_1372),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1385),
.A2(n_1284),
.B1(n_1352),
.B2(n_1276),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1408),
.B(n_1369),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1402),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1385),
.A2(n_1276),
.B1(n_1380),
.B2(n_1279),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1402),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1387),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1398),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1399),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1393),
.Y(n_1425)
);

OAI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1408),
.A2(n_1380),
.B1(n_1285),
.B2(n_1299),
.C(n_1330),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1393),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1399),
.Y(n_1428)
);

NOR4xp25_ASAP7_75t_SL g1429 ( 
.A(n_1404),
.B(n_1363),
.C(n_1372),
.D(n_1351),
.Y(n_1429)
);

OAI33xp33_ASAP7_75t_L g1430 ( 
.A1(n_1392),
.A2(n_1358),
.A3(n_1405),
.B1(n_1411),
.B2(n_1368),
.B3(n_1396),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1399),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1402),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1389),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1410),
.A2(n_1350),
.B1(n_1374),
.B2(n_1376),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1389),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_SL g1436 ( 
.A(n_1398),
.B(n_1346),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1400),
.A2(n_1376),
.B1(n_1350),
.B2(n_1382),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1389),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1401),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1401),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1400),
.A2(n_1297),
.B(n_1379),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1389),
.Y(n_1442)
);

AOI211xp5_ASAP7_75t_L g1443 ( 
.A1(n_1406),
.A2(n_1379),
.B(n_1303),
.C(n_1367),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1404),
.B(n_1369),
.Y(n_1444)
);

INVx5_ASAP7_75t_L g1445 ( 
.A(n_1407),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1401),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1386),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1422),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1418),
.B(n_1392),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1443),
.B(n_1397),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1424),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1416),
.B(n_1382),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1433),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1424),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1416),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1433),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1428),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1412),
.B(n_1402),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1433),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1428),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1435),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1441),
.B(n_1348),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1412),
.A2(n_1434),
.B(n_1417),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1431),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1413),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1436),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1445),
.B(n_1407),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1413),
.B(n_1392),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1443),
.B(n_1397),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1445),
.B(n_1407),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1415),
.Y(n_1472)
);

NOR2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1421),
.B(n_1403),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1413),
.B(n_1392),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1434),
.B(n_1403),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1438),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1413),
.B(n_1409),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1421),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1437),
.A2(n_1394),
.B(n_1395),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1444),
.B(n_1405),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1449),
.B(n_1480),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1450),
.B(n_1421),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1450),
.A2(n_1426),
.B1(n_1420),
.B2(n_1376),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1451),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1467),
.Y(n_1485)
);

AOI222xp33_ASAP7_75t_L g1486 ( 
.A1(n_1470),
.A2(n_1430),
.B1(n_1466),
.B2(n_1475),
.C1(n_1406),
.C2(n_1477),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

OAI33xp33_ASAP7_75t_L g1488 ( 
.A1(n_1469),
.A2(n_1405),
.A3(n_1446),
.B1(n_1440),
.B2(n_1439),
.B3(n_1411),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1451),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1470),
.A2(n_1400),
.B1(n_1366),
.B2(n_1362),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1454),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1467),
.B(n_1432),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1406),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1454),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1458),
.B(n_1406),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1473),
.B(n_1432),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1473),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1478),
.B(n_1432),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1453),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1453),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1457),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1472),
.B(n_1447),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1478),
.B(n_1464),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1463),
.A2(n_1400),
.B1(n_1366),
.B2(n_1362),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1464),
.A2(n_1463),
.B(n_1452),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1449),
.B(n_1405),
.Y(n_1507)
);

NAND4xp25_ASAP7_75t_L g1508 ( 
.A(n_1478),
.B(n_1427),
.C(n_1425),
.D(n_1415),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1419),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1469),
.B(n_1419),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1463),
.A2(n_1400),
.B1(n_1479),
.B2(n_1452),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1466),
.B(n_1425),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1457),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1427),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1468),
.B(n_1429),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_SL g1516 ( 
.A1(n_1477),
.A2(n_1438),
.B1(n_1442),
.B2(n_1386),
.C(n_1390),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1397),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1468),
.B(n_1429),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1461),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1461),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1468),
.B(n_1438),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1474),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1465),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1484),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1484),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1492),
.B(n_1471),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1485),
.B(n_1455),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1453),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1504),
.B(n_1455),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1490),
.A2(n_1455),
.B1(n_1414),
.B2(n_1460),
.C(n_1476),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1492),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1482),
.B(n_1471),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1482),
.B(n_1456),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1489),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1498),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1496),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1483),
.A2(n_1463),
.B1(n_1452),
.B2(n_1479),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1498),
.B(n_1471),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1499),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1516),
.B(n_1456),
.Y(n_1541)
);

INVx3_ASAP7_75t_SL g1542 ( 
.A(n_1497),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1489),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1491),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1491),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1494),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1509),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1514),
.B(n_1442),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1481),
.B(n_1456),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1481),
.B(n_1460),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1501),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1460),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1506),
.B(n_1445),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1505),
.A2(n_1463),
.B1(n_1455),
.B2(n_1452),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1514),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1500),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1531),
.B(n_1486),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1549),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1524),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1554),
.B(n_1503),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1542),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1515),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1539),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1542),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1552),
.B(n_1508),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1549),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1493),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1536),
.B(n_1510),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1515),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1550),
.B(n_1494),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1525),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1507),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1527),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1535),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1543),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1528),
.B(n_1507),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1538),
.A2(n_1511),
.B1(n_1463),
.B2(n_1488),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1558),
.B(n_1517),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1532),
.B(n_1518),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1549),
.Y(n_1585)
);

OAI21xp33_ASAP7_75t_L g1586 ( 
.A1(n_1560),
.A2(n_1558),
.B(n_1537),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1564),
.B(n_1537),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1580),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1577),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1577),
.A2(n_1530),
.B1(n_1541),
.B2(n_1555),
.C(n_1534),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1570),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1585),
.B(n_1550),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1526),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1580),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1579),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1573),
.B(n_1527),
.C(n_1544),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1574),
.B(n_1545),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1526),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1570),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1568),
.A2(n_1518),
.B(n_1556),
.Y(n_1600)
);

AOI211x1_ASAP7_75t_L g1601 ( 
.A1(n_1572),
.A2(n_1557),
.B(n_1547),
.C(n_1548),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1582),
.A2(n_1555),
.B(n_1559),
.C(n_1533),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1579),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1592),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1591),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1589),
.B(n_1566),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1589),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1563),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1597),
.B(n_1576),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1599),
.B(n_1566),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1598),
.B(n_1581),
.Y(n_1611)
);

OAI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1590),
.A2(n_1556),
.B1(n_1584),
.B2(n_1565),
.C1(n_1452),
.C2(n_1583),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1587),
.B(n_1569),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1609),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1604),
.B(n_1569),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_SL g1616 ( 
.A(n_1606),
.B(n_1596),
.C(n_1600),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1612),
.A2(n_1587),
.B(n_1570),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_R g1618 ( 
.A(n_1613),
.B(n_1588),
.Y(n_1618)
);

OAI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1607),
.A2(n_1601),
.B(n_1586),
.C(n_1569),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1610),
.A2(n_1590),
.B1(n_1602),
.B2(n_1595),
.C(n_1603),
.Y(n_1620)
);

AOI211xp5_ASAP7_75t_L g1621 ( 
.A1(n_1611),
.A2(n_1594),
.B(n_1584),
.C(n_1565),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1608),
.B(n_1571),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1616),
.A2(n_1605),
.B(n_1575),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1622),
.A2(n_1556),
.B1(n_1539),
.B2(n_1547),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1620),
.A2(n_1578),
.B(n_1562),
.C(n_1559),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1614),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1621),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1627),
.B(n_1617),
.Y(n_1628)
);

NAND2xp33_ASAP7_75t_SL g1629 ( 
.A(n_1624),
.B(n_1618),
.Y(n_1629)
);

OAI321xp33_ASAP7_75t_L g1630 ( 
.A1(n_1626),
.A2(n_1619),
.A3(n_1615),
.B1(n_1452),
.B2(n_1546),
.C(n_1533),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1623),
.B(n_1546),
.C(n_1540),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1625),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1626),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_R g1634 ( 
.A(n_1629),
.B(n_1551),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1628),
.B(n_1512),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_R g1636 ( 
.A(n_1633),
.B(n_1551),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1631),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1632),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1635),
.B(n_1540),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1638),
.Y(n_1640)
);

XNOR2xp5_ASAP7_75t_L g1641 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1640),
.B(n_1634),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1641),
.B1(n_1639),
.B2(n_1636),
.C(n_1523),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1643),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1643),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1644),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1645),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1646),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_SL g1649 ( 
.A1(n_1647),
.A2(n_1495),
.B1(n_1403),
.B2(n_1520),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1648),
.A2(n_1649),
.B1(n_1521),
.B2(n_1523),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1502),
.B(n_1520),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1651),
.B(n_1502),
.Y(n_1652)
);

AOI22x1_ASAP7_75t_L g1653 ( 
.A1(n_1652),
.A2(n_1519),
.B1(n_1513),
.B2(n_1521),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1653),
.A2(n_1519),
.B1(n_1513),
.B2(n_1476),
.Y(n_1654)
);

AOI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1403),
.B(n_1360),
.C(n_1462),
.Y(n_1655)
);


endmodule