module real_aes_6931_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_182;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g532 ( .A1(n_0), .A2(n_136), .B(n_533), .C(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_1), .B(n_477), .Y(n_537) );
INVx1_ASAP7_75t_L g421 ( .A(n_2), .Y(n_421) );
INVx1_ASAP7_75t_L g170 ( .A(n_3), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_4), .B(n_128), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_5), .A2(n_446), .B(n_471), .Y(n_470) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_6), .A2(n_113), .B(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_7), .A2(n_35), .B1(n_122), .B2(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_8), .B(n_113), .Y(n_139) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_10), .A2(n_137), .B(n_436), .C(n_438), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_11), .B(n_36), .Y(n_422) );
INVx1_ASAP7_75t_L g163 ( .A(n_12), .Y(n_163) );
INVx1_ASAP7_75t_L g118 ( .A(n_13), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_14), .B(n_126), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_15), .B(n_128), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_16), .B(n_114), .Y(n_175) );
AO32x2_ASAP7_75t_L g197 ( .A1(n_17), .A2(n_113), .A3(n_143), .B1(n_154), .B2(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_18), .B(n_122), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_19), .B(n_114), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_20), .A2(n_52), .B1(n_122), .B2(n_200), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_21), .A2(n_79), .B1(n_122), .B2(n_126), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_22), .B(n_122), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_23), .A2(n_154), .B(n_436), .C(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_24), .A2(n_154), .B(n_436), .C(n_465), .Y(n_464) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_25), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_26), .B(n_156), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_27), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_28), .A2(n_446), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_29), .B(n_156), .Y(n_194) );
INVx2_ASAP7_75t_L g124 ( .A(n_30), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_31), .A2(n_448), .B(n_456), .C(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_32), .B(n_122), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_33), .B(n_156), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_34), .B(n_208), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_37), .B(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_38), .Y(n_442) );
AOI222xp33_ASAP7_75t_SL g101 ( .A1(n_39), .A2(n_77), .B1(n_102), .B2(n_711), .C1(n_712), .C2(n_716), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g711 ( .A(n_39), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_40), .B(n_128), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_41), .B(n_446), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_42), .A2(n_100), .B1(n_720), .B2(n_730), .C1(n_744), .C2(n_750), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_42), .A2(n_76), .B1(n_416), .B2(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_42), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_43), .A2(n_448), .B(n_450), .C(n_456), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_44), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g534 ( .A(n_45), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_46), .A2(n_87), .B1(n_200), .B2(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g451 ( .A(n_47), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_48), .B(n_122), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_49), .B(n_122), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_50), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_51), .B(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_SL g179 ( .A1(n_53), .A2(n_57), .B1(n_122), .B2(n_126), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_54), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_55), .B(n_122), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_56), .B(n_122), .Y(n_205) );
INVx1_ASAP7_75t_L g138 ( .A(n_58), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_59), .B(n_446), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_60), .B(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_61), .A2(n_134), .B(n_166), .C(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_62), .B(n_122), .Y(n_171) );
INVx1_ASAP7_75t_L g117 ( .A(n_63), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_64), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_65), .B(n_128), .Y(n_487) );
AO32x2_ASAP7_75t_L g218 ( .A1(n_66), .A2(n_113), .A3(n_154), .B1(n_219), .B2(n_223), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_67), .B(n_129), .Y(n_439) );
INVx1_ASAP7_75t_L g149 ( .A(n_68), .Y(n_149) );
INVx1_ASAP7_75t_L g189 ( .A(n_69), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_70), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_71), .B(n_453), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_72), .A2(n_436), .B(n_456), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_73), .B(n_126), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_74), .Y(n_472) );
INVx1_ASAP7_75t_L g725 ( .A(n_75), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g104 ( .A1(n_76), .A2(n_105), .B1(n_415), .B2(n_416), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_76), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_78), .B(n_452), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_80), .B(n_200), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_81), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_82), .B(n_126), .Y(n_193) );
INVx2_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_84), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_85), .B(n_153), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_86), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g419 ( .A(n_88), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g710 ( .A(n_88), .Y(n_710) );
OR2x2_ASAP7_75t_L g729 ( .A(n_88), .B(n_719), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_89), .A2(n_98), .B1(n_126), .B2(n_127), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_90), .B(n_446), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_91), .Y(n_486) );
INVxp67_ASAP7_75t_L g475 ( .A(n_92), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_93), .B(n_126), .Y(n_147) );
INVx1_ASAP7_75t_L g432 ( .A(n_94), .Y(n_432) );
INVx1_ASAP7_75t_L g510 ( .A(n_95), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_96), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g458 ( .A(n_97), .B(n_156), .Y(n_458) );
INVxp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g102 ( .A1(n_103), .A2(n_417), .B1(n_423), .B2(n_707), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_104), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
INVx2_ASAP7_75t_L g415 ( .A(n_105), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_105), .A2(n_415), .B1(n_736), .B2(n_737), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g105 ( .A(n_106), .B(n_339), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_297), .Y(n_106) );
NOR4xp25_ASAP7_75t_L g107 ( .A(n_108), .B(n_237), .C(n_273), .D(n_287), .Y(n_107) );
OAI221xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_181), .B1(n_213), .B2(n_224), .C(n_228), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_109), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_157), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_140), .Y(n_111) );
AND2x2_ASAP7_75t_L g234 ( .A(n_112), .B(n_141), .Y(n_234) );
INVx3_ASAP7_75t_L g242 ( .A(n_112), .Y(n_242) );
AND2x2_ASAP7_75t_L g296 ( .A(n_112), .B(n_160), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_112), .B(n_159), .Y(n_332) );
AND2x2_ASAP7_75t_L g390 ( .A(n_112), .B(n_252), .Y(n_390) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_119), .B(n_139), .Y(n_112) );
INVx4_ASAP7_75t_L g180 ( .A(n_113), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_113), .A2(n_463), .B(n_464), .Y(n_462) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_113), .Y(n_469) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g143 ( .A(n_114), .Y(n_143) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_115), .B(n_116), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_131), .B(n_137), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_128), .Y(n_120) );
INVx3_ASAP7_75t_L g188 ( .A(n_122), .Y(n_188) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_122), .Y(n_512) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g200 ( .A(n_123), .Y(n_200) );
BUFx3_ASAP7_75t_L g221 ( .A(n_123), .Y(n_221) );
AND2x6_ASAP7_75t_L g436 ( .A(n_123), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g127 ( .A(n_124), .Y(n_127) );
INVx1_ASAP7_75t_L g135 ( .A(n_124), .Y(n_135) );
INVx2_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_128), .A2(n_146), .B(n_147), .Y(n_145) );
O2A1O1Ixp5_ASAP7_75t_SL g187 ( .A1(n_128), .A2(n_188), .B(n_189), .C(n_190), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_128), .B(n_475), .Y(n_474) );
INVx5_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g219 ( .A1(n_129), .A2(n_153), .B1(n_220), .B2(n_222), .Y(n_219) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_130), .Y(n_153) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
INVx1_ASAP7_75t_L g208 ( .A(n_130), .Y(n_208) );
AND2x2_ASAP7_75t_L g434 ( .A(n_130), .B(n_135), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_130), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_136), .Y(n_131) );
INVx2_ASAP7_75t_L g150 ( .A(n_134), .Y(n_150) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_136), .A2(n_150), .B(n_170), .C(n_171), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_136), .A2(n_153), .B1(n_178), .B2(n_179), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_136), .A2(n_153), .B1(n_199), .B2(n_201), .Y(n_198) );
BUFx3_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_137), .A2(n_162), .B(n_169), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_137), .A2(n_187), .B(n_191), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_137), .A2(n_204), .B(n_209), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_137), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g446 ( .A(n_137), .B(n_434), .Y(n_446) );
INVx4_ASAP7_75t_SL g457 ( .A(n_137), .Y(n_457) );
AND2x2_ASAP7_75t_L g225 ( .A(n_140), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g239 ( .A(n_140), .B(n_160), .Y(n_239) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_141), .B(n_160), .Y(n_254) );
AND2x2_ASAP7_75t_L g266 ( .A(n_141), .B(n_242), .Y(n_266) );
OR2x2_ASAP7_75t_L g268 ( .A(n_141), .B(n_226), .Y(n_268) );
AND2x2_ASAP7_75t_L g303 ( .A(n_141), .B(n_226), .Y(n_303) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_141), .Y(n_348) );
INVx1_ASAP7_75t_L g356 ( .A(n_141), .Y(n_356) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B(n_155), .Y(n_141) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_142), .A2(n_161), .B(n_172), .Y(n_160) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_143), .B(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_154), .Y(n_144) );
O2A1O1Ixp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_151), .C(n_152), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_150), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_152), .A2(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g535 ( .A(n_153), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g176 ( .A(n_154), .B(n_177), .C(n_180), .Y(n_176) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_156), .A2(n_186), .B(n_194), .Y(n_185) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_203), .B(n_212), .Y(n_202) );
INVx2_ASAP7_75t_L g223 ( .A(n_156), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_156), .A2(n_445), .B(n_447), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_156), .A2(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g503 ( .A(n_156), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g273 ( .A1(n_157), .A2(n_274), .B1(n_278), .B2(n_282), .C(n_283), .Y(n_273) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g233 ( .A(n_158), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_173), .Y(n_158) );
INVx2_ASAP7_75t_L g232 ( .A(n_159), .Y(n_232) );
AND2x2_ASAP7_75t_L g285 ( .A(n_159), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g304 ( .A(n_159), .B(n_242), .Y(n_304) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g367 ( .A(n_160), .B(n_242), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .C(n_166), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_164), .A2(n_439), .B(n_440), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_164), .A2(n_466), .B(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_166), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_167), .A2(n_192), .B(n_193), .Y(n_191) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g453 ( .A(n_168), .Y(n_453) );
AND2x2_ASAP7_75t_L g289 ( .A(n_173), .B(n_234), .Y(n_289) );
OAI322xp33_ASAP7_75t_L g357 ( .A1(n_173), .A2(n_313), .A3(n_358), .B1(n_360), .B2(n_363), .C1(n_365), .C2(n_369), .Y(n_357) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_174), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g253 ( .A(n_174), .Y(n_253) );
AND2x2_ASAP7_75t_L g362 ( .A(n_174), .B(n_242), .Y(n_362) );
AND2x2_ASAP7_75t_L g394 ( .A(n_174), .B(n_266), .Y(n_394) );
OR2x2_ASAP7_75t_L g397 ( .A(n_174), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
AO21x1_ASAP7_75t_L g226 ( .A1(n_177), .A2(n_180), .B(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_180), .A2(n_431), .B(n_441), .Y(n_430) );
INVx3_ASAP7_75t_L g477 ( .A(n_180), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_180), .B(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_180), .A2(n_507), .B(n_514), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_180), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_195), .Y(n_182) );
INVx1_ASAP7_75t_L g410 ( .A(n_183), .Y(n_410) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g215 ( .A(n_184), .B(n_202), .Y(n_215) );
INVx2_ASAP7_75t_L g250 ( .A(n_184), .Y(n_250) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_185), .Y(n_280) );
OR2x2_ASAP7_75t_L g404 ( .A(n_185), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g229 ( .A(n_195), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g269 ( .A(n_195), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g321 ( .A(n_195), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_202), .Y(n_195) );
AND2x2_ASAP7_75t_L g216 ( .A(n_196), .B(n_217), .Y(n_216) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_196), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g330 ( .A(n_196), .B(n_218), .Y(n_330) );
OR2x2_ASAP7_75t_L g338 ( .A(n_196), .B(n_272), .Y(n_338) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g247 ( .A(n_197), .Y(n_247) );
AND2x2_ASAP7_75t_L g257 ( .A(n_197), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g281 ( .A(n_197), .B(n_202), .Y(n_281) );
AND2x2_ASAP7_75t_L g345 ( .A(n_197), .B(n_218), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_202), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_202), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g258 ( .A(n_202), .Y(n_258) );
INVx1_ASAP7_75t_L g263 ( .A(n_202), .Y(n_263) );
AND2x2_ASAP7_75t_L g275 ( .A(n_202), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_202), .Y(n_353) );
INVx1_ASAP7_75t_L g405 ( .A(n_202), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
AND2x2_ASAP7_75t_L g382 ( .A(n_214), .B(n_291), .Y(n_382) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g309 ( .A(n_216), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g408 ( .A(n_216), .B(n_343), .Y(n_408) );
INVx1_ASAP7_75t_L g230 ( .A(n_217), .Y(n_230) );
AND2x2_ASAP7_75t_L g256 ( .A(n_217), .B(n_250), .Y(n_256) );
BUFx2_ASAP7_75t_L g315 ( .A(n_217), .Y(n_315) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_218), .Y(n_236) );
INVx1_ASAP7_75t_L g246 ( .A(n_218), .Y(n_246) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_221), .Y(n_455) );
INVx2_ASAP7_75t_L g536 ( .A(n_221), .Y(n_536) );
INVx1_ASAP7_75t_L g500 ( .A(n_223), .Y(n_500) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_224), .B(n_231), .Y(n_384) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI32xp33_ASAP7_75t_L g228 ( .A1(n_225), .A2(n_229), .A3(n_231), .B1(n_233), .B2(n_235), .Y(n_228) );
AND2x2_ASAP7_75t_L g368 ( .A(n_225), .B(n_241), .Y(n_368) );
AND2x2_ASAP7_75t_L g406 ( .A(n_225), .B(n_304), .Y(n_406) );
INVx1_ASAP7_75t_L g286 ( .A(n_226), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_230), .B(n_292), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_231), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_231), .B(n_234), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_231), .B(n_303), .Y(n_385) );
OR2x2_ASAP7_75t_L g399 ( .A(n_231), .B(n_268), .Y(n_399) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_234), .Y(n_326) );
OR2x2_ASAP7_75t_L g335 ( .A(n_232), .B(n_322), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_234), .B(n_285), .Y(n_307) );
INVx2_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
OR2x2_ASAP7_75t_L g337 ( .A(n_236), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g352 ( .A(n_236), .B(n_353), .Y(n_352) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_236), .A2(n_329), .B(n_410), .C(n_411), .Y(n_409) );
OAI321xp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_243), .A3(n_248), .B1(n_251), .B2(n_255), .C(n_259), .Y(n_237) );
INVx1_ASAP7_75t_L g350 ( .A(n_238), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g361 ( .A(n_239), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g313 ( .A(n_241), .Y(n_313) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_242), .B(n_356), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_243), .A2(n_381), .B1(n_383), .B2(n_385), .C(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
AND2x2_ASAP7_75t_L g318 ( .A(n_245), .B(n_292), .Y(n_318) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_246), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g291 ( .A(n_247), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_248), .A2(n_289), .B(n_334), .C(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g300 ( .A(n_250), .B(n_257), .Y(n_300) );
BUFx2_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
INVx1_ASAP7_75t_L g325 ( .A(n_250), .Y(n_325) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OR2x2_ASAP7_75t_L g331 ( .A(n_253), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g414 ( .A(n_253), .Y(n_414) );
INVx1_ASAP7_75t_L g407 ( .A(n_254), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g260 ( .A(n_256), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g364 ( .A(n_256), .B(n_281), .Y(n_364) );
INVx1_ASAP7_75t_L g293 ( .A(n_257), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_264), .B1(n_267), .B2(n_269), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_261), .B(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g329 ( .A(n_262), .B(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_SL g292 ( .A(n_263), .B(n_272), .Y(n_292) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g284 ( .A(n_266), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g294 ( .A(n_268), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_271), .A2(n_389), .B1(n_391), .B2(n_392), .C(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g277 ( .A(n_272), .Y(n_277) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_272), .Y(n_343) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_275), .B(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_276), .A2(n_281), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_279), .B(n_289), .Y(n_386) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g355 ( .A(n_280), .Y(n_355) );
AND2x2_ASAP7_75t_L g314 ( .A(n_281), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g403 ( .A(n_281), .Y(n_403) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
INVx1_ASAP7_75t_L g374 ( .A(n_285), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B1(n_293), .B2(n_294), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_291), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g359 ( .A(n_292), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_292), .B(n_330), .Y(n_396) );
OR2x2_ASAP7_75t_L g369 ( .A(n_293), .B(n_322), .Y(n_369) );
INVx1_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_296), .B(n_347), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_316), .C(n_327), .Y(n_297) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_305), .C(n_311), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_300), .A2(n_371), .B1(n_375), .B2(n_378), .C(n_380), .Y(n_370) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g312 ( .A(n_303), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g366 ( .A(n_303), .B(n_367), .Y(n_366) );
OAI211xp5_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_352), .B(n_354), .C(n_356), .Y(n_351) );
INVx2_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
OAI21xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_308), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g377 ( .A(n_310), .B(n_330), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
OAI21xp5_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_319), .B(n_320), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_323), .B(n_326), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_321), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_326), .B(n_413), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B(n_333), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g354 ( .A(n_330), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND4x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_370), .C(n_387), .D(n_409), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_357), .Y(n_340) );
OAI211xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_346), .B(n_349), .C(n_351), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_345), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_356), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g391 ( .A(n_366), .Y(n_391) );
INVx2_ASAP7_75t_SL g379 ( .A(n_367), .Y(n_379) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g392 ( .A(n_377), .Y(n_392) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_SL g387 ( .A(n_388), .B(n_395), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
OAI221xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B1(n_399), .B2(n_400), .C(n_401), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g713 ( .A(n_418), .Y(n_713) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g709 ( .A(n_420), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g719 ( .A(n_420), .Y(n_719) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_L g714 ( .A(n_423), .Y(n_714) );
OR3x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_605), .C(n_670), .Y(n_423) );
NAND4xp25_ASAP7_75t_SL g424 ( .A(n_425), .B(n_546), .C(n_572), .D(n_595), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_478), .B1(n_516), .B2(n_523), .C(n_538), .Y(n_425) );
CKINVDCx14_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_427), .A2(n_539), .B1(n_563), .B2(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_459), .Y(n_427) );
INVx1_ASAP7_75t_SL g599 ( .A(n_428), .Y(n_599) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_443), .Y(n_428) );
OR2x2_ASAP7_75t_L g521 ( .A(n_429), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g541 ( .A(n_429), .B(n_460), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_429), .B(n_468), .Y(n_554) );
AND2x2_ASAP7_75t_L g571 ( .A(n_429), .B(n_443), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_429), .B(n_519), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_429), .B(n_570), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_429), .B(n_459), .Y(n_692) );
AOI211xp5_ASAP7_75t_SL g703 ( .A1(n_429), .A2(n_609), .B(n_704), .C(n_705), .Y(n_703) );
INVx5_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_430), .B(n_460), .Y(n_575) );
AND2x2_ASAP7_75t_L g578 ( .A(n_430), .B(n_461), .Y(n_578) );
OR2x2_ASAP7_75t_L g623 ( .A(n_430), .B(n_460), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_430), .B(n_468), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_435), .Y(n_431) );
INVx5_ASAP7_75t_L g449 ( .A(n_436), .Y(n_449) );
INVx5_ASAP7_75t_SL g522 ( .A(n_443), .Y(n_522) );
AND2x2_ASAP7_75t_L g540 ( .A(n_443), .B(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_443), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g626 ( .A(n_443), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g658 ( .A(n_443), .B(n_468), .Y(n_658) );
OR2x2_ASAP7_75t_L g664 ( .A(n_443), .B(n_554), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_443), .B(n_614), .Y(n_673) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_458), .Y(n_443) );
BUFx2_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_449), .A2(n_457), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_449), .A2(n_457), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_454), .C(n_455), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_452), .A2(n_455), .B(n_486), .C(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_468), .Y(n_459) );
AND2x2_ASAP7_75t_L g555 ( .A(n_460), .B(n_522), .Y(n_555) );
INVx1_ASAP7_75t_SL g568 ( .A(n_460), .Y(n_568) );
OR2x2_ASAP7_75t_L g603 ( .A(n_460), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g609 ( .A(n_460), .B(n_468), .Y(n_609) );
AND2x2_ASAP7_75t_L g667 ( .A(n_460), .B(n_519), .Y(n_667) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_461), .B(n_522), .Y(n_594) );
INVx3_ASAP7_75t_L g519 ( .A(n_468), .Y(n_519) );
OR2x2_ASAP7_75t_L g560 ( .A(n_468), .B(n_522), .Y(n_560) );
AND2x2_ASAP7_75t_L g570 ( .A(n_468), .B(n_568), .Y(n_570) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_468), .Y(n_618) );
AND2x2_ASAP7_75t_L g627 ( .A(n_468), .B(n_541), .Y(n_627) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_476), .Y(n_468) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_477), .A2(n_529), .B(n_537), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_478), .A2(n_644), .B1(n_646), .B2(n_648), .C(n_651), .Y(n_643) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_490), .Y(n_479) );
AND2x2_ASAP7_75t_L g617 ( .A(n_480), .B(n_598), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_480), .B(n_676), .Y(n_680) );
OR2x2_ASAP7_75t_L g701 ( .A(n_480), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_480), .B(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx5_ASAP7_75t_L g548 ( .A(n_481), .Y(n_548) );
AND2x2_ASAP7_75t_L g625 ( .A(n_481), .B(n_492), .Y(n_625) );
AND2x2_ASAP7_75t_L g686 ( .A(n_481), .B(n_565), .Y(n_686) );
AND2x2_ASAP7_75t_L g699 ( .A(n_481), .B(n_519), .Y(n_699) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_488), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_504), .Y(n_490) );
AND2x4_ASAP7_75t_L g526 ( .A(n_491), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g544 ( .A(n_491), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
AND2x2_ASAP7_75t_L g620 ( .A(n_491), .B(n_598), .Y(n_620) );
AND2x2_ASAP7_75t_L g630 ( .A(n_491), .B(n_548), .Y(n_630) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_491), .Y(n_638) );
AND2x2_ASAP7_75t_L g650 ( .A(n_491), .B(n_528), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_491), .B(n_582), .Y(n_654) );
AND2x2_ASAP7_75t_L g691 ( .A(n_491), .B(n_686), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_491), .B(n_565), .Y(n_702) );
OR2x2_ASAP7_75t_L g704 ( .A(n_491), .B(n_640), .Y(n_704) );
INVx5_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g590 ( .A(n_492), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g600 ( .A(n_492), .B(n_545), .Y(n_600) );
AND2x2_ASAP7_75t_L g612 ( .A(n_492), .B(n_528), .Y(n_612) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_492), .Y(n_642) );
AND2x4_ASAP7_75t_L g676 ( .A(n_492), .B(n_527), .Y(n_676) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
AOI21xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B(n_500), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
BUFx2_ASAP7_75t_L g525 ( .A(n_504), .Y(n_525) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
AND2x2_ASAP7_75t_L g598 ( .A(n_505), .B(n_528), .Y(n_598) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g545 ( .A(n_506), .B(n_528), .Y(n_545) );
BUFx2_ASAP7_75t_L g591 ( .A(n_506), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_518), .B(n_599), .Y(n_678) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_519), .B(n_541), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_519), .B(n_522), .Y(n_580) );
AND2x2_ASAP7_75t_L g635 ( .A(n_519), .B(n_571), .Y(n_635) );
AOI221xp5_ASAP7_75t_SL g572 ( .A1(n_520), .A2(n_573), .B1(n_581), .B2(n_583), .C(n_587), .Y(n_572) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g567 ( .A(n_521), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g608 ( .A(n_521), .B(n_609), .Y(n_608) );
OAI321xp33_ASAP7_75t_L g615 ( .A1(n_521), .A2(n_574), .A3(n_616), .B1(n_618), .B2(n_619), .C(n_621), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_522), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_525), .B(n_676), .Y(n_694) );
AND2x2_ASAP7_75t_L g581 ( .A(n_526), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_526), .B(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_527), .Y(n_557) );
AND2x2_ASAP7_75t_L g564 ( .A(n_527), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_527), .B(n_639), .Y(n_669) );
INVx1_ASAP7_75t_L g706 ( .A(n_527), .Y(n_706) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_542), .B(n_543), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_540), .A2(n_650), .B(n_699), .C(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_541), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_541), .B(n_579), .Y(n_645) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g588 ( .A(n_545), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_545), .B(n_548), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_545), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_545), .B(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_549), .B1(n_561), .B2(n_566), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g562 ( .A(n_548), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g585 ( .A(n_548), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g597 ( .A(n_548), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_548), .B(n_591), .Y(n_633) );
OR2x2_ASAP7_75t_L g640 ( .A(n_548), .B(n_565), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_548), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g690 ( .A(n_548), .B(n_676), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_552), .B1(n_556), .B2(n_558), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g596 ( .A(n_551), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_554), .A2(n_569), .B1(n_637), .B2(n_641), .Y(n_636) );
INVx1_ASAP7_75t_L g684 ( .A(n_555), .Y(n_684) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_559), .A2(n_596), .B1(n_599), .B2(n_600), .C(n_601), .Y(n_595) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g574 ( .A(n_560), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_564), .B(n_630), .Y(n_662) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_565), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_565), .Y(n_586) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
AND2x2_ASAP7_75t_L g613 ( .A(n_571), .B(n_614), .Y(n_613) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx2_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x2_ASAP7_75t_L g657 ( .A(n_578), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_581), .A2(n_607), .B1(n_610), .B2(n_613), .C(n_615), .Y(n_606) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_585), .B(n_642), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B(n_592), .Y(n_587) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
CKINVDCx16_ASAP7_75t_R g689 ( .A(n_592), .Y(n_689) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g631 ( .A(n_594), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g652 ( .A(n_597), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_597), .B(n_657), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_600), .B(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_606), .B(n_624), .C(n_643), .D(n_656), .Y(n_605) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g614 ( .A(n_609), .Y(n_614) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g647 ( .A(n_618), .B(n_623), .Y(n_647) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI211xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_628), .C(n_636), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_626), .A2(n_668), .B(n_696), .C(n_703), .Y(n_695) );
INVx1_ASAP7_75t_SL g655 ( .A(n_627), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_628) );
INVx1_ASAP7_75t_L g659 ( .A(n_633), .Y(n_659) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_639), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_639), .B(n_650), .Y(n_683) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g660 ( .A(n_650), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_655), .Y(n_651) );
INVxp33_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .A3(n_660), .B1(n_661), .B2(n_663), .C1(n_665), .C2(n_668), .Y(n_656) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND3xp33_ASAP7_75t_SL g670 ( .A(n_671), .B(n_688), .C(n_695), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_677), .B2(n_679), .C(n_681), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g687 ( .A(n_676), .Y(n_687) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_688) );
NAND2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g715 ( .A(n_708), .Y(n_715) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_710), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .Y(n_722) );
NOR2xp33_ASAP7_75t_SL g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_SL g749 ( .A(n_724), .Y(n_749) );
INVx1_ASAP7_75t_L g748 ( .A(n_726), .Y(n_748) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_726), .A2(n_749), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g740 ( .A(n_729), .Y(n_740) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_729), .Y(n_742) );
BUFx2_ASAP7_75t_L g752 ( .A(n_729), .Y(n_752) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_739), .B(n_741), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_SL g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
CKINVDCx6p67_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
endmodule