module fake_aes_4564_n_485 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_485);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_485;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_73;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_393;
wire n_135;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g67 ( .A(n_23), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_6), .Y(n_68) );
INVx2_ASAP7_75t_L g69 ( .A(n_5), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_44), .Y(n_70) );
BUFx6f_ASAP7_75t_L g71 ( .A(n_38), .Y(n_71) );
INVxp67_ASAP7_75t_SL g72 ( .A(n_66), .Y(n_72) );
INVxp67_ASAP7_75t_L g73 ( .A(n_17), .Y(n_73) );
INVxp67_ASAP7_75t_SL g74 ( .A(n_1), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_17), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_40), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_42), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_20), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_26), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_61), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_16), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_24), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_9), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_59), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_8), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_28), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_30), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_13), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_35), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_1), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_32), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_50), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_22), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_7), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
CKINVDCx14_ASAP7_75t_R g97 ( .A(n_36), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_13), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_3), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_78), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
INVx3_ASAP7_75t_L g105 ( .A(n_69), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_68), .B(n_0), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_67), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_81), .Y(n_111) );
INVx5_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_81), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_93), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_70), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_84), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_68), .B(n_0), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_84), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
BUFx10_ASAP7_75t_L g126 ( .A(n_107), .Y(n_126) );
INVx2_ASAP7_75t_SL g127 ( .A(n_108), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_108), .B(n_80), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_117), .B(n_85), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_115), .B(n_98), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_115), .B(n_98), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_117), .B(n_97), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_119), .B(n_73), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_102), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_109), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_107), .B(n_89), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_107), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_111), .B(n_87), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_109), .Y(n_143) );
BUFx4f_ASAP7_75t_L g144 ( .A(n_123), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_112), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_121), .B(n_73), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_113), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_112), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_132), .B(n_123), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_148), .B(n_121), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_148), .B(n_125), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_144), .A2(n_124), .B1(n_118), .B2(n_110), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_132), .B(n_125), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_130), .Y(n_158) );
OR2x2_ASAP7_75t_SL g159 ( .A(n_128), .B(n_75), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_127), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_144), .B(n_123), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_141), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_131), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_141), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_133), .B(n_123), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_142), .B(n_88), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_128), .B(n_122), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
NOR2xp33_ASAP7_75t_R g173 ( .A(n_126), .B(n_100), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
NOR3xp33_ASAP7_75t_SL g175 ( .A(n_129), .B(n_95), .C(n_86), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_149), .A2(n_91), .B1(n_74), .B2(n_86), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
NOR2xp33_ASAP7_75t_R g179 ( .A(n_126), .B(n_79), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_126), .B(n_72), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_129), .B(n_122), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_149), .B(n_105), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_139), .B(n_89), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_139), .B(n_96), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g185 ( .A(n_136), .B(n_72), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_134), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_169), .B(n_127), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_181), .B(n_136), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_174), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_167), .A2(n_136), .B1(n_134), .B2(n_150), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_167), .A2(n_152), .B1(n_137), .B2(n_150), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_158), .B(n_96), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_182), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
AOI222xp33_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_99), .B1(n_106), .B2(n_104), .C1(n_105), .C2(n_143), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_187), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_177), .B(n_137), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_154), .A2(n_152), .B(n_147), .C(n_138), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_167), .B(n_138), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_164), .B(n_99), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
OR2x6_ASAP7_75t_L g208 ( .A(n_183), .B(n_90), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_153), .B(n_76), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_172), .A2(n_147), .B1(n_143), .B2(n_76), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_160), .A2(n_178), .B(n_161), .Y(n_211) );
INVxp67_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
INVx3_ASAP7_75t_SL g213 ( .A(n_164), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_153), .A2(n_120), .B(n_114), .C(n_116), .Y(n_214) );
INVxp67_ASAP7_75t_SL g215 ( .A(n_162), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_156), .Y(n_216) );
INVx3_ASAP7_75t_SL g217 ( .A(n_162), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_168), .B(n_92), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_191), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_202), .Y(n_223) );
NOR2xp33_ASAP7_75t_R g224 ( .A(n_213), .B(n_180), .Y(n_224) );
CKINVDCx6p67_ASAP7_75t_R g225 ( .A(n_213), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_200), .B(n_153), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_191), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_192), .A2(n_186), .B1(n_183), .B2(n_184), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_201), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_202), .Y(n_230) );
INVx4_ASAP7_75t_SL g231 ( .A(n_217), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_208), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g233 ( .A1(n_216), .A2(n_185), .B1(n_179), .B2(n_183), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_212), .B(n_184), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_196), .B(n_184), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_202), .Y(n_236) );
OAI211xp5_ASAP7_75t_SL g237 ( .A1(n_199), .A2(n_175), .B(n_176), .C(n_106), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_216), .A2(n_159), .B1(n_165), .B2(n_162), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_209), .A2(n_165), .B1(n_171), .B2(n_163), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_190), .Y(n_241) );
OAI22xp33_ASAP7_75t_L g242 ( .A1(n_208), .A2(n_165), .B1(n_159), .B2(n_177), .Y(n_242) );
AND2x6_ASAP7_75t_L g243 ( .A(n_191), .B(n_165), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_201), .B(n_177), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_198), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_217), .Y(n_246) );
NOR2x1_ASAP7_75t_SL g247 ( .A(n_208), .B(n_165), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_191), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_229), .B(n_208), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_229), .B(n_209), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_248), .A2(n_211), .B(n_203), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_239), .A2(n_195), .B1(n_206), .B2(n_209), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_226), .B(n_194), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_226), .B(n_188), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_245), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_233), .B(n_214), .C(n_220), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_223), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_243), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_244), .A2(n_189), .B(n_218), .C(n_197), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_237), .A2(n_218), .B1(n_197), .B2(n_210), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_242), .A2(n_232), .B1(n_234), .B2(n_224), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_234), .B(n_205), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_225), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_231), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_232), .A2(n_193), .B1(n_219), .B2(n_204), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g267 ( .A1(n_247), .A2(n_92), .B1(n_105), .B2(n_204), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_230), .A2(n_198), .B1(n_207), .B2(n_120), .Y(n_268) );
NAND2x1_ASAP7_75t_L g269 ( .A(n_243), .B(n_204), .Y(n_269) );
AND2x4_ASAP7_75t_SL g270 ( .A(n_223), .B(n_221), .Y(n_270) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_256), .A2(n_235), .B(n_230), .C(n_246), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_244), .B1(n_228), .B2(n_236), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_254), .B(n_225), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_258), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_262), .A2(n_104), .B1(n_105), .B2(n_241), .C(n_116), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_264), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_255), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_255), .B(n_245), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_253), .A2(n_236), .B1(n_223), .B2(n_246), .Y(n_280) );
AOI33xp33_ASAP7_75t_L g281 ( .A1(n_261), .A2(n_90), .A3(n_94), .B1(n_101), .B2(n_240), .B3(n_219), .Y(n_281) );
OAI21xp33_ASAP7_75t_SL g282 ( .A1(n_249), .A2(n_223), .B(n_236), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_249), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_265), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_263), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_256), .A2(n_244), .B1(n_236), .B2(n_246), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_251), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_262), .B(n_244), .Y(n_288) );
OAI33xp33_ASAP7_75t_L g289 ( .A1(n_250), .A2(n_94), .A3(n_101), .B1(n_207), .B2(n_6), .B3(n_7), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_268), .Y(n_290) );
OAI221xp5_ASAP7_75t_L g291 ( .A1(n_260), .A2(n_82), .B1(n_221), .B2(n_215), .C(n_178), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_251), .A2(n_248), .B(n_247), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_251), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_283), .B(n_257), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
AND4x1_ASAP7_75t_L g296 ( .A(n_281), .B(n_259), .C(n_266), .D(n_231), .Y(n_296) );
AND2x2_ASAP7_75t_SL g297 ( .A(n_276), .B(n_265), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_257), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_287), .Y(n_301) );
OAI33xp33_ASAP7_75t_L g302 ( .A1(n_280), .A2(n_250), .A3(n_268), .B1(n_253), .B2(n_8), .B3(n_9), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_270), .Y(n_304) );
OAI33xp33_ASAP7_75t_L g305 ( .A1(n_280), .A2(n_2), .A3(n_4), .B1(n_5), .B2(n_10), .B3(n_11), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_276), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_293), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_278), .B(n_269), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_271), .B(n_254), .Y(n_311) );
AOI21xp33_ASAP7_75t_L g312 ( .A1(n_271), .A2(n_269), .B(n_267), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_278), .B(n_270), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_292), .B(n_258), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_284), .B(n_270), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_284), .B(n_258), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_284), .B(n_267), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_290), .B(n_248), .Y(n_319) );
AOI22x1_ASAP7_75t_L g320 ( .A1(n_274), .A2(n_290), .B1(n_231), .B2(n_293), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_292), .B(n_71), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_286), .B(n_243), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
NOR2xp33_ASAP7_75t_R g325 ( .A(n_297), .B(n_273), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_300), .B(n_275), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_322), .B(n_292), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_300), .B(n_288), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_295), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_314), .B(n_292), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_297), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_298), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_303), .B(n_275), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_303), .B(n_281), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_297), .B(n_282), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_310), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
OAI211xp5_ASAP7_75t_L g340 ( .A1(n_311), .A2(n_282), .B(n_273), .C(n_286), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_307), .B(n_288), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_310), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_299), .B(n_274), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_311), .A2(n_272), .B1(n_289), .B2(n_291), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_296), .B(n_289), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_314), .B(n_274), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_304), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_294), .B(n_272), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_294), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_296), .B(n_291), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_319), .B(n_2), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_302), .A2(n_231), .B1(n_285), .B2(n_243), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_319), .B(n_4), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_304), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_312), .A2(n_227), .B(n_222), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_314), .B(n_71), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_313), .B(n_10), .Y(n_359) );
NAND3x1_ASAP7_75t_L g360 ( .A(n_313), .B(n_238), .C(n_12), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_318), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_306), .B(n_103), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_306), .B(n_103), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_318), .Y(n_364) );
OA21x2_ASAP7_75t_L g365 ( .A1(n_337), .A2(n_320), .B(n_309), .Y(n_365) );
NOR3xp33_ASAP7_75t_SL g366 ( .A(n_340), .B(n_305), .C(n_312), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_348), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
OAI22xp33_ASAP7_75t_SL g370 ( .A1(n_337), .A2(n_321), .B1(n_315), .B2(n_320), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g371 ( .A1(n_332), .A2(n_316), .B(n_317), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_338), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_333), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_361), .A2(n_305), .B1(n_103), .B2(n_324), .C(n_323), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_341), .B(n_321), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_359), .B(n_11), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_355), .B(n_321), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_364), .B(n_315), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_315), .B1(n_323), .B2(n_309), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_343), .B(n_315), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_360), .A2(n_309), .B1(n_308), .B2(n_238), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_351), .A2(n_308), .B1(n_238), .B2(n_227), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_308), .B1(n_243), .B2(n_238), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_103), .B1(n_112), .B2(n_146), .C(n_16), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_350), .B(n_12), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_343), .B(n_14), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_345), .A2(n_227), .B1(n_222), .B2(n_112), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_357), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_329), .B(n_14), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_356), .A2(n_227), .B(n_222), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_352), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_325), .A2(n_243), .B1(n_227), .B2(n_222), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_349), .B(n_15), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_353), .A2(n_227), .B1(n_222), .B2(n_243), .Y(n_398) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_354), .B(n_222), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_325), .Y(n_400) );
AOI32xp33_ASAP7_75t_L g401 ( .A1(n_328), .A2(n_331), .A3(n_346), .B1(n_335), .B2(n_326), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_344), .B(n_18), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_336), .B(n_18), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_362), .B(n_146), .C(n_160), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_400), .A2(n_331), .B1(n_328), .B2(n_363), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_393), .B(n_363), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_401), .B(n_362), .C(n_358), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_358), .B(n_347), .Y(n_408) );
XNOR2x1_ASAP7_75t_L g409 ( .A(n_367), .B(n_19), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_395), .B(n_21), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_402), .B(n_25), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_372), .B(n_27), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_368), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_369), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_373), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_389), .Y(n_417) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_365), .B(n_146), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_382), .B(n_31), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_388), .Y(n_421) );
NOR2x1_ASAP7_75t_SL g422 ( .A(n_371), .B(n_33), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_379), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g424 ( .A(n_400), .B(n_34), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_375), .Y(n_425) );
INVxp33_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_370), .A2(n_171), .B(n_151), .Y(n_427) );
NAND2xp33_ASAP7_75t_SL g428 ( .A(n_380), .B(n_37), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_397), .B(n_39), .Y(n_429) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_404), .B(n_41), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_404), .B(n_43), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_407), .A2(n_377), .B1(n_403), .B2(n_392), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_417), .B(n_383), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_428), .A2(n_386), .B1(n_370), .B2(n_374), .Y(n_436) );
XNOR2x1_ASAP7_75t_L g437 ( .A(n_409), .B(n_387), .Y(n_437) );
XNOR2xp5_ASAP7_75t_L g438 ( .A(n_424), .B(n_385), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_414), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_417), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g441 ( .A1(n_405), .A2(n_396), .B(n_398), .C(n_390), .Y(n_441) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_430), .B(n_384), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_410), .B(n_394), .Y(n_443) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_426), .B(n_45), .Y(n_444) );
AOI322xp5_ASAP7_75t_L g445 ( .A1(n_421), .A2(n_171), .A3(n_47), .B1(n_48), .B2(n_49), .C1(n_53), .C2(n_54), .Y(n_445) );
XOR2x2_ASAP7_75t_L g446 ( .A(n_422), .B(n_46), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_432), .A2(n_55), .B(n_56), .C(n_57), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_408), .A2(n_146), .B1(n_60), .B2(n_62), .C(n_63), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_415), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_425), .A2(n_146), .B1(n_64), .B2(n_65), .Y(n_452) );
OAI21xp33_ASAP7_75t_SL g453 ( .A1(n_433), .A2(n_58), .B(n_135), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_423), .B(n_135), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_412), .B(n_140), .C(n_145), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_443), .B(n_431), .Y(n_457) );
INVx4_ASAP7_75t_L g458 ( .A(n_446), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_440), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_442), .B(n_418), .Y(n_460) );
NOR2xp33_ASAP7_75t_R g461 ( .A(n_444), .B(n_420), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_453), .B(n_412), .C(n_411), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_436), .B(n_413), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_435), .A2(n_426), .B(n_429), .C(n_427), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_448), .Y(n_465) );
OAI211xp5_ASAP7_75t_SL g466 ( .A1(n_445), .A2(n_145), .B(n_441), .C(n_449), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_456), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_437), .A2(n_438), .B1(n_439), .B2(n_450), .Y(n_468) );
OAI311xp33_ASAP7_75t_L g469 ( .A1(n_454), .A2(n_447), .A3(n_451), .B1(n_455), .C1(n_452), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_434), .A2(n_436), .B(n_453), .C(n_401), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_440), .A2(n_367), .B1(n_400), .B2(n_348), .Y(n_471) );
OAI211xp5_ASAP7_75t_SL g472 ( .A1(n_434), .A2(n_436), .B(n_453), .C(n_401), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_457), .B(n_459), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_460), .B(n_458), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_472), .B(n_470), .C(n_468), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_465), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_458), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_476), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_475), .A2(n_463), .B1(n_466), .B2(n_462), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_473), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_478), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_479), .A2(n_474), .B(n_477), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_481), .Y(n_483) );
AOI22xp5_ASAP7_75t_SL g484 ( .A1(n_483), .A2(n_482), .B1(n_480), .B2(n_467), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_484), .A2(n_469), .B1(n_471), .B2(n_464), .C(n_461), .Y(n_485) );
endmodule