module real_aes_7497_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1106;
wire n_800;
wire n_778;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_1067;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_1034;
wire n_694;
wire n_491;
wire n_549;
wire n_923;
wire n_894;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_994;
wire n_892;
wire n_495;
wire n_1072;
wire n_528;
wire n_1078;
wire n_744;
wire n_384;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_875;
wire n_951;
wire n_467;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_872;
wire n_636;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_1025;
wire n_755;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_973;
wire n_960;
wire n_455;
wire n_671;
wire n_1084;
wire n_725;
wire n_1081;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_1006;
wire n_754;
wire n_417;
wire n_449;
wire n_607;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_713;
wire n_728;
wire n_735;
wire n_598;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1014;
wire n_1003;
wire n_1000;
wire n_727;
wire n_1083;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_1136;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_679;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_1045;
wire n_566;
wire n_967;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g1045 ( .A(n_0), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_1), .A2(n_287), .B1(n_610), .B2(n_745), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_2), .A2(n_154), .B1(n_518), .B2(n_521), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_3), .A2(n_160), .B1(n_468), .B2(n_597), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_4), .Y(n_604) );
INVx1_ASAP7_75t_L g937 ( .A(n_5), .Y(n_937) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_6), .A2(n_349), .B1(n_571), .B2(n_668), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g1130 ( .A(n_7), .Y(n_1130) );
OA22x2_ASAP7_75t_L g1131 ( .A1(n_7), .A2(n_1130), .B1(n_1132), .B2(n_1148), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_8), .A2(n_126), .B1(n_521), .B2(n_770), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_9), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_10), .A2(n_97), .B1(n_520), .B2(n_682), .Y(n_1073) );
AO22x2_ASAP7_75t_L g404 ( .A1(n_11), .A2(n_218), .B1(n_405), .B2(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g1097 ( .A(n_11), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_12), .A2(n_144), .B1(n_503), .B2(n_567), .Y(n_764) );
AOI222xp33_ASAP7_75t_L g874 ( .A1(n_13), .A2(n_325), .B1(n_335), .B2(n_733), .C1(n_875), .C2(n_876), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_14), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_15), .A2(n_211), .B1(n_520), .B2(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g721 ( .A(n_16), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_17), .A2(n_49), .B1(n_756), .B2(n_951), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_18), .A2(n_191), .B1(n_500), .B2(n_828), .C(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g701 ( .A(n_19), .Y(n_701) );
INVx1_ASAP7_75t_L g709 ( .A(n_20), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_21), .A2(n_240), .B1(n_575), .B2(n_576), .Y(n_1058) );
INVx1_ASAP7_75t_L g1003 ( .A(n_22), .Y(n_1003) );
AOI22xp5_ASAP7_75t_SL g669 ( .A1(n_23), .A2(n_187), .B1(n_597), .B2(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_24), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_25), .A2(n_361), .B1(n_848), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_26), .A2(n_87), .B1(n_875), .B2(n_876), .Y(n_1109) );
AOI22xp33_ASAP7_75t_SL g1076 ( .A1(n_27), .A2(n_200), .B1(n_575), .B2(n_576), .Y(n_1076) );
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_28), .A2(n_188), .B1(n_423), .B2(n_533), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_29), .A2(n_314), .B1(n_529), .B2(n_1001), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_30), .A2(n_148), .B1(n_483), .B2(n_821), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_31), .A2(n_109), .B1(n_459), .B2(n_746), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_32), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g1075 ( .A1(n_33), .A2(n_130), .B1(n_464), .B2(n_819), .Y(n_1075) );
AO22x2_ASAP7_75t_L g408 ( .A1(n_34), .A2(n_116), .B1(n_405), .B2(n_409), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_35), .A2(n_261), .B1(n_479), .B2(n_503), .Y(n_791) );
AOI222xp33_ASAP7_75t_L g774 ( .A1(n_36), .A2(n_185), .B1(n_291), .B2(n_533), .C1(n_641), .C2(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g1018 ( .A(n_37), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_38), .B(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_39), .A2(n_203), .B1(n_500), .B2(n_570), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_40), .A2(n_72), .B1(n_479), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g987 ( .A(n_41), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_42), .B(n_553), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_43), .Y(n_1024) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_44), .A2(n_122), .B1(n_641), .B2(n_740), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_45), .A2(n_318), .B1(n_651), .B2(n_872), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_46), .A2(n_93), .B1(n_479), .B2(n_744), .Y(n_919) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_47), .A2(n_76), .B1(n_129), .B2(n_619), .C1(n_622), .C2(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g695 ( .A(n_48), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_50), .A2(n_138), .B1(n_459), .B2(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g647 ( .A(n_51), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_52), .B(n_622), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_53), .A2(n_105), .B1(n_561), .B2(n_563), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_54), .A2(n_273), .B1(n_632), .B2(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_55), .A2(n_226), .B1(n_479), .B2(n_654), .Y(n_949) );
AO22x1_ASAP7_75t_L g1005 ( .A1(n_56), .A2(n_1006), .B1(n_1033), .B2(n_1034), .Y(n_1005) );
INVx1_ASAP7_75t_L g1033 ( .A(n_56), .Y(n_1033) );
AOI222xp33_ASAP7_75t_L g854 ( .A1(n_57), .A2(n_173), .B1(n_344), .B2(n_432), .C1(n_687), .C2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_58), .A2(n_89), .B1(n_864), .B2(n_865), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_59), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_60), .A2(n_310), .B1(n_654), .B2(n_1001), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_61), .A2(n_181), .B1(n_516), .B2(n_520), .Y(n_515) );
INVx1_ASAP7_75t_L g796 ( .A(n_62), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_63), .B(n_509), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_64), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_65), .A2(n_379), .B1(n_674), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_66), .A2(n_155), .B1(n_818), .B2(n_819), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_67), .A2(n_222), .B1(n_563), .B2(n_744), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_68), .A2(n_290), .B1(n_744), .B2(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_69), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_70), .A2(n_339), .B1(n_828), .B2(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g1108 ( .A(n_71), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_73), .A2(n_374), .B1(n_516), .B2(n_641), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g993 ( .A(n_74), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_75), .A2(n_103), .B1(n_529), .B2(n_844), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_77), .A2(n_252), .B1(n_572), .B2(n_766), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_78), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_79), .A2(n_201), .B1(n_753), .B2(n_754), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_80), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_81), .A2(n_192), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_82), .A2(n_248), .B1(n_479), .B2(n_483), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_83), .Y(n_836) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_84), .A2(n_253), .B1(n_405), .B2(n_406), .Y(n_412) );
INVx1_ASAP7_75t_L g1094 ( .A(n_84), .Y(n_1094) );
CKINVDCx20_ASAP7_75t_R g1144 ( .A(n_85), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_86), .A2(n_232), .B1(n_570), .B2(n_572), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_88), .A2(n_212), .B1(n_682), .B2(n_683), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_90), .A2(n_274), .B1(n_481), .B2(n_654), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_91), .A2(n_123), .B1(n_612), .B2(n_639), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_92), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_94), .A2(n_264), .B1(n_423), .B2(n_518), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_95), .A2(n_182), .B1(n_508), .B2(n_512), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_96), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_98), .A2(n_832), .B1(n_856), .B2(n_857), .Y(n_831) );
CKINVDCx16_ASAP7_75t_R g856 ( .A(n_98), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_99), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_100), .A2(n_371), .B1(n_656), .B2(n_770), .Y(n_769) );
AOI222xp33_ASAP7_75t_L g921 ( .A1(n_101), .A2(n_111), .B1(n_174), .B2(n_431), .C1(n_876), .C2(n_922), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g1038 ( .A1(n_102), .A2(n_1039), .B1(n_1059), .B2(n_1060), .Y(n_1038) );
INVx1_ASAP7_75t_L g1059 ( .A(n_102), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_104), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_106), .A2(n_255), .B1(n_561), .B2(n_563), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_107), .A2(n_1101), .B1(n_1120), .B2(n_1121), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g1120 ( .A(n_107), .Y(n_1120) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_108), .Y(n_888) );
INVx1_ASAP7_75t_L g685 ( .A(n_110), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_112), .A2(n_269), .B1(n_590), .B2(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_113), .A2(n_204), .B1(n_814), .B2(n_1072), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_114), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_115), .A2(n_259), .B1(n_484), .B2(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g1098 ( .A(n_116), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_117), .A2(n_294), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_118), .A2(n_267), .B1(n_677), .B2(n_706), .Y(n_1118) );
CKINVDCx20_ASAP7_75t_R g1009 ( .A(n_119), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_120), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_121), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_124), .A2(n_142), .B1(n_505), .B2(n_848), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_125), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_127), .A2(n_348), .B1(n_481), .B2(n_571), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g1104 ( .A(n_128), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_131), .A2(n_136), .B1(n_590), .B2(n_872), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_132), .Y(n_896) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_133), .A2(n_243), .B1(n_641), .B2(n_740), .Y(n_1146) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_134), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1139 ( .A1(n_135), .A2(n_208), .B1(n_473), .B2(n_698), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_137), .A2(n_272), .B1(n_597), .B2(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_139), .A2(n_153), .B1(n_753), .B2(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_140), .A2(n_345), .B1(n_502), .B2(n_504), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_141), .A2(n_221), .B1(n_972), .B2(n_973), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_143), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_145), .A2(n_198), .B1(n_641), .B2(n_770), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_146), .A2(n_298), .B1(n_525), .B2(n_746), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g1116 ( .A1(n_147), .A2(n_245), .B1(n_502), .B2(n_865), .Y(n_1116) );
AND2x6_ASAP7_75t_L g385 ( .A(n_149), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1091 ( .A(n_149), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_150), .A2(n_277), .B1(n_468), .B2(n_504), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_151), .A2(n_329), .B1(n_533), .B2(n_656), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g1068 ( .A1(n_152), .A2(n_256), .B1(n_553), .B2(n_717), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_156), .A2(n_334), .B1(n_597), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_157), .A2(n_323), .B1(n_468), .B2(n_473), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_158), .A2(n_236), .B1(n_251), .B2(n_432), .C1(n_553), .C2(n_656), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_159), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_161), .A2(n_309), .B1(n_459), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g657 ( .A(n_162), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g1081 ( .A1(n_163), .A2(n_340), .B1(n_677), .B2(n_703), .Y(n_1081) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_164), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_165), .A2(n_359), .B1(n_766), .B2(n_848), .Y(n_947) );
INVx1_ASAP7_75t_L g1032 ( .A(n_166), .Y(n_1032) );
INVx1_ASAP7_75t_L g720 ( .A(n_167), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_168), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_169), .A2(n_315), .B1(n_500), .B2(n_677), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_170), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_171), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_172), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_175), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_176), .A2(n_346), .B1(n_590), .B2(n_946), .Y(n_1002) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_177), .A2(n_244), .B1(n_405), .B2(n_409), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_177), .B(n_1096), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g1142 ( .A(n_178), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_179), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_180), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_183), .A2(n_369), .B1(n_527), .B2(n_529), .Y(n_526) );
INVx1_ASAP7_75t_L g1067 ( .A(n_184), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_186), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_189), .B(n_438), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_190), .A2(n_247), .B1(n_524), .B2(n_525), .Y(n_523) );
XOR2x2_ASAP7_75t_L g908 ( .A(n_193), .B(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_194), .A2(n_302), .B1(n_512), .B2(n_680), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_195), .Y(n_776) );
OA22x2_ASAP7_75t_L g690 ( .A1(n_196), .A2(n_691), .B1(n_692), .B2(n_724), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_196), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_197), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_199), .A2(n_288), .B1(n_459), .B2(n_561), .C(n_1028), .Y(n_1027) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_202), .A2(n_205), .B1(n_744), .B2(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g649 ( .A(n_206), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_207), .A2(n_296), .B1(n_680), .B2(n_787), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_209), .B(n_680), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_210), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_213), .A2(n_258), .B1(n_571), .B2(n_848), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_214), .B(n_512), .Y(n_1070) );
INVx1_ASAP7_75t_L g907 ( .A(n_215), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_216), .A2(n_285), .B1(n_572), .B2(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_217), .A2(n_242), .B1(n_438), .B2(n_520), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_219), .A2(n_313), .B1(n_521), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_220), .A2(n_276), .B1(n_464), .B2(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_223), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_224), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_225), .A2(n_278), .B1(n_563), .B2(n_651), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_227), .A2(n_368), .B1(n_505), .B2(n_668), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_228), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_229), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_230), .Y(n_958) );
INVx1_ASAP7_75t_L g644 ( .A(n_231), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_233), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_234), .A2(n_333), .B1(n_656), .B2(n_770), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_235), .A2(n_254), .B1(n_505), .B2(n_848), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_237), .A2(n_381), .B1(n_508), .B2(n_612), .C(n_613), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_238), .A2(n_350), .B1(n_362), .B2(n_423), .C1(n_432), .C2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_239), .A2(n_378), .B1(n_508), .B2(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g390 ( .A(n_241), .Y(n_390) );
XNOR2xp5_ASAP7_75t_L g802 ( .A(n_246), .B(n_803), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_249), .A2(n_292), .B1(n_533), .B2(n_687), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_250), .Y(n_548) );
INVx1_ASAP7_75t_L g994 ( .A(n_257), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_260), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_262), .A2(n_539), .B1(n_577), .B2(n_578), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_262), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g1106 ( .A(n_263), .Y(n_1106) );
INVx1_ASAP7_75t_L g696 ( .A(n_265), .Y(n_696) );
XOR2x2_ASAP7_75t_L g1063 ( .A(n_266), .B(n_1064), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_268), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_270), .Y(n_614) );
OA22x2_ASAP7_75t_L g727 ( .A1(n_271), .A2(n_728), .B1(n_729), .B2(n_757), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_271), .Y(n_728) );
INVx1_ASAP7_75t_L g405 ( .A(n_275), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_275), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_279), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_280), .A2(n_341), .B1(n_706), .B2(n_707), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_281), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_282), .Y(n_959) );
INVx1_ASAP7_75t_L g723 ( .A(n_283), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_284), .B(n_787), .Y(n_940) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_286), .A2(n_367), .B1(n_706), .B2(n_916), .Y(n_1135) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_289), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_293), .Y(n_806) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_295), .A2(n_383), .B(n_391), .C(n_1099), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_297), .Y(n_608) );
INVx1_ASAP7_75t_L g712 ( .A(n_299), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_300), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_301), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_303), .Y(n_840) );
INVx1_ASAP7_75t_L g1029 ( .A(n_304), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_305), .A2(n_331), .B1(n_570), .B2(n_756), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_306), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_307), .B(n_639), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_308), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_311), .A2(n_376), .B1(n_509), .B2(n_514), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_312), .A2(n_352), .B1(n_486), .B2(n_490), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_316), .Y(n_466) );
AND2x2_ASAP7_75t_L g389 ( .A(n_317), .B(n_390), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_319), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_320), .B(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_321), .Y(n_962) );
INVx1_ASAP7_75t_L g386 ( .A(n_322), .Y(n_386) );
INVx1_ASAP7_75t_L g688 ( .A(n_324), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_326), .A2(n_332), .B1(n_563), .B2(n_668), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g990 ( .A(n_327), .Y(n_990) );
INVx1_ASAP7_75t_L g652 ( .A(n_328), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_330), .Y(n_600) );
AO22x2_ASAP7_75t_L g581 ( .A1(n_336), .A2(n_582), .B1(n_624), .B2(n_625), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_336), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_337), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g967 ( .A(n_338), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_342), .A2(n_360), .B1(n_468), .B2(n_823), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_343), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_347), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_351), .Y(n_906) );
INVx1_ASAP7_75t_L g635 ( .A(n_353), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_354), .B(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_355), .B(n_532), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_356), .A2(n_373), .B1(n_524), .B2(n_946), .Y(n_945) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_357), .B(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_358), .A2(n_396), .B1(n_493), .B2(n_494), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_358), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_363), .B(n_638), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_364), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g1111 ( .A(n_365), .Y(n_1111) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_366), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_370), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_372), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_375), .A2(n_955), .B1(n_979), .B2(n_980), .Y(n_954) );
INVx1_ASAP7_75t_L g979 ( .A(n_375), .Y(n_979) );
INVx1_ASAP7_75t_L g704 ( .A(n_377), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_380), .Y(n_988) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_386), .Y(n_1090) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_387), .A2(n_1089), .B(n_1129), .Y(n_1128) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_660), .B1(n_1084), .B2(n_1085), .C(n_1086), .Y(n_391) );
INVx1_ASAP7_75t_L g1085 ( .A(n_392), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_535), .B2(n_536), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_495), .B1(n_496), .B2(n_534), .Y(n_394) );
INVx1_ASAP7_75t_L g534 ( .A(n_395), .Y(n_534) );
INVx1_ASAP7_75t_L g494 ( .A(n_396), .Y(n_494) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_456), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_421), .C(n_442), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_415), .B2(n_416), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g850 ( .A1(n_400), .A2(n_416), .B1(n_851), .B2(n_852), .C(n_853), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_400), .A2(n_958), .B1(n_959), .B2(n_960), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_400), .A2(n_960), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g544 ( .A(n_401), .Y(n_544) );
BUFx3_ASAP7_75t_L g905 ( .A(n_401), .Y(n_905) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_410), .Y(n_401) );
INVx2_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_408), .Y(n_402) );
AND2x2_ASAP7_75t_L g420 ( .A(n_403), .B(n_408), .Y(n_420) );
AND2x2_ASAP7_75t_L g461 ( .A(n_403), .B(n_427), .Y(n_461) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g428 ( .A(n_404), .B(n_414), .Y(n_428) );
AND2x2_ASAP7_75t_L g433 ( .A(n_404), .B(n_408), .Y(n_433) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_407), .Y(n_409) );
INVx2_ASAP7_75t_L g427 ( .A(n_408), .Y(n_427) );
INVx1_ASAP7_75t_L g475 ( .A(n_408), .Y(n_475) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_411), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g465 ( .A(n_411), .B(n_461), .Y(n_465) );
AND2x4_ASAP7_75t_L g511 ( .A(n_411), .B(n_482), .Y(n_511) );
AND2x6_ASAP7_75t_L g514 ( .A(n_411), .B(n_420), .Y(n_514) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g426 ( .A(n_412), .Y(n_426) );
INVx1_ASAP7_75t_L g435 ( .A(n_412), .Y(n_435) );
INVx1_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_412), .B(n_414), .Y(n_476) );
AND2x2_ASAP7_75t_L g434 ( .A(n_413), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g472 ( .A(n_414), .B(n_455), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_416), .A2(n_542), .B1(n_543), .B2(n_545), .Y(n_541) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g636 ( .A(n_418), .Y(n_636) );
BUFx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g711 ( .A(n_419), .Y(n_711) );
AND2x2_ASAP7_75t_L g471 ( .A(n_420), .B(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g484 ( .A(n_420), .B(n_434), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_420), .B(n_472), .Y(n_594) );
OAI222xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_429), .B1(n_430), .B2(n_436), .C1(n_437), .C2(n_441), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g549 ( .A(n_423), .Y(n_549) );
BUFx4f_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_424), .Y(n_622) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_424), .Y(n_656) );
BUFx2_ASAP7_75t_L g687 ( .A(n_424), .Y(n_687) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_424), .Y(n_719) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g440 ( .A(n_426), .Y(n_440) );
INVx1_ASAP7_75t_L g447 ( .A(n_427), .Y(n_447) );
AND2x4_ASAP7_75t_L g439 ( .A(n_428), .B(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_428), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g518 ( .A(n_428), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g547 ( .A(n_431), .Y(n_547) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx4_ASAP7_75t_L g621 ( .A(n_432), .Y(n_621) );
BUFx3_ASAP7_75t_L g775 ( .A(n_432), .Y(n_775) );
INVx2_ASAP7_75t_L g781 ( .A(n_432), .Y(n_781) );
AND2x6_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g452 ( .A(n_433), .Y(n_452) );
AND2x4_ASAP7_75t_L g521 ( .A(n_433), .B(n_454), .Y(n_521) );
AND2x2_ASAP7_75t_L g460 ( .A(n_434), .B(n_461), .Y(n_460) );
AND2x6_ASAP7_75t_L g481 ( .A(n_434), .B(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_437), .A2(n_621), .B1(n_900), .B2(n_901), .C(n_902), .Y(n_899) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g623 ( .A(n_438), .Y(n_623) );
BUFx2_ASAP7_75t_L g855 ( .A(n_438), .Y(n_855) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx12f_ASAP7_75t_L g533 ( .A(n_439), .Y(n_533) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_439), .Y(n_553) );
INVx1_ASAP7_75t_L g809 ( .A(n_439), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_448), .B2(n_449), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_444), .A2(n_1018), .B1(n_1019), .B2(n_1020), .Y(n_1017) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_SL g897 ( .A(n_445), .Y(n_897) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_446), .Y(n_556) );
BUFx3_ASAP7_75t_L g615 ( .A(n_446), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_446), .A2(n_617), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AND2x2_ASAP7_75t_L g766 ( .A(n_447), .B(n_492), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_449), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_554) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g1020 ( .A(n_450), .Y(n_1020) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g617 ( .A(n_451), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_451), .A2(n_896), .B1(n_897), .B2(n_898), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_451), .A2(n_615), .B1(n_993), .B2(n_994), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_451), .A2(n_556), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_477), .Y(n_456) );
OAI221xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_462), .B1(n_463), .B2(n_466), .C(n_467), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_460), .Y(n_571) );
INVx2_ASAP7_75t_L g586 ( .A(n_460), .Y(n_586) );
BUFx2_ASAP7_75t_SL g872 ( .A(n_460), .Y(n_872) );
AND2x2_ASAP7_75t_L g489 ( .A(n_461), .B(n_472), .Y(n_489) );
AND2x4_ASAP7_75t_L g491 ( .A(n_461), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_461), .B(n_472), .Y(n_607) );
INVx4_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
INVx3_ASAP7_75t_L g632 ( .A(n_463), .Y(n_632) );
OAI221xp5_ASAP7_75t_SL g693 ( .A1(n_463), .A2(n_694), .B1(n_695), .B2(n_696), .C(n_697), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_463), .A2(n_891), .B1(n_892), .B2(n_893), .Y(n_890) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g573 ( .A(n_465), .Y(n_573) );
BUFx3_ASAP7_75t_L g590 ( .A(n_465), .Y(n_590) );
BUFx3_ASAP7_75t_L g756 ( .A(n_465), .Y(n_756) );
BUFx3_ASAP7_75t_L g977 ( .A(n_465), .Y(n_977) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx5_ASAP7_75t_L g503 ( .A(n_470), .Y(n_503) );
INVx4_ASAP7_75t_L g671 ( .A(n_470), .Y(n_671) );
INVx1_ASAP7_75t_L g749 ( .A(n_470), .Y(n_749) );
INVx2_ASAP7_75t_L g848 ( .A(n_470), .Y(n_848) );
INVx3_ASAP7_75t_L g864 ( .A(n_470), .Y(n_864) );
INVx8_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx6_ASAP7_75t_SL g505 ( .A(n_474), .Y(n_505) );
INVx1_ASAP7_75t_SL g823 ( .A(n_474), .Y(n_823) );
INVx1_ASAP7_75t_L g886 ( .A(n_474), .Y(n_886) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
INVx1_ASAP7_75t_L g492 ( .A(n_476), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_478), .B(n_485), .Y(n_477) );
INVx4_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_480), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_599) );
INVx3_ASAP7_75t_L g651 ( .A(n_480), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_480), .A2(n_701), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_700) );
INVx2_ASAP7_75t_SL g972 ( .A(n_480), .Y(n_972) );
INVx4_ASAP7_75t_L g1031 ( .A(n_480), .Y(n_1031) );
INVx11_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx11_ASAP7_75t_L g528 ( .A(n_481), .Y(n_528) );
INVx1_ASAP7_75t_L g602 ( .A(n_483), .Y(n_602) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx6_ASAP7_75t_L g530 ( .A(n_484), .Y(n_530) );
BUFx3_ASAP7_75t_L g567 ( .A(n_484), .Y(n_567) );
BUFx3_ASAP7_75t_L g744 ( .A(n_484), .Y(n_744) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx4f_ASAP7_75t_SL g706 ( .A(n_488), .Y(n_706) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g524 ( .A(n_489), .Y(n_524) );
BUFx3_ASAP7_75t_L g668 ( .A(n_489), .Y(n_668) );
BUFx3_ASAP7_75t_L g746 ( .A(n_489), .Y(n_746) );
BUFx2_ASAP7_75t_L g610 ( .A(n_490), .Y(n_610) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g525 ( .A(n_491), .Y(n_525) );
BUFx3_ASAP7_75t_L g563 ( .A(n_491), .Y(n_563) );
BUFx2_ASAP7_75t_SL g677 ( .A(n_491), .Y(n_677) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_491), .Y(n_707) );
BUFx3_ASAP7_75t_L g828 ( .A(n_491), .Y(n_828) );
INVx1_ASAP7_75t_L g917 ( .A(n_491), .Y(n_917) );
BUFx2_ASAP7_75t_L g946 ( .A(n_491), .Y(n_946) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_496), .B(n_628), .Y(n_627) );
NAND4xp75_ASAP7_75t_L g497 ( .A(n_498), .B(n_506), .C(n_522), .D(n_531), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g576 ( .A(n_505), .Y(n_576) );
BUFx2_ASAP7_75t_L g597 ( .A(n_505), .Y(n_597) );
BUFx2_ASAP7_75t_L g865 ( .A(n_505), .Y(n_865) );
BUFx4f_ASAP7_75t_SL g1026 ( .A(n_505), .Y(n_1026) );
AND2x2_ASAP7_75t_SL g506 ( .A(n_507), .B(n_515), .Y(n_506) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx5_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g639 ( .A(n_510), .Y(n_639) );
INVx2_ASAP7_75t_L g680 ( .A(n_510), .Y(n_680) );
INVx2_ASAP7_75t_L g1072 ( .A(n_510), .Y(n_1072) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g814 ( .A(n_513), .Y(n_814) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g612 ( .A(n_514), .Y(n_612) );
BUFx4f_ASAP7_75t_L g787 ( .A(n_514), .Y(n_787) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g714 ( .A(n_517), .Y(n_714) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g682 ( .A(n_518), .Y(n_682) );
BUFx2_ASAP7_75t_L g740 ( .A(n_518), .Y(n_740) );
BUFx3_ASAP7_75t_L g770 ( .A(n_518), .Y(n_770) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g641 ( .A(n_521), .Y(n_641) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_521), .Y(n_683) );
BUFx2_ASAP7_75t_SL g922 ( .A(n_521), .Y(n_922) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
BUFx2_ASAP7_75t_L g826 ( .A(n_524), .Y(n_826) );
INVxp67_ASAP7_75t_L g646 ( .A(n_525), .Y(n_646) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g675 ( .A(n_528), .Y(n_675) );
INVx2_ASAP7_75t_SL g821 ( .A(n_528), .Y(n_821) );
INVx5_ASAP7_75t_SL g846 ( .A(n_528), .Y(n_846) );
INVx4_ASAP7_75t_L g1001 ( .A(n_528), .Y(n_1001) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g654 ( .A(n_530), .Y(n_654) );
INVx2_ASAP7_75t_L g703 ( .A(n_530), .Y(n_703) );
INVx2_ASAP7_75t_L g973 ( .A(n_530), .Y(n_973) );
INVx1_ASAP7_75t_L g722 ( .A(n_532), .Y(n_722) );
BUFx4f_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g877 ( .A(n_533), .Y(n_877) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_579), .B1(n_658), .B2(n_659), .Y(n_537) );
INVx1_ASAP7_75t_L g658 ( .A(n_538), .Y(n_658) );
INVx2_ASAP7_75t_L g578 ( .A(n_539), .Y(n_578) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_558), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_546), .C(n_554), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_543), .A2(n_709), .B1(n_710), .B2(n_712), .C(n_713), .Y(n_708) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_544), .Y(n_1010) );
INVx2_ASAP7_75t_L g1105 ( .A(n_544), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .C(n_551), .Y(n_546) );
OAI222xp33_ASAP7_75t_L g805 ( .A1(n_547), .A2(n_806), .B1(n_807), .B2(n_808), .C1(n_809), .C2(n_810), .Y(n_805) );
OAI221xp5_ASAP7_75t_L g1044 ( .A1(n_547), .A2(n_1045), .B1(n_1046), .B2(n_1047), .C(n_1048), .Y(n_1044) );
OAI222xp33_ASAP7_75t_L g1141 ( .A1(n_547), .A2(n_549), .B1(n_809), .B2(n_1142), .C1(n_1143), .C2(n_1144), .Y(n_1141) );
OAI222xp33_ASAP7_75t_L g731 ( .A1(n_549), .A2(n_732), .B1(n_734), .B2(n_735), .C1(n_736), .C2(n_737), .Y(n_731) );
OAI221xp5_ASAP7_75t_SL g961 ( .A1(n_549), .A2(n_620), .B1(n_962), .B2(n_963), .C(n_964), .Y(n_961) );
BUFx4f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g736 ( .A(n_553), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_568), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_574), .Y(n_568) );
BUFx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_571), .Y(n_674) );
INVx3_ASAP7_75t_L g694 ( .A(n_571), .Y(n_694) );
BUFx3_ASAP7_75t_L g753 ( .A(n_571), .Y(n_753) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g659 ( .A(n_579), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_626), .B2(n_627), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g625 ( .A(n_582), .Y(n_625) );
AND4x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_598), .C(n_611), .D(n_618), .Y(n_582) );
NOR2xp33_ASAP7_75t_SL g583 ( .A(n_584), .B(n_591), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_584) );
INVx3_ASAP7_75t_L g951 ( .A(n_586), .Y(n_951) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g841 ( .A(n_590), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_593), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
BUFx2_ASAP7_75t_R g593 ( .A(n_594), .Y(n_593) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_603), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_608), .B2(n_609), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g645 ( .A(n_606), .Y(n_645) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_616), .B2(n_617), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_617), .A2(n_897), .B1(n_966), .B2(n_967), .Y(n_965) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_620), .A2(n_685), .B(n_686), .Y(n_684) );
OAI21xp5_ASAP7_75t_SL g1107 ( .A1(n_620), .A2(n_1108), .B(n_1109), .Y(n_1107) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g715 ( .A1(n_621), .A2(n_716), .B1(n_720), .B2(n_721), .C1(n_722), .C2(n_723), .Y(n_715) );
INVx4_ASAP7_75t_L g733 ( .A(n_621), .Y(n_733) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
XOR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_657), .Y(n_628) );
NAND4xp75_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .C(n_642), .D(n_655), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
OA211x2_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B(n_637), .C(n_640), .Y(n_634) );
OA211x2_ASAP7_75t_L g866 ( .A1(n_636), .A2(n_867), .B(n_868), .C(n_869), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_636), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_648), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_646), .B2(n_647), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_645), .A2(n_702), .B1(n_835), .B2(n_836), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_645), .A2(n_653), .B1(n_888), .B2(n_889), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_656), .Y(n_875) );
INVx1_ASAP7_75t_L g1084 ( .A(n_660), .Y(n_1084) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_929), .Y(n_660) );
XOR2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_801), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_689), .B2(n_800), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
XOR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_688), .Y(n_664) );
NOR4xp75_ASAP7_75t_L g665 ( .A(n_666), .B(n_672), .C(n_678), .D(n_684), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g1080 ( .A(n_668), .Y(n_1080) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g699 ( .A(n_671), .Y(n_699) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_SL g839 ( .A(n_674), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g800 ( .A(n_689), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_725), .B1(n_798), .B2(n_799), .Y(n_689) );
INVx1_ASAP7_75t_L g798 ( .A(n_690), .Y(n_798) );
INVx1_ASAP7_75t_L g724 ( .A(n_692), .Y(n_724) );
OR4x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_700), .C(n_708), .D(n_715), .Y(n_692) );
INVx2_ASAP7_75t_L g818 ( .A(n_694), .Y(n_818) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_702), .A2(n_1029), .B1(n_1030), .B2(n_1032), .Y(n_1028) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g893 ( .A(n_707), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_710), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_710), .A2(n_905), .B1(n_987), .B2(n_988), .Y(n_986) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g960 ( .A(n_711), .Y(n_960) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx4_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g807 ( .A(n_719), .Y(n_807) );
INVx1_ASAP7_75t_L g799 ( .A(n_725), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_758), .B2(n_759), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g757 ( .A(n_729), .Y(n_757) );
NAND3x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_742), .C(n_750), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_738), .Y(n_730) );
OAI21xp5_ASAP7_75t_SL g1066 ( .A1(n_732), .A2(n_1067), .B(n_1068), .Y(n_1066) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
BUFx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AO22x2_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_777), .B2(n_797), .Y(n_759) );
INVx2_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
XOR2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_776), .Y(n_761) );
NAND4xp75_ASAP7_75t_L g762 ( .A(n_763), .B(n_767), .C(n_771), .D(n_774), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AND2x2_ASAP7_75t_SL g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx3_ASAP7_75t_L g936 ( .A(n_775), .Y(n_936) );
INVx2_ASAP7_75t_L g797 ( .A(n_777), .Y(n_797) );
XOR2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_796), .Y(n_777) );
NAND2x1_ASAP7_75t_L g778 ( .A(n_779), .B(n_789), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_784), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_782), .B(n_783), .Y(n_780) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .C(n_788), .Y(n_784) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_793), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_829), .B1(n_927), .B2(n_928), .Y(n_801) );
INVx1_ASAP7_75t_L g927 ( .A(n_802), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_815), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_811), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_824), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_822), .Y(n_816) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g928 ( .A(n_829), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_858), .B1(n_925), .B2(n_926), .Y(n_829) );
INVx1_ASAP7_75t_L g926 ( .A(n_830), .Y(n_926) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_SL g857 ( .A(n_832), .Y(n_857) );
AND4x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_842), .C(n_849), .D(n_854), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_837), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_837) );
AND2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_847), .Y(n_842) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g925 ( .A(n_858), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_879), .B1(n_923), .B2(n_924), .Y(n_858) );
INVx3_ASAP7_75t_SL g924 ( .A(n_859), .Y(n_924) );
XOR2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_878), .Y(n_859) );
NAND4xp75_ASAP7_75t_L g860 ( .A(n_861), .B(n_866), .C(n_870), .D(n_874), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_873), .Y(n_870) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_875), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_875), .Y(n_1046) );
INVx3_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g923 ( .A(n_879), .Y(n_923) );
XOR2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_908), .Y(n_879) );
XOR2xp5_ASAP7_75t_SL g880 ( .A(n_881), .B(n_907), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_894), .Y(n_881) );
NOR3xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_887), .C(n_890), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
NOR3xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_899), .C(n_903), .Y(n_894) );
NAND4xp75_ASAP7_75t_L g909 ( .A(n_910), .B(n_913), .C(n_918), .D(n_921), .Y(n_909) );
AND2x2_ASAP7_75t_SL g910 ( .A(n_911), .B(n_912), .Y(n_910) );
AND2x2_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_981), .B1(n_1082), .B2(n_1083), .Y(n_929) );
INVx1_ASAP7_75t_L g1082 ( .A(n_930), .Y(n_1082) );
OAI22xp5_ASAP7_75t_SL g930 ( .A1(n_931), .A2(n_932), .B1(n_953), .B2(n_954), .Y(n_930) );
INVx3_ASAP7_75t_SL g931 ( .A(n_932), .Y(n_931) );
XNOR2xp5_ASAP7_75t_L g1062 ( .A(n_932), .B(n_1063), .Y(n_1062) );
XOR2x2_ASAP7_75t_L g932 ( .A(n_933), .B(n_952), .Y(n_932) );
NAND2xp5_ASAP7_75t_SL g933 ( .A(n_934), .B(n_943), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_939), .Y(n_934) );
OAI21xp5_ASAP7_75t_SL g935 ( .A1(n_936), .A2(n_937), .B(n_938), .Y(n_935) );
OAI21xp33_ASAP7_75t_L g989 ( .A1(n_936), .A2(n_990), .B(n_991), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g1012 ( .A1(n_936), .A2(n_1013), .B1(n_1014), .B2(n_1015), .C(n_1016), .Y(n_1012) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .C(n_942), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_948), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_947), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx2_ASAP7_75t_L g980 ( .A(n_955), .Y(n_980) );
AND2x2_ASAP7_75t_SL g955 ( .A(n_956), .B(n_968), .Y(n_955) );
NOR3xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_961), .C(n_965), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_960), .A2(n_1009), .B1(n_1010), .B2(n_1011), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_969), .B(n_974), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_978), .Y(n_974) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g1083 ( .A(n_981), .Y(n_1083) );
XOR2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_1036), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_1004), .B1(n_1005), .B2(n_1035), .Y(n_982) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_983), .Y(n_1035) );
XOR2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_1003), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_995), .Y(n_984) );
NOR3xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .C(n_992), .Y(n_985) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_996), .B(n_999), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1002), .Y(n_999) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1006), .Y(n_1034) );
AND3x1_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1021), .C(n_1027), .Y(n_1006) );
NOR3xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1012), .C(n_1017), .Y(n_1007) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1038), .B1(n_1061), .B2(n_1062), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1039), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1052), .Y(n_1039) );
NOR3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1044), .C(n_1049), .Y(n_1040) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1056), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .Y(n_1056) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
NAND3x2_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1074), .C(n_1077), .Y(n_1064) );
NOR2x1_ASAP7_75t_SL g1065 ( .A(n_1066), .B(n_1069), .Y(n_1065) );
NAND3xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1071), .C(n_1073), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1076), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1081), .Y(n_1077) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_SL g1086 ( .A(n_1087), .Y(n_1086) );
NOR2x1_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1092), .Y(n_1087) );
OR2x2_ASAP7_75t_SL g1151 ( .A(n_1088), .B(n_1093), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1091), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1090), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1090), .B(n_1126), .Y(n_1129) );
CKINVDCx16_ASAP7_75t_R g1126 ( .A(n_1091), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g1092 ( .A(n_1093), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1098), .Y(n_1096) );
OAI322xp33_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1122), .A3(n_1123), .B1(n_1127), .B2(n_1130), .C1(n_1131), .C2(n_1149), .Y(n_1099) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1101), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1113), .Y(n_1101) );
NOR3xp33_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1107), .C(n_1110), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1117), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1116), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1119), .Y(n_1117) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
CKINVDCx20_ASAP7_75t_R g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1132), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1140), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1137), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1139), .Y(n_1137) );
NOR2xp33_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1145), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1147), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_1150), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_1151), .Y(n_1150) );
endmodule