module real_aes_18099_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_0), .Y(n_797) );
AND2x4_ASAP7_75t_L g830 ( .A(n_1), .B(n_831), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_2), .A2(n_4), .B1(n_179), .B2(n_506), .Y(n_505) );
OAI22x1_ASAP7_75t_R g115 ( .A1(n_3), .A2(n_45), .B1(n_116), .B2(n_117), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_3), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_5), .A2(n_43), .B1(n_136), .B2(n_159), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_6), .A2(n_26), .B1(n_159), .B2(n_235), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_7), .A2(n_17), .B1(n_178), .B2(n_214), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_8), .A2(n_60), .B1(n_196), .B2(n_237), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_9), .A2(n_18), .B1(n_135), .B2(n_136), .Y(n_522) );
INVx1_ASAP7_75t_L g831 ( .A(n_10), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_11), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_12), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_13), .A2(n_19), .B1(n_195), .B2(n_198), .Y(n_194) );
OR2x2_ASAP7_75t_L g113 ( .A(n_14), .B(n_39), .Y(n_113) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_15), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_16), .Y(n_218) );
INVx2_ASAP7_75t_L g820 ( .A(n_20), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_21), .A2(n_97), .B1(n_178), .B2(n_179), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_22), .A2(n_40), .B1(n_144), .B2(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_23), .B(n_139), .Y(n_138) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_24), .A2(n_57), .B(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_25), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_27), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_28), .B(n_141), .Y(n_492) );
INVx4_ASAP7_75t_R g534 ( .A(n_29), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_30), .A2(n_48), .B1(n_164), .B2(n_165), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_31), .A2(n_54), .B1(n_165), .B2(n_178), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_32), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_33), .B(n_144), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_34), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_35), .B(n_159), .Y(n_499) );
INVx1_ASAP7_75t_L g508 ( .A(n_36), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_SL g574 ( .A1(n_37), .A2(n_136), .B(n_140), .C(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_38), .A2(n_55), .B1(n_136), .B2(n_165), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_41), .A2(n_85), .B1(n_136), .B2(n_234), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_42), .A2(n_47), .B1(n_135), .B2(n_136), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_44), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_45), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_46), .A2(n_59), .B1(n_178), .B2(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g496 ( .A(n_49), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_50), .B(n_136), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_51), .Y(n_555) );
INVx2_ASAP7_75t_L g108 ( .A(n_52), .Y(n_108) );
BUFx3_ASAP7_75t_L g111 ( .A(n_53), .Y(n_111) );
INVx1_ASAP7_75t_L g816 ( .A(n_53), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_56), .A2(n_86), .B1(n_136), .B2(n_165), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_58), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_61), .A2(n_74), .B1(n_164), .B2(n_182), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_62), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_63), .A2(n_76), .B1(n_135), .B2(n_136), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_64), .A2(n_95), .B1(n_178), .B2(n_198), .Y(n_224) );
INVx1_ASAP7_75t_L g131 ( .A(n_65), .Y(n_131) );
AND2x4_ASAP7_75t_L g150 ( .A(n_66), .B(n_151), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_67), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_67), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_68), .A2(n_88), .B1(n_164), .B2(n_165), .Y(n_504) );
AO22x1_ASAP7_75t_L g513 ( .A1(n_69), .A2(n_75), .B1(n_211), .B2(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g151 ( .A(n_70), .Y(n_151) );
AND2x2_ASAP7_75t_L g577 ( .A(n_71), .B(n_153), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_72), .B(n_237), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_73), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_77), .B(n_159), .Y(n_556) );
INVx2_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_79), .B(n_153), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_80), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_81), .A2(n_96), .B1(n_165), .B2(n_237), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_82), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_83), .B(n_186), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_84), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_87), .B(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_89), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_90), .B(n_153), .Y(n_552) );
INVx1_ASAP7_75t_L g468 ( .A(n_91), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_91), .B(n_815), .Y(n_814) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_92), .B(n_139), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_93), .A2(n_201), .B(n_237), .C(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g536 ( .A(n_94), .B(n_537), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g823 ( .A(n_98), .Y(n_823) );
NAND2xp33_ASAP7_75t_L g560 ( .A(n_99), .B(n_145), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_805), .B(n_825), .C(n_833), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_114), .B(n_796), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx12f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x6_ASAP7_75t_SL g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_108), .B(n_802), .Y(n_801) );
INVx3_ASAP7_75t_L g808 ( .A(n_108), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_108), .B(n_843), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1_ASAP7_75t_L g804 ( .A(n_111), .B(n_113), .Y(n_804) );
AND2x6_ASAP7_75t_SL g813 ( .A(n_112), .B(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
XNOR2x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
AOI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_465), .B1(n_469), .B2(n_793), .Y(n_118) );
XNOR2x1_ASAP7_75t_SL g817 ( .A(n_119), .B(n_818), .Y(n_817) );
NAND2x1p5_ASAP7_75t_L g119 ( .A(n_120), .B(n_409), .Y(n_119) );
NOR3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_327), .C(n_364), .Y(n_120) );
NAND4xp75_ASAP7_75t_L g121 ( .A(n_122), .B(n_247), .C(n_281), .D(n_311), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI32xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_169), .A3(n_219), .B1(n_228), .B2(n_242), .Y(n_123) );
OR2x2_ASAP7_75t_L g228 ( .A(n_124), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_125), .A2(n_439), .B(n_441), .Y(n_438) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_154), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_126), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g310 ( .A(n_126), .B(n_256), .Y(n_310) );
AND2x2_ASAP7_75t_L g405 ( .A(n_126), .B(n_221), .Y(n_405) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx2_ASAP7_75t_L g254 ( .A(n_127), .Y(n_254) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_152), .Y(n_127) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_128), .A2(n_132), .B(n_152), .Y(n_287) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g153 ( .A(n_129), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_129), .B(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g216 ( .A(n_129), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_129), .B(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_129), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g500 ( .A(n_129), .B(n_483), .Y(n_500) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g186 ( .A(n_130), .Y(n_186) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_142), .B(n_148), .Y(n_132) );
O2A1O1Ixp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_138), .C(n_140), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_135), .A2(n_555), .B(n_556), .C(n_557), .Y(n_554) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
INVx1_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_137), .Y(n_139) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx1_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx1_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
INVx1_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_137), .Y(n_215) );
INVx2_ASAP7_75t_L g235 ( .A(n_137), .Y(n_235) );
INVx1_ASAP7_75t_L g237 ( .A(n_137), .Y(n_237) );
INVx3_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_139), .Y(n_514) );
INVx6_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_140), .A2(n_513), .B(n_515), .C(n_518), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_140), .A2(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_140), .B(n_513), .Y(n_586) );
BUFx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g162 ( .A(n_141), .Y(n_162) );
INVx1_ASAP7_75t_L g201 ( .A(n_141), .Y(n_201) );
INVx1_ASAP7_75t_L g495 ( .A(n_141), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_147), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g164 ( .A(n_145), .Y(n_164) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_145), .A2(n_215), .B1(n_534), .B2(n_535), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_147), .A2(n_158), .B1(n_160), .B2(n_163), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_147), .A2(n_160), .B1(n_177), .B2(n_181), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_147), .A2(n_194), .B1(n_199), .B2(n_200), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_147), .A2(n_160), .B1(n_210), .B2(n_213), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_147), .A2(n_200), .B1(n_224), .B2(n_225), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_147), .A2(n_233), .B1(n_236), .B2(n_238), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_147), .A2(n_160), .B1(n_272), .B2(n_273), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_147), .A2(n_480), .B1(n_481), .B2(n_482), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_147), .A2(n_238), .B1(n_504), .B2(n_505), .Y(n_503) );
OAI22x1_ASAP7_75t_L g521 ( .A1(n_147), .A2(n_238), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_SL g239 ( .A(n_149), .Y(n_239) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx10_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
BUFx10_ASAP7_75t_L g483 ( .A(n_150), .Y(n_483) );
INVx1_ASAP7_75t_L g519 ( .A(n_150), .Y(n_519) );
INVx2_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_153), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g278 ( .A(n_154), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_154), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_155), .Y(n_265) );
INVx1_ASAP7_75t_L g309 ( .A(n_155), .Y(n_309) );
AND2x2_ASAP7_75t_L g353 ( .A(n_155), .B(n_287), .Y(n_353) );
OR2x2_ASAP7_75t_L g407 ( .A(n_155), .B(n_231), .Y(n_407) );
AO31x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .A3(n_166), .B(n_167), .Y(n_155) );
INVx2_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
AO31x2_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_193), .A3(n_202), .B(n_204), .Y(n_192) );
AO31x2_ASAP7_75t_L g208 ( .A1(n_156), .A2(n_209), .A3(n_216), .B(n_217), .Y(n_208) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_156), .A2(n_189), .A3(n_521), .B(n_524), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_159), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g482 ( .A(n_161), .Y(n_482) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g558 ( .A(n_162), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_165), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g506 ( .A(n_165), .Y(n_506) );
AO31x2_ASAP7_75t_L g478 ( .A1(n_166), .A2(n_479), .A3(n_483), .B(n_484), .Y(n_478) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_170), .A2(n_333), .B1(n_425), .B2(n_427), .Y(n_424) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_190), .Y(n_170) );
INVx4_ASAP7_75t_L g250 ( .A(n_171), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_171), .A2(n_230), .B1(n_262), .B2(n_264), .Y(n_261) );
OR2x2_ASAP7_75t_L g267 ( .A(n_171), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g386 ( .A(n_171), .B(n_285), .Y(n_386) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g306 ( .A(n_172), .B(n_191), .Y(n_306) );
AND2x2_ASAP7_75t_L g397 ( .A(n_172), .B(n_269), .Y(n_397) );
AND2x2_ASAP7_75t_L g452 ( .A(n_172), .B(n_208), .Y(n_452) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g246 ( .A(n_173), .Y(n_246) );
AND2x4_ASAP7_75t_L g373 ( .A(n_173), .B(n_269), .Y(n_373) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .A3(n_183), .B(n_187), .Y(n_173) );
AO31x2_ASAP7_75t_L g222 ( .A1(n_174), .A2(n_202), .A3(n_223), .B(n_226), .Y(n_222) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_175), .A2(n_529), .B(n_532), .Y(n_528) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_180), .B(n_572), .Y(n_571) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_183), .A2(n_239), .A3(n_271), .B(n_274), .Y(n_270) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_183), .A2(n_528), .B(n_536), .Y(n_527) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g204 ( .A(n_185), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_185), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g189 ( .A(n_186), .Y(n_189) );
INVx2_ASAP7_75t_L g203 ( .A(n_186), .Y(n_203) );
OAI21xp33_ASAP7_75t_L g518 ( .A1(n_186), .A2(n_517), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_189), .B(n_275), .Y(n_274) );
NAND2x1_ASAP7_75t_L g249 ( .A(n_190), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_190), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_206), .Y(n_190) );
INVx2_ASAP7_75t_L g244 ( .A(n_191), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_191), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g292 ( .A(n_191), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_191), .B(n_294), .Y(n_319) );
AND2x2_ASAP7_75t_L g322 ( .A(n_191), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g382 ( .A(n_191), .Y(n_382) );
INVx4_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_192), .B(n_207), .Y(n_260) );
BUFx2_ASAP7_75t_L g298 ( .A(n_192), .Y(n_298) );
AND2x2_ASAP7_75t_L g347 ( .A(n_192), .B(n_208), .Y(n_347) );
AND2x2_ASAP7_75t_L g389 ( .A(n_192), .B(n_270), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_192), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_197), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g238 ( .A(n_201), .Y(n_238) );
AO31x2_ASAP7_75t_L g502 ( .A1(n_202), .A2(n_239), .A3(n_503), .B(n_507), .Y(n_502) );
AOI21x1_ASAP7_75t_L g566 ( .A1(n_202), .A2(n_567), .B(n_577), .Y(n_566) );
BUFx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_203), .B(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_203), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_203), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g537 ( .A(n_203), .Y(n_537) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_208), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g300 ( .A(n_208), .B(n_270), .Y(n_300) );
INVx1_ASAP7_75t_L g323 ( .A(n_208), .Y(n_323) );
INVx2_ASAP7_75t_L g343 ( .A(n_208), .Y(n_343) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_208), .Y(n_388) );
OAI21xp33_ASAP7_75t_SL g491 ( .A1(n_211), .A2(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AO31x2_ASAP7_75t_L g231 ( .A1(n_216), .A2(n_232), .A3(n_239), .B(n_240), .Y(n_231) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g307 ( .A(n_220), .B(n_308), .Y(n_307) );
NOR2x1p5_ASAP7_75t_L g413 ( .A(n_220), .B(n_407), .Y(n_413) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x4_ASAP7_75t_L g230 ( .A(n_221), .B(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g263 ( .A(n_221), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_221), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_221), .B(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g255 ( .A(n_222), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g313 ( .A(n_222), .B(n_231), .Y(n_313) );
BUFx2_ASAP7_75t_L g426 ( .A(n_222), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_228), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g464 ( .A(n_228), .Y(n_464) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g400 ( .A(n_230), .Y(n_400) );
AND2x4_ASAP7_75t_L g423 ( .A(n_230), .B(n_353), .Y(n_423) );
AND2x2_ASAP7_75t_L g447 ( .A(n_230), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g256 ( .A(n_231), .Y(n_256) );
BUFx2_ASAP7_75t_L g280 ( .A(n_231), .Y(n_280) );
INVx1_ASAP7_75t_L g336 ( .A(n_231), .Y(n_336) );
OR2x2_ASAP7_75t_L g458 ( .A(n_231), .B(n_315), .Y(n_458) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_235), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_238), .B(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_245), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_245), .Y(n_325) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g266 ( .A(n_246), .Y(n_266) );
OR2x2_ASAP7_75t_L g303 ( .A(n_246), .B(n_295), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_251), .B(n_257), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_252), .A2(n_346), .B1(n_348), .B2(n_351), .Y(n_345) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
OR2x2_ASAP7_75t_L g391 ( .A(n_254), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g399 ( .A(n_254), .Y(n_399) );
AND2x2_ASAP7_75t_L g412 ( .A(n_254), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g374 ( .A(n_255), .B(n_353), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B1(n_267), .B2(n_276), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g326 ( .A(n_260), .Y(n_326) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g284 ( .A(n_263), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g352 ( .A(n_263), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g361 ( .A(n_263), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_263), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_264), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g349 ( .A(n_266), .B(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g363 ( .A(n_266), .Y(n_363) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
AND2x4_ASAP7_75t_L g342 ( .A(n_270), .B(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_270), .Y(n_358) );
INVx1_ASAP7_75t_L g422 ( .A(n_270), .Y(n_422) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
AND2x4_ASAP7_75t_L g314 ( .A(n_278), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g331 ( .A(n_278), .Y(n_331) );
INVx1_ASAP7_75t_L g289 ( .A(n_280), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_290), .B1(n_301), .B2(n_307), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_286), .Y(n_339) );
INVx1_ASAP7_75t_L g315 ( .A(n_287), .Y(n_315) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_291), .B(n_296), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_292), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g444 ( .A(n_293), .Y(n_444) );
INVx1_ASAP7_75t_L g463 ( .A(n_293), .Y(n_463) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_297), .B(n_363), .Y(n_440) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g456 ( .A(n_298), .Y(n_456) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
INVx2_ASAP7_75t_L g394 ( .A(n_302), .Y(n_394) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g383 ( .A(n_303), .Y(n_383) );
AND2x4_ASAP7_75t_L g385 ( .A(n_304), .B(n_342), .Y(n_385) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_308), .A2(n_454), .B1(n_457), .B2(n_459), .Y(n_453) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g378 ( .A(n_309), .Y(n_378) );
INVx1_ASAP7_75t_L g332 ( .A(n_310), .Y(n_332) );
AND2x4_ASAP7_75t_L g425 ( .A(n_310), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g433 ( .A(n_310), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .Y(n_311) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_SL g376 ( .A(n_313), .Y(n_376) );
INVx2_ASAP7_75t_L g392 ( .A(n_313), .Y(n_392) );
INVx1_ASAP7_75t_L g419 ( .A(n_314), .Y(n_419) );
AND2x2_ASAP7_75t_L g450 ( .A(n_314), .B(n_361), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .C(n_324), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_321), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g362 ( .A(n_322), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_322), .B(n_397), .Y(n_430) );
INVx1_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_325), .B(n_389), .Y(n_415) );
INVx1_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
NAND3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_344), .C(n_354), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_333), .B(n_340), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g448 ( .A(n_331), .Y(n_448) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI32xp33_ASAP7_75t_L g384 ( .A1(n_335), .A2(n_385), .A3(n_386), .B1(n_387), .B2(n_390), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_335), .B(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_342), .B(n_363), .Y(n_403) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_347), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g408 ( .A(n_347), .B(n_357), .Y(n_408) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g436 ( .A(n_350), .Y(n_436) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_352), .A2(n_355), .B1(n_359), .B2(n_362), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_353), .B(n_361), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_355), .A2(n_413), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g451 ( .A(n_357), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_402), .B1(n_404), .B2(n_408), .Y(n_401) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g443 ( .A(n_363), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_365), .B(n_384), .C(n_393), .D(n_401), .Y(n_364) );
O2A1O1Ixp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_371), .B(n_374), .C(n_375), .Y(n_365) );
NOR2x1_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g429 ( .A(n_373), .B(n_388), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_373), .B(n_456), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_379), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_380), .A2(n_418), .B1(n_420), .B2(n_423), .Y(n_417) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_385), .A2(n_390), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_398), .Y(n_393) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_R g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_408), .A2(n_425), .B1(n_462), .B2(n_464), .Y(n_461) );
NOR3x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_431), .C(n_445), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_424), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g437 ( .A(n_412), .Y(n_437) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
INVx1_ASAP7_75t_L g434 ( .A(n_426), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_428), .A2(n_432), .B1(n_435), .B2(n_437), .C(n_438), .Y(n_431) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
NAND4xp25_ASAP7_75t_SL g445 ( .A(n_446), .B(n_449), .C(n_453), .D(n_461), .Y(n_445) );
AND2x2_ASAP7_75t_L g459 ( .A(n_452), .B(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_467), .Y(n_795) );
AND2x2_ASAP7_75t_L g803 ( .A(n_467), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_670), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_618), .Y(n_471) );
OAI211xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_509), .B(n_538), .C(n_603), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_475), .A2(n_539), .B(n_754), .Y(n_753) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
INVx2_ASAP7_75t_L g599 ( .A(n_476), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_476), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g710 ( .A(n_477), .B(n_488), .Y(n_710) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g578 ( .A(n_478), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_478), .B(n_502), .Y(n_615) );
AND2x2_ASAP7_75t_L g648 ( .A(n_478), .B(n_565), .Y(n_648) );
OR2x2_ASAP7_75t_L g653 ( .A(n_478), .B(n_502), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_482), .A2(n_498), .B(n_499), .Y(n_497) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_482), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g563 ( .A(n_483), .Y(n_563) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g792 ( .A(n_487), .Y(n_792) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_501), .Y(n_487) );
AND2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_502), .Y(n_593) );
INVx3_ASAP7_75t_L g601 ( .A(n_488), .Y(n_601) );
NAND2x1p5_ASAP7_75t_SL g633 ( .A(n_488), .B(n_617), .Y(n_633) );
INVx1_ASAP7_75t_L g651 ( .A(n_488), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_488), .B(n_596), .Y(n_676) );
BUFx2_ASAP7_75t_L g762 ( .A(n_488), .Y(n_762) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_497), .B(n_500), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g546 ( .A(n_502), .Y(n_546) );
INVx1_ASAP7_75t_L g602 ( .A(n_502), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_502), .B(n_578), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_502), .B(n_565), .Y(n_711) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_526), .Y(n_509) );
INVx1_ASAP7_75t_L g769 ( .A(n_510), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
OR2x2_ASAP7_75t_L g541 ( .A(n_511), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g606 ( .A(n_511), .Y(n_606) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g585 ( .A(n_515), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_518), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_519), .A2(n_568), .B(n_574), .Y(n_567) );
INVx2_ASAP7_75t_L g542 ( .A(n_520), .Y(n_542) );
OR2x2_ASAP7_75t_L g607 ( .A(n_520), .B(n_527), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_520), .B(n_527), .Y(n_612) );
INVx2_ASAP7_75t_L g657 ( .A(n_520), .Y(n_657) );
AND2x2_ASAP7_75t_L g698 ( .A(n_520), .B(n_551), .Y(n_698) );
AND2x2_ASAP7_75t_L g732 ( .A(n_520), .B(n_629), .Y(n_732) );
INVx1_ASAP7_75t_L g543 ( .A(n_526), .Y(n_543) );
INVx1_ASAP7_75t_L g662 ( .A(n_526), .Y(n_662) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g582 ( .A(n_527), .B(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g623 ( .A(n_527), .B(n_584), .Y(n_623) );
INVx2_ASAP7_75t_L g629 ( .A(n_527), .Y(n_629) );
AND2x2_ASAP7_75t_L g684 ( .A(n_527), .B(n_551), .Y(n_684) );
AND2x2_ASAP7_75t_L g741 ( .A(n_527), .B(n_550), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_544), .B1(n_579), .B2(n_590), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_541), .B(n_720), .C(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g638 ( .A(n_542), .Y(n_638) );
AND2x2_ASAP7_75t_L g688 ( .A(n_542), .B(n_550), .Y(n_688) );
INVx1_ASAP7_75t_L g788 ( .A(n_543), .Y(n_788) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_545), .B(n_743), .Y(n_779) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g634 ( .A(n_546), .Y(n_634) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_564), .Y(n_548) );
INVx1_ASAP7_75t_L g622 ( .A(n_549), .Y(n_622) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g702 ( .A(n_550), .B(n_583), .Y(n_702) );
AND2x2_ASAP7_75t_L g721 ( .A(n_550), .B(n_628), .Y(n_721) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g589 ( .A(n_551), .Y(n_589) );
BUFx3_ASAP7_75t_L g627 ( .A(n_551), .Y(n_627) );
AND2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_657), .Y(n_656) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_559), .B(n_562), .Y(n_553) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g749 ( .A(n_564), .Y(n_749) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_578), .Y(n_564) );
INVx2_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .B(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g597 ( .A(n_578), .Y(n_597) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x6_ASAP7_75t_L g580 ( .A(n_581), .B(n_588), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g636 ( .A(n_582), .B(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g766 ( .A(n_582), .Y(n_766) );
INVx1_ASAP7_75t_L g611 ( .A(n_583), .Y(n_611) );
AND2x2_ASAP7_75t_L g691 ( .A(n_583), .B(n_629), .Y(n_691) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g628 ( .A(n_584), .B(n_629), .Y(n_628) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_589), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g724 ( .A(n_589), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_598), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_591), .A2(n_632), .B1(n_635), .B2(n_639), .Y(n_631) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_592), .A2(n_612), .B1(n_644), .B2(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
BUFx2_ASAP7_75t_SL g630 ( .A(n_593), .Y(n_630) );
AND2x4_ASAP7_75t_L g748 ( .A(n_593), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g757 ( .A(n_593), .Y(n_757) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g669 ( .A(n_595), .Y(n_669) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_596), .B(n_601), .Y(n_727) );
INVxp67_ASAP7_75t_L g756 ( .A(n_596), .Y(n_756) );
AND2x2_ASAP7_75t_L g761 ( .A(n_596), .B(n_627), .Y(n_761) );
OR2x2_ASAP7_75t_L g743 ( .A(n_597), .B(n_617), .Y(n_743) );
INVx1_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_599), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g663 ( .A(n_600), .B(n_648), .Y(n_663) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_601), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g647 ( .A(n_601), .Y(n_647) );
OR2x2_ASAP7_75t_L g742 ( .A(n_601), .B(n_743), .Y(n_742) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_613), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g660 ( .A(n_606), .B(n_657), .Y(n_660) );
INVx2_ASAP7_75t_L g784 ( .A(n_606), .Y(n_784) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g713 ( .A(n_610), .B(n_656), .Y(n_713) );
AND2x2_ASAP7_75t_L g738 ( .A(n_610), .B(n_684), .Y(n_738) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g641 ( .A(n_611), .Y(n_641) );
AND2x2_ASAP7_75t_L g668 ( .A(n_612), .B(n_622), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_612), .B(n_667), .Y(n_680) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g765 ( .A(n_615), .Y(n_765) );
OR2x2_ASAP7_75t_L g781 ( .A(n_615), .B(n_676), .Y(n_781) );
INVx1_ASAP7_75t_L g705 ( .A(n_617), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_642), .C(n_664), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_624), .B1(n_625), .B2(n_630), .C(n_631), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g644 ( .A(n_623), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_623), .B(n_688), .Y(n_772) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g667 ( .A(n_627), .Y(n_667) );
AND3x1_ASAP7_75t_L g763 ( .A(n_627), .B(n_764), .C(n_765), .Y(n_763) );
AND2x2_ASAP7_75t_L g750 ( .A(n_628), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g760 ( .A(n_628), .Y(n_760) );
INVxp67_ASAP7_75t_L g774 ( .A(n_630), .Y(n_774) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
OR2x2_ASAP7_75t_L g729 ( .A(n_633), .B(n_653), .Y(n_729) );
INVx2_ASAP7_75t_L g764 ( .A(n_633), .Y(n_764) );
INVx1_ASAP7_75t_L g682 ( .A(n_634), .Y(n_682) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_636), .A2(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_637), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g645 ( .A(n_638), .Y(n_645) );
OR2x2_ASAP7_75t_L g739 ( .A(n_638), .B(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g699 ( .A(n_641), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_641), .B(n_698), .Y(n_778) );
AND3x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_649), .C(n_654), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
AND2x2_ASAP7_75t_L g693 ( .A(n_645), .B(n_684), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_646), .A2(n_713), .B1(n_714), .B2(n_716), .Y(n_712) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
OAI321xp33_ASAP7_75t_L g735 ( .A1(n_647), .A2(n_736), .A3(n_737), .B1(n_739), .B2(n_742), .C(n_744), .Y(n_735) );
AND2x2_ASAP7_75t_L g787 ( .A(n_647), .B(n_652), .Y(n_787) );
AND2x2_ASAP7_75t_L g685 ( .A(n_648), .B(n_651), .Y(n_685) );
INVx2_ASAP7_75t_L g694 ( .A(n_650), .Y(n_694) );
AND2x2_ASAP7_75t_L g703 ( .A(n_650), .B(n_704), .Y(n_703) );
AND2x4_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g715 ( .A(n_653), .B(n_705), .Y(n_715) );
INVx2_ASAP7_75t_L g747 ( .A(n_653), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B(n_663), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g751 ( .A(n_657), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_660), .B(n_667), .Y(n_677) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B(n_669), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_667), .B(n_691), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_667), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g768 ( .A(n_667), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g736 ( .A(n_669), .Y(n_736) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_671), .B(n_733), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_695), .C(n_718), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_686), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B1(n_678), .B2(n_681), .C(n_683), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OR2x2_ASAP7_75t_L g726 ( .A(n_675), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_692), .B(n_694), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g723 ( .A(n_691), .B(n_724), .Y(n_723) );
OAI21xp33_ASAP7_75t_SL g706 ( .A1(n_692), .A2(n_707), .B(n_712), .Y(n_706) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_700), .B(n_703), .C(n_706), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_697), .B(n_772), .Y(n_771) );
NAND2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_705), .B(n_747), .Y(n_746) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_708), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_725), .B1(n_728), .B2(n_730), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_727), .Y(n_790) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_770), .C(n_785), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_752), .Y(n_734) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B(n_750), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_758), .C(n_767), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
AOI32xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_761), .A3(n_762), .B1(n_763), .B2(n_766), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g786 ( .A(n_761), .B(n_787), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_773), .B(n_775), .Y(n_770) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AOI22x1_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B1(n_780), .B2(n_782), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AOI21xp33_ASAP7_75t_L g789 ( .A1(n_778), .A2(n_790), .B(n_791), .Y(n_789) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .B(n_789), .Y(n_785) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx8_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
BUFx12f_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
BUFx10_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR2x1_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
BUFx3_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx8_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_808), .B(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_809), .A2(n_821), .B1(n_834), .B2(n_844), .Y(n_833) );
NOR2x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_822), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_817), .Y(n_810) );
BUFx12f_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx12f_ASAP7_75t_L g824 ( .A(n_812), .Y(n_824) );
INVx4_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx5_ASAP7_75t_L g832 ( .A(n_813), .Y(n_832) );
INVx3_ASAP7_75t_L g843 ( .A(n_813), .Y(n_843) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_832), .Y(n_829) );
INVx2_ASAP7_75t_SL g842 ( .A(n_830), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx8_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
OR2x6_ASAP7_75t_L g838 ( .A(n_839), .B(n_843), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OR2x4_ASAP7_75t_L g846 ( .A(n_841), .B(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx4_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
BUFx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
endmodule