module fake_netlist_5_1310_n_1152 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1152);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1152;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_1104;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1020;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_897;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_1064;
wire n_858;
wire n_829;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_1069;
wire n_969;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_1058;
wire n_358;
wire n_838;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_1116;
wire n_627;
wire n_954;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_707;
wire n_710;
wire n_857;
wire n_695;
wire n_795;
wire n_832;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_1004;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1032;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_132),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_162),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_24),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_66),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_189),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_51),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_68),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_122),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_34),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_26),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_63),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_124),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_109),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_136),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_106),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_203),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_119),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_140),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_170),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_152),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_9),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_158),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_91),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_47),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_84),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_23),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_141),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_175),
.Y(n_253)
);

INVxp33_ASAP7_75t_R g254 ( 
.A(n_39),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_144),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_102),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_217),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_32),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_52),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_183),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_147),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_107),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_77),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_74),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_138),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_182),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_23),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_31),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_108),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_94),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_115),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_155),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_116),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_173),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_101),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_156),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_37),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_199),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_12),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_213),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_10),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_50),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_290),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_222),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_239),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_266),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_246),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_251),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_237),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_247),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_0),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_261),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_261),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_219),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_220),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_221),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_223),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_224),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_257),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_225),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_226),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_228),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_234),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_318),
.Y(n_341)
);

OA21x2_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_313),
.B(n_329),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_235),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_233),
.B(n_229),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_274),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_236),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_240),
.Y(n_347)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_241),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g363 ( 
.A1(n_298),
.A2(n_301),
.B(n_300),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_276),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_319),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_305),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_320),
.B(n_282),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_291),
.A2(n_285),
.B1(n_288),
.B2(n_283),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_242),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_337),
.Y(n_373)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_302),
.A2(n_244),
.B(n_243),
.Y(n_374)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_302),
.A2(n_249),
.B(n_248),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_307),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_310),
.B(n_252),
.Y(n_384)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_304),
.A2(n_280),
.B1(n_273),
.B2(n_272),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_309),
.A2(n_255),
.B(n_253),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_338),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_311),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_292),
.A2(n_268),
.B1(n_267),
.B2(n_265),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_390),
.B(n_391),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_369),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_336),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_388),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_390),
.B(n_315),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_345),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_343),
.B(n_336),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_341),
.Y(n_411)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_390),
.B(n_315),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_341),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_390),
.B(n_316),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_391),
.B(n_316),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_366),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_384),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_323),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_384),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_325),
.Y(n_432)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_346),
.B(n_295),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_346),
.Y(n_440)
);

CKINVDCx6p67_ASAP7_75t_R g441 ( 
.A(n_394),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

AOI21x1_ASAP7_75t_L g443 ( 
.A1(n_363),
.A2(n_376),
.B(n_374),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_345),
.B(n_256),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_349),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_368),
.B(n_364),
.Y(n_448)
);

NOR2x1p5_ASAP7_75t_L g449 ( 
.A(n_394),
.B(n_254),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_363),
.A2(n_259),
.B(n_258),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_356),
.B(n_335),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_346),
.B(n_262),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_358),
.B(n_264),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_354),
.Y(n_457)
);

INVxp67_ASAP7_75t_R g458 ( 
.A(n_344),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_368),
.A2(n_392),
.B1(n_387),
.B2(n_345),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_379),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_364),
.B(n_263),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_394),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_459),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_411),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_422),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_438),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_439),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_442),
.B(n_394),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_400),
.B(n_356),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_367),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_365),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_386),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_345),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_428),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_428),
.B(n_387),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_407),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_396),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_452),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_401),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_434),
.B(n_350),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_441),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_455),
.B(n_345),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_441),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_387),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_352),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_382),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_398),
.B(n_365),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_454),
.B(n_456),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_414),
.B(n_374),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_395),
.B(n_347),
.Y(n_520)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_443),
.A2(n_376),
.B(n_374),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_404),
.B(n_358),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_417),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_448),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_418),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_418),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_449),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_420),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_420),
.B(n_376),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_421),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_451),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_404),
.B(n_358),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_398),
.B(n_375),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_415),
.B(n_347),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_450),
.A2(n_409),
.B(n_344),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVxp33_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_430),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_415),
.B(n_375),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_430),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_463),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

XNOR2x2_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_348),
.Y(n_552)
);

INVx8_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_469),
.B(n_424),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_494),
.B(n_448),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_488),
.A2(n_458),
.B1(n_444),
.B2(n_419),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_479),
.Y(n_558)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_472),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_495),
.B(n_419),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_524),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_490),
.A2(n_419),
.B1(n_433),
.B2(n_370),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_375),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_482),
.B(n_385),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_472),
.B(n_370),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_528),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_484),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_511),
.A2(n_370),
.B1(n_347),
.B2(n_460),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_518),
.Y(n_572)
);

NOR2x1p5_ASAP7_75t_L g573 ( 
.A(n_515),
.B(n_348),
.Y(n_573)
);

NOR3xp33_ASAP7_75t_SL g574 ( 
.A(n_536),
.B(n_389),
.C(n_348),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_491),
.B(n_405),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_485),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_481),
.B(n_457),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_491),
.B(n_405),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_499),
.B(n_385),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_511),
.B(n_405),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_516),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_502),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_486),
.B(n_385),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_385),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_552),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_496),
.B(n_447),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_498),
.B(n_447),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_509),
.B(n_389),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_427),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_503),
.B(n_379),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_531),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_501),
.B(n_427),
.Y(n_592)
);

NOR2x2_ASAP7_75t_L g593 ( 
.A(n_517),
.B(n_389),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_549),
.B(n_427),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_509),
.B(n_433),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_507),
.B(n_435),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_512),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_477),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_510),
.B(n_383),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_435),
.Y(n_601)
);

A2O1A1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_545),
.A2(n_437),
.B(n_435),
.C(n_453),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_489),
.B(n_437),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_489),
.B(n_437),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_523),
.B(n_355),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_493),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_471),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_537),
.B(n_355),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_504),
.B(n_457),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_505),
.B(n_379),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_528),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_513),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_522),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_542),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_508),
.B(n_453),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_517),
.B(n_355),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_546),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_508),
.A2(n_383),
.B(n_453),
.C(n_460),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_527),
.A2(n_465),
.B1(n_462),
.B2(n_399),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_520),
.B(n_525),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_562),
.B(n_487),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_SL g624 ( 
.A(n_585),
.B(n_474),
.C(n_473),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_SL g625 ( 
.A(n_565),
.B(n_476),
.C(n_475),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_554),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_569),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_R g628 ( 
.A(n_572),
.B(n_478),
.Y(n_628)
);

AND2x6_ASAP7_75t_SL g629 ( 
.A(n_588),
.B(n_470),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_581),
.B(n_520),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_611),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_591),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_555),
.B(n_584),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_570),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_597),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_SL g636 ( 
.A(n_595),
.B(n_550),
.C(n_540),
.Y(n_636)
);

AND2x6_ASAP7_75t_SL g637 ( 
.A(n_579),
.B(n_551),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_583),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_577),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_600),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_598),
.Y(n_642)
);

NOR3xp33_ASAP7_75t_SL g643 ( 
.A(n_566),
.B(n_540),
.C(n_533),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_555),
.B(n_529),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_612),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_R g646 ( 
.A(n_559),
.B(n_526),
.Y(n_646)
);

AND3x2_ASAP7_75t_SL g647 ( 
.A(n_593),
.B(n_465),
.C(n_462),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_567),
.B(n_355),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_561),
.A2(n_553),
.B(n_533),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_607),
.B(n_526),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_571),
.A2(n_519),
.B1(n_553),
.B2(n_547),
.Y(n_651)
);

BUFx5_ASAP7_75t_L g652 ( 
.A(n_586),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_559),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_SL g654 ( 
.A(n_590),
.B(n_519),
.C(n_530),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_613),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_617),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_R g657 ( 
.A(n_582),
.B(n_521),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_586),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_558),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_SL g660 ( 
.A(n_605),
.B(n_548),
.C(n_534),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_557),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_564),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_621),
.B(n_532),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_557),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_568),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_621),
.B(n_535),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_573),
.B(n_541),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_576),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_568),
.B(n_544),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_599),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_606),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_614),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_601),
.B(n_497),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_SL g674 ( 
.A(n_574),
.B(n_399),
.C(n_1),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_596),
.B(n_601),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_594),
.B(n_497),
.Y(n_677)
);

INVx3_ASAP7_75t_SL g678 ( 
.A(n_610),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_575),
.B(n_497),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_594),
.B(n_497),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_615),
.Y(n_681)
);

BUFx4f_ASAP7_75t_L g682 ( 
.A(n_586),
.Y(n_682)
);

AOI22x1_ASAP7_75t_L g683 ( 
.A1(n_618),
.A2(n_399),
.B1(n_446),
.B2(n_423),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_608),
.B(n_379),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_589),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_620),
.B(n_497),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_586),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_633),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_633),
.A2(n_556),
.B(n_580),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_638),
.B(n_609),
.Y(n_690)
);

O2A1O1Ixp5_ASAP7_75t_L g691 ( 
.A1(n_649),
.A2(n_563),
.B(n_602),
.C(n_578),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_683),
.A2(n_619),
.B(n_604),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_643),
.A2(n_604),
.B(n_603),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_642),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_626),
.B(n_592),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_686),
.B(n_563),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_673),
.A2(n_616),
.B(n_603),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_679),
.A2(n_561),
.B(n_616),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_623),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_673),
.A2(n_587),
.B(n_446),
.Y(n_700)
);

NOR2x1_ASAP7_75t_L g701 ( 
.A(n_632),
.B(n_423),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_651),
.A2(n_587),
.B(n_446),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_651),
.A2(n_587),
.B(n_446),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_631),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_645),
.Y(n_705)
);

OAI21x1_ASAP7_75t_SL g706 ( 
.A1(n_644),
.A2(n_587),
.B(n_29),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_656),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_675),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_708)
);

AOI21x1_ASAP7_75t_L g709 ( 
.A1(n_677),
.A2(n_423),
.B(n_412),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_631),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_646),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_666),
.A2(n_412),
.B(n_423),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_655),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_622),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_631),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_662),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_639),
.B(n_2),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_641),
.B(n_28),
.Y(n_718)
);

OAI21x1_ASAP7_75t_L g719 ( 
.A1(n_677),
.A2(n_412),
.B(n_35),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_661),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_681),
.B(n_4),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_667),
.Y(n_722)
);

AOI221xp5_ASAP7_75t_L g723 ( 
.A1(n_624),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_636),
.A2(n_412),
.B(n_36),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_668),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_670),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_676),
.B(n_5),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_661),
.Y(n_729)
);

AO21x1_ASAP7_75t_L g730 ( 
.A1(n_680),
.A2(n_6),
.B(n_7),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_681),
.B(n_8),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_680),
.A2(n_412),
.B(n_38),
.Y(n_733)
);

O2A1O1Ixp5_ASAP7_75t_L g734 ( 
.A1(n_682),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_644),
.A2(n_40),
.B(n_33),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_630),
.B(n_11),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_638),
.B(n_13),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_663),
.A2(n_42),
.B(n_41),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_659),
.B(n_13),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_652),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_652),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_640),
.B(n_14),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_640),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_684),
.A2(n_44),
.B(n_43),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_627),
.B(n_14),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_634),
.B(n_15),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_637),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_685),
.B(n_15),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_664),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_696),
.A2(n_682),
.B(n_658),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_694),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_696),
.A2(n_658),
.B(n_648),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_SL g753 ( 
.A1(n_723),
.A2(n_674),
.B(n_629),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_708),
.A2(n_625),
.B(n_678),
.C(n_660),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_745),
.B(n_635),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_712),
.A2(n_658),
.B(n_669),
.Y(n_756)
);

BUFx4f_ASAP7_75t_L g757 ( 
.A(n_729),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_747),
.A2(n_653),
.B1(n_650),
.B2(n_671),
.Y(n_758)
);

AO21x1_ASAP7_75t_L g759 ( 
.A1(n_688),
.A2(n_669),
.B(n_650),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_688),
.B(n_672),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_695),
.B(n_629),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_SL g762 ( 
.A1(n_708),
.A2(n_647),
.B(n_665),
.C(n_628),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_689),
.A2(n_698),
.B(n_691),
.Y(n_764)
);

AO32x2_ASAP7_75t_L g765 ( 
.A1(n_730),
.A2(n_637),
.A3(n_654),
.B1(n_657),
.B2(n_652),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_746),
.B(n_664),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_SL g767 ( 
.A1(n_738),
.A2(n_665),
.B(n_652),
.C(n_687),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_724),
.A2(n_664),
.B(n_17),
.C(n_18),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_709),
.A2(n_46),
.B(n_45),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_SL g770 ( 
.A1(n_748),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_694),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_705),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_690),
.B(n_722),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_714),
.B(n_48),
.Y(n_774)
);

AOI21x1_ASAP7_75t_L g775 ( 
.A1(n_702),
.A2(n_703),
.B(n_692),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_715),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_749),
.B(n_715),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_700),
.A2(n_692),
.B(n_702),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_713),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_726),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_693),
.A2(n_16),
.B(n_19),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_717),
.B(n_19),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_713),
.B(n_20),
.Y(n_783)
);

AO32x2_ASAP7_75t_L g784 ( 
.A1(n_734),
.A2(n_21),
.A3(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_699),
.Y(n_785)
);

AO31x2_ASAP7_75t_L g786 ( 
.A1(n_728),
.A2(n_133),
.A3(n_216),
.B(n_215),
.Y(n_786)
);

OAI22x1_ASAP7_75t_L g787 ( 
.A1(n_721),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_749),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_703),
.A2(n_134),
.B(n_214),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_719),
.A2(n_131),
.B(n_212),
.Y(n_790)
);

AO31x2_ASAP7_75t_L g791 ( 
.A1(n_728),
.A2(n_130),
.A3(n_211),
.B(n_49),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_716),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_719),
.A2(n_135),
.B(n_210),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_735),
.A2(n_26),
.B(n_27),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_697),
.A2(n_218),
.B(n_53),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_697),
.A2(n_209),
.B(n_54),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_727),
.B(n_27),
.Y(n_797)
);

AO31x2_ASAP7_75t_L g798 ( 
.A1(n_740),
.A2(n_55),
.A3(n_56),
.B(n_57),
.Y(n_798)
);

INVx8_ASAP7_75t_L g799 ( 
.A(n_729),
.Y(n_799)
);

AO21x1_ASAP7_75t_L g800 ( 
.A1(n_737),
.A2(n_58),
.B(n_59),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_744),
.A2(n_208),
.B(n_61),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_740),
.A2(n_741),
.B(n_690),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_733),
.A2(n_60),
.B(n_64),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_711),
.Y(n_804)
);

BUFx4f_ASAP7_75t_L g805 ( 
.A(n_729),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_721),
.B(n_207),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_732),
.A2(n_65),
.B(n_67),
.C(n_69),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_SL g808 ( 
.A1(n_742),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_718),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_736),
.A2(n_739),
.B(n_725),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_690),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_741),
.A2(n_81),
.B(n_82),
.Y(n_812)
);

AOI211x1_ASAP7_75t_L g813 ( 
.A1(n_743),
.A2(n_83),
.B(n_86),
.C(n_87),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_733),
.A2(n_88),
.B(n_89),
.Y(n_814)
);

OA21x2_ASAP7_75t_L g815 ( 
.A1(n_706),
.A2(n_743),
.B(n_707),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_731),
.A2(n_205),
.B(n_93),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_701),
.A2(n_92),
.B(n_95),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_704),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_714),
.B(n_204),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_710),
.B(n_96),
.Y(n_820)
);

CKINVDCx11_ASAP7_75t_R g821 ( 
.A(n_804),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_780),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_799),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_781),
.A2(n_794),
.B1(n_806),
.B2(n_810),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_787),
.A2(n_720),
.B1(n_731),
.B2(n_99),
.Y(n_825)
);

INVx6_ASAP7_75t_L g826 ( 
.A(n_763),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_761),
.A2(n_720),
.B1(n_731),
.B2(n_100),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_751),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_763),
.B(n_731),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_792),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_772),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_785),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_777),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_776),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_771),
.Y(n_835)
);

BUFx4f_ASAP7_75t_SL g836 ( 
.A(n_788),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_753),
.A2(n_97),
.B1(n_98),
.B2(n_103),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_799),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_760),
.B(n_104),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_768),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_779),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_783),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_797),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_843)
);

INVx4_ASAP7_75t_SL g844 ( 
.A(n_782),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_818),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_759),
.Y(n_846)
);

CKINVDCx11_ASAP7_75t_R g847 ( 
.A(n_774),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_755),
.Y(n_848)
);

INVx6_ASAP7_75t_L g849 ( 
.A(n_763),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_784),
.Y(n_850)
);

BUFx2_ASAP7_75t_SL g851 ( 
.A(n_766),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_758),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_802),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_800),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_764),
.A2(n_127),
.B(n_128),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_SL g856 ( 
.A1(n_801),
.A2(n_129),
.B1(n_137),
.B2(n_139),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_784),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_815),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_765),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_773),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_820),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_813),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_757),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_805),
.Y(n_865)
);

OAI22xp33_ASAP7_75t_L g866 ( 
.A1(n_819),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_765),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_754),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_765),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_786),
.Y(n_870)
);

AOI22x1_ASAP7_75t_SL g871 ( 
.A1(n_762),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_817),
.Y(n_872)
);

OAI22xp33_ASAP7_75t_L g873 ( 
.A1(n_750),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

BUFx2_ASAP7_75t_SL g875 ( 
.A(n_756),
.Y(n_875)
);

INVx8_ASAP7_75t_L g876 ( 
.A(n_811),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_808),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_809),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_816),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_752),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_786),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_791),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_830),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_870),
.B(n_778),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_860),
.B(n_775),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_828),
.Y(n_886)
);

CKINVDCx6p67_ASAP7_75t_R g887 ( 
.A(n_821),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_835),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_882),
.A2(n_814),
.B(n_803),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_858),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_882),
.A2(n_793),
.B(n_790),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_841),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_855),
.A2(n_769),
.B(n_789),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_859),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_846),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_831),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_848),
.B(n_767),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_867),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_869),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_868),
.A2(n_876),
.B1(n_824),
.B2(n_840),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_848),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_853),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_881),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_850),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_842),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_857),
.Y(n_906)
);

CKINVDCx11_ASAP7_75t_R g907 ( 
.A(n_847),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_833),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_837),
.A2(n_807),
.B1(n_812),
.B2(n_796),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_875),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_872),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_862),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_826),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_874),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_874),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_839),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_855),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_861),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_845),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_851),
.B(n_791),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_868),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_877),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_834),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_844),
.B(n_798),
.Y(n_924)
);

AO31x2_ASAP7_75t_L g925 ( 
.A1(n_863),
.A2(n_795),
.A3(n_840),
.B(n_878),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_826),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_849),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_849),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_906),
.B(n_844),
.Y(n_929)
);

AO21x2_ASAP7_75t_L g930 ( 
.A1(n_917),
.A2(n_863),
.B(n_837),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_894),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_894),
.Y(n_932)
);

OA21x2_ASAP7_75t_L g933 ( 
.A1(n_893),
.A2(n_854),
.B(n_879),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_921),
.Y(n_934)
);

AO21x1_ASAP7_75t_SL g935 ( 
.A1(n_917),
.A2(n_825),
.B(n_827),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_890),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_890),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_900),
.A2(n_876),
.B1(n_878),
.B2(n_852),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_884),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_883),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_906),
.B(n_822),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_883),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_889),
.A2(n_852),
.B(n_880),
.Y(n_943)
);

AO21x2_ASAP7_75t_L g944 ( 
.A1(n_889),
.A2(n_866),
.B(n_873),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_898),
.Y(n_945)
);

AO21x2_ASAP7_75t_L g946 ( 
.A1(n_891),
.A2(n_832),
.B(n_876),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_904),
.B(n_885),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_888),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_898),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_899),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_899),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_886),
.B(n_836),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_892),
.Y(n_953)
);

AO21x2_ASAP7_75t_L g954 ( 
.A1(n_891),
.A2(n_871),
.B(n_798),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_926),
.Y(n_955)
);

INVx4_ASAP7_75t_SL g956 ( 
.A(n_925),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_887),
.B(n_823),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_931),
.Y(n_958)
);

NOR4xp25_ASAP7_75t_SL g959 ( 
.A(n_936),
.B(n_915),
.C(n_914),
.D(n_895),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_939),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_939),
.B(n_895),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_931),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_939),
.B(n_904),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_939),
.B(n_956),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_946),
.A2(n_903),
.B(n_911),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_932),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_956),
.B(n_885),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_902),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_932),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_956),
.B(n_896),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_934),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_938),
.A2(n_909),
.B1(n_921),
.B2(n_916),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_945),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_941),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_930),
.A2(n_916),
.B1(n_856),
.B2(n_910),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_936),
.B(n_901),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_941),
.B(n_905),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_934),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_945),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_949),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_963),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_956),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_967),
.B(n_956),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_958),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_974),
.B(n_929),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_971),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_964),
.B(n_947),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_968),
.B(n_937),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_971),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_964),
.B(n_934),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_973),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_979),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_958),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_963),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_960),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_961),
.B(n_978),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_990),
.B(n_970),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_986),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_992),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_985),
.B(n_977),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_991),
.B(n_970),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_987),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_993),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_989),
.B(n_976),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_989),
.B(n_979),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_981),
.Y(n_1007)
);

NAND2xp67_ASAP7_75t_L g1008 ( 
.A(n_982),
.B(n_952),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_990),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1002),
.B(n_997),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1003),
.B(n_995),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_998),
.Y(n_1013)
);

AND2x4_ASAP7_75t_SL g1014 ( 
.A(n_998),
.B(n_887),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_1009),
.B(n_997),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_999),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1007),
.B(n_991),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1015),
.Y(n_1018)
);

OAI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_1013),
.A2(n_1005),
.B1(n_1001),
.B2(n_996),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_1014),
.A2(n_1017),
.B1(n_1010),
.B2(n_1012),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_1014),
.B(n_907),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_1011),
.B(n_922),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1018),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1022),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1020),
.B(n_1012),
.Y(n_1026)
);

CKINVDCx16_ASAP7_75t_R g1027 ( 
.A(n_1021),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_1023),
.B(n_1016),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_1019),
.B(n_957),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1018),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1018),
.B(n_1000),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1020),
.A2(n_930),
.B1(n_922),
.B2(n_972),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_1025),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1033),
.A2(n_975),
.B(n_915),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1030),
.A2(n_996),
.B1(n_914),
.B2(n_1006),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1024),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1029),
.B(n_988),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1028),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1031),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1032),
.A2(n_930),
.B1(n_983),
.B2(n_982),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_1034),
.B(n_919),
.C(n_923),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1039),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1040),
.B(n_1006),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_1037),
.B(n_984),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1038),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_SL g1047 ( 
.A1(n_1035),
.A2(n_983),
.B(n_918),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_1041),
.B(n_976),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1036),
.B(n_988),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1047),
.A2(n_996),
.B(n_943),
.C(n_971),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1046),
.B(n_996),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_1043),
.A2(n_1049),
.B1(n_1048),
.B2(n_1044),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1045),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1042),
.B(n_984),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_1042),
.A2(n_930),
.B1(n_996),
.B2(n_955),
.Y(n_1055)
);

OAI321xp33_ASAP7_75t_L g1056 ( 
.A1(n_1043),
.A2(n_913),
.A3(n_918),
.B1(n_843),
.B2(n_910),
.C(n_927),
.Y(n_1056)
);

INVxp33_ASAP7_75t_L g1057 ( 
.A(n_1051),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1053),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1054),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1052),
.B(n_994),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1055),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1056),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1050),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1053),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1053),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1053),
.Y(n_1067)
);

XNOR2x2_ASAP7_75t_L g1068 ( 
.A(n_1065),
.B(n_959),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1062),
.A2(n_935),
.B1(n_944),
.B2(n_933),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_1060),
.B(n_968),
.Y(n_1070)
);

NOR3x1_ASAP7_75t_L g1071 ( 
.A(n_1062),
.B(n_865),
.C(n_913),
.Y(n_1071)
);

OAI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_1063),
.A2(n_959),
.B(n_864),
.C(n_955),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1058),
.B(n_994),
.Y(n_1073)
);

AOI211x1_ASAP7_75t_L g1074 ( 
.A1(n_1066),
.A2(n_1067),
.B(n_1059),
.C(n_1057),
.Y(n_1074)
);

NOR4xp75_ASAP7_75t_L g1075 ( 
.A(n_1064),
.B(n_1061),
.C(n_978),
.D(n_960),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1058),
.B(n_980),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1058),
.Y(n_1077)
);

NAND4xp75_ASAP7_75t_L g1078 ( 
.A(n_1065),
.B(n_929),
.C(n_927),
.D(n_924),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_905),
.Y(n_1079)
);

OAI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1074),
.A2(n_864),
.B(n_955),
.C(n_838),
.Y(n_1080)
);

NAND5xp2_ASAP7_75t_L g1081 ( 
.A(n_1073),
.B(n_829),
.C(n_924),
.D(n_935),
.E(n_902),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_L g1082 ( 
.A(n_1076),
.B(n_955),
.C(n_838),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1072),
.A2(n_944),
.B(n_864),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_1070),
.B(n_168),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1069),
.A2(n_944),
.B1(n_946),
.B2(n_960),
.C(n_928),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_1078),
.B(n_928),
.C(n_943),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1084),
.B(n_1071),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1080),
.Y(n_1088)
);

AOI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1082),
.A2(n_1075),
.B(n_1068),
.C(n_926),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1079),
.B(n_946),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_SL g1091 ( 
.A(n_1083),
.B(n_897),
.C(n_961),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_1081),
.B(n_911),
.C(n_912),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1086),
.B(n_926),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1085),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1084),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_L g1096 ( 
.A(n_1095),
.B(n_960),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1088),
.Y(n_1097)
);

OAI32xp33_ASAP7_75t_L g1098 ( 
.A1(n_1094),
.A2(n_1093),
.A3(n_1090),
.B1(n_1092),
.B2(n_1089),
.Y(n_1098)
);

XOR2x1_ASAP7_75t_L g1099 ( 
.A(n_1087),
.B(n_933),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1091),
.B(n_912),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_SL g1101 ( 
.A(n_1089),
.B(n_937),
.C(n_980),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1095),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1095),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1095),
.B(n_926),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1087),
.A2(n_944),
.B(n_933),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_1097),
.B(n_926),
.C(n_908),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1102),
.A2(n_933),
.B1(n_908),
.B2(n_962),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_1098),
.B(n_169),
.C(n_171),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1104),
.B(n_908),
.Y(n_1109)
);

NOR2x1_ASAP7_75t_L g1110 ( 
.A(n_1103),
.B(n_965),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1096),
.B(n_966),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_L g1112 ( 
.A(n_1101),
.B(n_893),
.C(n_174),
.Y(n_1112)
);

XNOR2xp5_ASAP7_75t_L g1113 ( 
.A(n_1099),
.B(n_172),
.Y(n_1113)
);

AND4x1_ASAP7_75t_L g1114 ( 
.A(n_1105),
.B(n_176),
.C(n_177),
.D(n_178),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1100),
.B(n_965),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1097),
.Y(n_1116)
);

NOR2x2_ASAP7_75t_L g1117 ( 
.A(n_1102),
.B(n_179),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1097),
.B(n_965),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1113),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1116),
.B(n_965),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1109),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1112),
.A2(n_966),
.B1(n_962),
.B2(n_958),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1117),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1111),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1106),
.A2(n_969),
.B1(n_966),
.B2(n_962),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1118),
.Y(n_1126)
);

AND4x1_ASAP7_75t_L g1127 ( 
.A(n_1108),
.B(n_180),
.C(n_181),
.D(n_184),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1123),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1121),
.A2(n_1115),
.B1(n_1110),
.B2(n_1107),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1119),
.A2(n_1114),
.B1(n_969),
.B2(n_951),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1124),
.A2(n_969),
.B1(n_954),
.B2(n_953),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1120),
.A2(n_954),
.B1(n_953),
.B2(n_920),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1122),
.A2(n_951),
.B1(n_950),
.B2(n_949),
.Y(n_1133)
);

OAI22x1_ASAP7_75t_L g1134 ( 
.A1(n_1127),
.A2(n_920),
.B1(n_950),
.B2(n_903),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1128),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1129),
.Y(n_1136)
);

XNOR2xp5_ASAP7_75t_L g1137 ( 
.A(n_1134),
.B(n_1126),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1138),
.Y(n_1139)
);

AOI22x1_ASAP7_75t_L g1140 ( 
.A1(n_1139),
.A2(n_1136),
.B1(n_1137),
.B2(n_1126),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1140),
.A2(n_1130),
.B1(n_1133),
.B2(n_1132),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1140),
.A2(n_1131),
.B1(n_1125),
.B2(n_942),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1140),
.A2(n_942),
.B1(n_940),
.B2(n_948),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_1141),
.B(n_185),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1142),
.B(n_186),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1143),
.A2(n_187),
.B(n_188),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_190),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1145),
.A2(n_191),
.B(n_192),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_193),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1147),
.A2(n_954),
.B1(n_194),
.B2(n_195),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1149),
.A2(n_954),
.B1(n_197),
.B2(n_198),
.Y(n_1151)
);

AOI211xp5_ASAP7_75t_L g1152 ( 
.A1(n_1150),
.A2(n_1148),
.B(n_1151),
.C(n_200),
.Y(n_1152)
);


endmodule