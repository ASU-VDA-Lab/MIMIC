module fake_jpeg_3223_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx3_ASAP7_75t_SL g44 ( 
.A(n_19),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_11),
.B(n_34),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_61),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_43),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_47),
.B1(n_43),
.B2(n_52),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_53),
.B1(n_50),
.B2(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_54),
.B1(n_40),
.B2(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_0),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_55),
.B1(n_59),
.B2(n_41),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_86),
.B1(n_60),
.B2(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_47),
.B1(n_38),
.B2(n_52),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_57),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_64),
.B(n_71),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_21),
.B(n_18),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_68),
.B1(n_67),
.B2(n_73),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_7),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_68),
.B1(n_73),
.B2(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_60),
.B1(n_45),
.B2(n_2),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_17),
.B1(n_16),
.B2(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_3),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_29),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_110),
.C(n_119),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_24),
.C(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_15),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_4),
.C(n_6),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_120),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_102),
.B(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_130),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_7),
.C(n_9),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_128),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_9),
.B(n_10),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_119),
.B1(n_112),
.B2(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_138),
.Y(n_143)
);

OAI321xp33_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_114),
.A3(n_117),
.B1(n_15),
.B2(n_13),
.C(n_14),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_142),
.A2(n_140),
.B1(n_122),
.B2(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_144),
.B(n_145),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_137),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_127),
.B(n_126),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_125),
.B(n_123),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_125),
.Y(n_151)
);


endmodule