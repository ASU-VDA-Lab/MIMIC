module fake_jpeg_1256_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_R g14 ( 
.A(n_7),
.B(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVxp33_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_6),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_12),
.B(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_11),
.B1(n_12),
.B2(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_14),
.B(n_16),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_11),
.B(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_18),
.B1(n_19),
.B2(n_3),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_5),
.Y(n_40)
);

NOR4xp25_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_27),
.C(n_28),
.D(n_31),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_39),
.C(n_40),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_37),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_37),
.B(n_43),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B(n_28),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_38),
.B(n_35),
.Y(n_55)
);


endmodule