module real_aes_10088_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_2086, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_2086;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_2043;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_2014;
wire n_1279;
wire n_2003;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_2035;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_2031;
wire n_1160;
wire n_2040;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_2049;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_1987;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_2063;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_2004;
wire n_1201;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_2067;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_2064;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_2082;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_2038;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_2041;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_2058;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_2068;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_2057;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_2050;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_2012;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_1712;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_2069;
wire n_1568;
wire n_1368;
wire n_994;
wire n_2059;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2045;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_2036;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_2072;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_2033;
wire n_1985;
wire n_1812;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_2061;
wire n_1163;
wire n_1278;
wire n_2039;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_2023;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_2081;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_2052;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_2070;
wire n_862;
wire n_869;
wire n_2019;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_2042;
wire n_1066;
wire n_2046;
wire n_2080;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_2062;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_2084;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_2065;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_936;
wire n_581;
wire n_2048;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_2032;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_2078;
wire n_377;
wire n_1169;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_2053;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_2034;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_2060;
wire n_1710;
wire n_2074;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_2066;
wire n_1156;
wire n_988;
wire n_2011;
wire n_2055;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1691;
wire n_1176;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_2079;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_2037;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_2030;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_2076;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_2044;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_2075;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1277;
wire n_1049;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_2047;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_2056;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_2083;
wire n_1963;
wire n_1958;
wire n_969;
wire n_2010;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_2077;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_2071;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_2051;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_2073;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_2054;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_0), .Y(n_716) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1), .Y(n_1697) );
OA22x2_ASAP7_75t_L g1115 ( .A1(n_2), .A2(n_1116), .B1(n_1172), .B2(n_1173), .Y(n_1115) );
INVxp67_ASAP7_75t_SL g1173 ( .A(n_2), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1726 ( .A1(n_3), .A2(n_362), .B1(n_1727), .B2(n_1735), .Y(n_1726) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_4), .Y(n_1261) );
INVx1_ASAP7_75t_L g755 ( .A(n_5), .Y(n_755) );
INVx1_ASAP7_75t_L g1262 ( .A(n_6), .Y(n_1262) );
INVx1_ASAP7_75t_L g1639 ( .A(n_7), .Y(n_1639) );
OAI221xp5_ASAP7_75t_L g1685 ( .A1(n_8), .A2(n_340), .B1(n_591), .B2(n_596), .C(n_889), .Y(n_1685) );
OAI22xp33_ASAP7_75t_SL g1706 ( .A1(n_8), .A2(n_340), .B1(n_670), .B2(n_672), .Y(n_1706) );
INVx1_ASAP7_75t_L g894 ( .A(n_9), .Y(n_894) );
AOI221xp5_ASAP7_75t_SL g919 ( .A1(n_9), .A2(n_150), .B1(n_653), .B2(n_920), .C(n_922), .Y(n_919) );
INVxp33_ASAP7_75t_L g1403 ( .A(n_10), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_10), .A2(n_104), .B1(n_1472), .B2(n_1473), .Y(n_1483) );
INVx1_ASAP7_75t_L g887 ( .A(n_11), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_11), .A2(n_241), .B1(n_934), .B2(n_936), .C(n_937), .Y(n_933) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_12), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_12), .A2(n_334), .B1(n_742), .B2(n_744), .Y(n_741) );
INVxp33_ASAP7_75t_L g1681 ( .A(n_13), .Y(n_1681) );
AOI221xp5_ASAP7_75t_L g1702 ( .A1(n_13), .A2(n_103), .B1(n_665), .B2(n_743), .C(n_1703), .Y(n_1702) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_14), .A2(n_100), .B1(n_665), .B2(n_1252), .C(n_1253), .Y(n_1251) );
INVx1_ASAP7_75t_L g1269 ( .A(n_14), .Y(n_1269) );
INVx1_ASAP7_75t_L g1695 ( .A(n_15), .Y(n_1695) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_16), .A2(n_285), .B1(n_440), .B2(n_445), .C(n_447), .Y(n_439) );
INVx1_ASAP7_75t_L g575 ( .A(n_16), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g1603 ( .A1(n_17), .A2(n_63), .B1(n_1069), .B2(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1621 ( .A(n_17), .Y(n_1621) );
AOI22xp5_ASAP7_75t_L g1738 ( .A1(n_18), .A2(n_311), .B1(n_1739), .B2(n_1743), .Y(n_1738) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_19), .A2(n_255), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_19), .Y(n_1166) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_20), .Y(n_1073) );
CKINVDCx16_ASAP7_75t_R g1776 ( .A(n_21), .Y(n_1776) );
INVxp33_ASAP7_75t_L g1409 ( .A(n_22), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_22), .A2(n_215), .B1(n_1390), .B2(n_1476), .Y(n_1482) );
INVx1_ASAP7_75t_L g1988 ( .A(n_23), .Y(n_1988) );
AOI22xp33_ASAP7_75t_L g2016 ( .A1(n_23), .A2(n_125), .B1(n_659), .B2(n_2017), .Y(n_2016) );
INVxp33_ASAP7_75t_L g1642 ( .A(n_24), .Y(n_1642) );
AOI221xp5_ASAP7_75t_L g1662 ( .A1(n_24), .A2(n_81), .B1(n_553), .B2(n_838), .C(n_1663), .Y(n_1662) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_25), .A2(n_69), .B1(n_939), .B2(n_1017), .C(n_1020), .Y(n_1016) );
INVx1_ASAP7_75t_L g1052 ( .A(n_25), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1589 ( .A1(n_26), .A2(n_364), .B1(n_974), .B2(n_1561), .C(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1613 ( .A(n_26), .Y(n_1613) );
CKINVDCx5p33_ASAP7_75t_R g2040 ( .A(n_27), .Y(n_2040) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_28), .A2(n_360), .B1(n_733), .B2(n_734), .Y(n_1499) );
INVxp67_ASAP7_75t_SL g1532 ( .A(n_28), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_29), .A2(n_375), .B1(n_423), .B2(n_433), .Y(n_422) );
INVx1_ASAP7_75t_L g518 ( .A(n_29), .Y(n_518) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_30), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_30), .A2(n_354), .B1(n_649), .B2(n_652), .C(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1651 ( .A1(n_31), .A2(n_357), .B1(n_800), .B2(n_1652), .Y(n_1651) );
INVxp67_ASAP7_75t_SL g1668 ( .A(n_31), .Y(n_1668) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_32), .A2(n_243), .B1(n_653), .B2(n_664), .C(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1279 ( .A(n_32), .Y(n_1279) );
INVx1_ASAP7_75t_L g1037 ( .A(n_33), .Y(n_1037) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_34), .A2(n_324), .B1(n_591), .B2(n_693), .C(n_889), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_34), .A2(n_324), .B1(n_931), .B2(n_932), .Y(n_930) );
INVxp33_ASAP7_75t_SL g765 ( .A(n_35), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_35), .A2(n_144), .B1(n_553), .B2(n_836), .C(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g383 ( .A(n_36), .Y(n_383) );
INVx1_ASAP7_75t_L g468 ( .A(n_37), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_37), .A2(n_335), .B1(n_550), .B2(n_553), .Y(n_549) );
INVxp33_ASAP7_75t_SL g687 ( .A(n_38), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_38), .A2(n_295), .B1(n_445), .B2(n_729), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g2064 ( .A(n_39), .Y(n_2064) );
AOI22xp5_ASAP7_75t_L g1762 ( .A1(n_40), .A2(n_172), .B1(n_1727), .B2(n_1735), .Y(n_1762) );
INVx1_ASAP7_75t_L g1346 ( .A(n_41), .Y(n_1346) );
OAI221xp5_ASAP7_75t_L g1124 ( .A1(n_42), .A2(n_70), .B1(n_691), .B2(n_693), .C(n_889), .Y(n_1124) );
OAI222xp33_ASAP7_75t_L g1150 ( .A1(n_42), .A2(n_70), .B1(n_239), .B2(n_931), .C1(n_932), .C2(n_1036), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_43), .A2(n_235), .B1(n_1764), .B2(n_1795), .Y(n_1794) );
AOI21xp33_ASAP7_75t_L g1084 ( .A1(n_44), .A2(n_1085), .B(n_1086), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_44), .A2(n_91), .B1(n_577), .B2(n_623), .C(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1502 ( .A(n_45), .Y(n_1502) );
OAI221xp5_ASAP7_75t_L g1514 ( .A1(n_45), .A2(n_317), .B1(n_682), .B2(n_684), .C(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1646 ( .A(n_46), .Y(n_1646) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_47), .A2(n_356), .B1(n_574), .B2(n_1558), .Y(n_1557) );
OAI22xp5_ASAP7_75t_L g1578 ( .A1(n_47), .A2(n_264), .B1(n_1069), .B2(n_1579), .Y(n_1578) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_48), .Y(n_911) );
INVx1_ASAP7_75t_L g494 ( .A(n_49), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_49), .A2(n_343), .B1(n_536), .B2(n_546), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g1998 ( .A(n_50), .Y(n_1998) );
AOI22xp5_ASAP7_75t_L g1746 ( .A1(n_51), .A2(n_140), .B1(n_1727), .B2(n_1735), .Y(n_1746) );
AO221x2_ASAP7_75t_L g1752 ( .A1(n_52), .A2(n_265), .B1(n_1739), .B2(n_1743), .C(n_1753), .Y(n_1752) );
CKINVDCx16_ASAP7_75t_R g1492 ( .A(n_53), .Y(n_1492) );
CKINVDCx5p33_ASAP7_75t_R g1601 ( .A(n_54), .Y(n_1601) );
AOI22xp5_ASAP7_75t_SL g1781 ( .A1(n_55), .A2(n_254), .B1(n_1743), .B2(n_1764), .Y(n_1781) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_56), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_56), .A2(n_224), .B1(n_656), .B2(n_659), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g1134 ( .A(n_57), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1655 ( .A1(n_58), .A2(n_210), .B1(n_1357), .B2(n_1656), .Y(n_1655) );
OAI22xp5_ASAP7_75t_L g1672 ( .A1(n_58), .A2(n_210), .B1(n_869), .B2(n_871), .Y(n_1672) );
INVx1_ASAP7_75t_L g711 ( .A(n_59), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g1355 ( .A1(n_60), .A2(n_102), .B1(n_440), .B2(n_652), .C(n_653), .Y(n_1355) );
INVxp67_ASAP7_75t_L g1388 ( .A(n_60), .Y(n_1388) );
INVxp67_ASAP7_75t_L g1186 ( .A(n_61), .Y(n_1186) );
INVx1_ASAP7_75t_L g1549 ( .A(n_62), .Y(n_1549) );
INVx1_ASAP7_75t_L g1623 ( .A(n_63), .Y(n_1623) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_64), .A2(n_168), .B1(n_1046), .B2(n_1552), .Y(n_1551) );
AOI221xp5_ASAP7_75t_L g1560 ( .A1(n_64), .A2(n_228), .B1(n_927), .B2(n_1561), .C(n_1563), .Y(n_1560) );
CKINVDCx14_ASAP7_75t_R g1833 ( .A(n_65), .Y(n_1833) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_66), .A2(n_216), .B1(n_742), .B2(n_744), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g1523 ( .A1(n_66), .A2(n_216), .B1(n_550), .B2(n_1524), .Y(n_1523) );
OAI221xp5_ASAP7_75t_L g1075 ( .A1(n_67), .A2(n_157), .B1(n_1071), .B2(n_1076), .C(n_1077), .Y(n_1075) );
INVx1_ASAP7_75t_L g1114 ( .A(n_67), .Y(n_1114) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_68), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_68), .A2(n_112), .B1(n_663), .B2(n_927), .Y(n_1236) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_69), .A2(n_217), .B1(n_1048), .B2(n_1050), .C(n_1051), .Y(n_1047) );
INVx1_ASAP7_75t_L g770 ( .A(n_71), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g1132 ( .A(n_72), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_73), .A2(n_96), .B1(n_803), .B2(n_805), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_73), .A2(n_96), .B1(n_869), .B2(n_871), .Y(n_868) );
AOI21xp33_ASAP7_75t_L g961 ( .A1(n_74), .A2(n_455), .B(n_727), .Y(n_961) );
INVxp33_ASAP7_75t_L g984 ( .A(n_74), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_75), .A2(n_209), .B1(n_724), .B2(n_1318), .Y(n_1317) );
INVxp67_ASAP7_75t_SL g1331 ( .A(n_75), .Y(n_1331) );
XOR2x2_ASAP7_75t_L g1634 ( .A(n_76), .B(n_1635), .Y(n_1634) );
OAI22xp33_ASAP7_75t_L g1255 ( .A1(n_77), .A2(n_225), .B1(n_672), .B2(n_1230), .Y(n_1255) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_77), .A2(n_225), .B1(n_599), .B2(n_693), .C(n_1274), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1792 ( .A1(n_78), .A2(n_220), .B1(n_1727), .B2(n_1793), .Y(n_1792) );
INVx1_ASAP7_75t_L g782 ( .A(n_79), .Y(n_782) );
INVx1_ASAP7_75t_L g1361 ( .A(n_80), .Y(n_1361) );
INVxp33_ASAP7_75t_L g1643 ( .A(n_81), .Y(n_1643) );
INVx1_ASAP7_75t_L g1215 ( .A(n_82), .Y(n_1215) );
INVx1_ASAP7_75t_L g1321 ( .A(n_83), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_84), .Y(n_813) );
XNOR2x2_ASAP7_75t_L g1586 ( .A(n_85), .B(n_1587), .Y(n_1586) );
INVxp33_ASAP7_75t_L g1680 ( .A(n_86), .Y(n_1680) );
AOI22xp33_ASAP7_75t_L g1705 ( .A1(n_86), .A2(n_292), .B1(n_470), .B2(n_1318), .Y(n_1705) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_87), .A2(n_286), .B1(n_720), .B2(n_800), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_87), .A2(n_286), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
INVx1_ASAP7_75t_L g1544 ( .A(n_88), .Y(n_1544) );
CKINVDCx5p33_ASAP7_75t_R g2004 ( .A(n_89), .Y(n_2004) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_90), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_91), .A2(n_250), .B1(n_796), .B2(n_1018), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_92), .A2(n_189), .B1(n_445), .B2(n_801), .Y(n_1034) );
INVx1_ASAP7_75t_L g1060 ( .A(n_92), .Y(n_1060) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_93), .A2(n_295), .B1(n_682), .B2(n_684), .C(n_686), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_93), .A2(n_316), .B1(n_720), .B2(n_724), .C(n_727), .Y(n_719) );
INVxp33_ASAP7_75t_SL g1512 ( .A(n_94), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_94), .A2(n_358), .B1(n_1524), .B2(n_1526), .Y(n_1528) );
CKINVDCx14_ASAP7_75t_R g1754 ( .A(n_95), .Y(n_1754) );
INVx1_ASAP7_75t_L g674 ( .A(n_97), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_98), .Y(n_913) );
BUFx2_ASAP7_75t_L g410 ( .A(n_99), .Y(n_410) );
OR2x2_ASAP7_75t_L g501 ( .A(n_99), .B(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g505 ( .A(n_99), .Y(n_505) );
INVx1_ASAP7_75t_L g558 ( .A(n_99), .Y(n_558) );
INVx1_ASAP7_75t_L g1271 ( .A(n_100), .Y(n_1271) );
AOI221xp5_ASAP7_75t_L g2061 ( .A1(n_101), .A2(n_320), .B1(n_574), .B2(n_604), .C(n_1473), .Y(n_2061) );
INVx1_ASAP7_75t_L g2073 ( .A(n_101), .Y(n_2073) );
INVxp33_ASAP7_75t_SL g1386 ( .A(n_102), .Y(n_1386) );
INVxp33_ASAP7_75t_L g1683 ( .A(n_103), .Y(n_1683) );
INVxp67_ASAP7_75t_L g1421 ( .A(n_104), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g2002 ( .A(n_105), .Y(n_2002) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_106), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g1979 ( .A(n_107), .Y(n_1979) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_108), .A2(n_240), .B1(n_965), .B2(n_967), .C(n_970), .Y(n_964) );
INVxp67_ASAP7_75t_SL g998 ( .A(n_108), .Y(n_998) );
INVx1_ASAP7_75t_L g898 ( .A(n_109), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_109), .A2(n_296), .B1(n_925), .B2(n_926), .Y(n_924) );
AOI221xp5_ASAP7_75t_SL g1026 ( .A1(n_110), .A2(n_116), .B1(n_727), .B2(n_743), .C(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1045 ( .A(n_110), .Y(n_1045) );
INVxp33_ASAP7_75t_L g1455 ( .A(n_111), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_111), .A2(n_322), .B1(n_800), .B2(n_1227), .Y(n_1463) );
INVxp33_ASAP7_75t_L g1199 ( .A(n_112), .Y(n_1199) );
INVx1_ASAP7_75t_L g1022 ( .A(n_113), .Y(n_1022) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_114), .A2(n_139), .B1(n_791), .B2(n_1301), .C(n_1303), .Y(n_1300) );
INVxp33_ASAP7_75t_L g1325 ( .A(n_114), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_115), .A2(n_193), .B1(n_599), .B2(n_691), .C(n_692), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_115), .A2(n_193), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g1044 ( .A(n_116), .Y(n_1044) );
XOR2x2_ASAP7_75t_L g1064 ( .A(n_117), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1368 ( .A(n_118), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g2065 ( .A(n_119), .Y(n_2065) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_120), .A2(n_239), .B1(n_500), .B2(n_1122), .Y(n_1121) );
CKINVDCx5p33_ASAP7_75t_R g1164 ( .A(n_120), .Y(n_1164) );
OA22x2_ASAP7_75t_L g1291 ( .A1(n_121), .A2(n_1292), .B1(n_1293), .B2(n_1340), .Y(n_1291) );
CKINVDCx16_ASAP7_75t_R g1340 ( .A(n_121), .Y(n_1340) );
INVxp33_ASAP7_75t_L g1448 ( .A(n_122), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_122), .A2(n_302), .B1(n_1465), .B2(n_1466), .Y(n_1464) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_123), .Y(n_909) );
INVx1_ASAP7_75t_L g1221 ( .A(n_124), .Y(n_1221) );
INVx1_ASAP7_75t_L g1993 ( .A(n_125), .Y(n_1993) );
INVxp67_ASAP7_75t_L g1195 ( .A(n_126), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_126), .A2(n_162), .B1(n_445), .B2(n_738), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_127), .A2(n_279), .B1(n_660), .B2(n_792), .Y(n_1092) );
OAI211xp5_ASAP7_75t_L g1094 ( .A1(n_127), .A2(n_1095), .B(n_1097), .C(n_1099), .Y(n_1094) );
INVx1_ASAP7_75t_L g2038 ( .A(n_128), .Y(n_2038) );
AOI221xp5_ASAP7_75t_L g2050 ( .A1(n_128), .A2(n_152), .B1(n_577), .B2(n_2051), .C(n_2052), .Y(n_2050) );
INVx1_ASAP7_75t_L g1240 ( .A(n_129), .Y(n_1240) );
OAI22xp33_ASAP7_75t_SL g1605 ( .A1(n_130), .A2(n_167), .B1(n_448), .B2(n_935), .Y(n_1605) );
INVx1_ASAP7_75t_L g1624 ( .A(n_130), .Y(n_1624) );
CKINVDCx5p33_ASAP7_75t_R g1250 ( .A(n_131), .Y(n_1250) );
INVx1_ASAP7_75t_L g1694 ( .A(n_132), .Y(n_1694) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_133), .A2(n_344), .B1(n_795), .B2(n_797), .Y(n_794) );
INVxp67_ASAP7_75t_SL g863 ( .A(n_133), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_134), .A2(n_198), .B1(n_652), .B2(n_653), .C(n_667), .Y(n_1033) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_134), .A2(n_189), .B1(n_1055), .B2(n_1057), .C(n_1059), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g2031 ( .A(n_135), .B(n_2032), .Y(n_2031) );
CKINVDCx5p33_ASAP7_75t_R g1598 ( .A(n_136), .Y(n_1598) );
INVx1_ASAP7_75t_L g1576 ( .A(n_137), .Y(n_1576) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_138), .Y(n_916) );
INVxp33_ASAP7_75t_L g1327 ( .A(n_139), .Y(n_1327) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_141), .A2(n_326), .B1(n_470), .B2(n_473), .C(n_477), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_141), .A2(n_232), .B1(n_536), .B2(n_541), .Y(n_535) );
OAI22xp33_ASAP7_75t_L g1070 ( .A1(n_142), .A2(n_329), .B1(n_484), .B2(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_142), .A2(n_196), .B1(n_529), .B2(n_554), .Y(n_1108) );
INVxp67_ASAP7_75t_L g1194 ( .A(n_143), .Y(n_1194) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_143), .A2(n_203), .B1(n_455), .B2(n_727), .C(n_1227), .Y(n_1226) );
INVxp33_ASAP7_75t_SL g760 ( .A(n_144), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_145), .A2(n_196), .B1(n_935), .B2(n_1069), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_145), .A2(n_329), .B1(n_542), .B2(n_1107), .Y(n_1106) );
AOI21xp5_ASAP7_75t_L g1093 ( .A1(n_146), .A2(n_663), .B(n_665), .Y(n_1093) );
INVx1_ASAP7_75t_L g1100 ( .A(n_146), .Y(n_1100) );
XNOR2xp5_ASAP7_75t_L g750 ( .A(n_147), .B(n_751), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g1247 ( .A(n_148), .Y(n_1247) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_149), .A2(n_187), .B1(n_591), .B2(n_596), .C(n_599), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_149), .A2(n_187), .B1(n_670), .B2(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g896 ( .A(n_150), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g1508 ( .A1(n_151), .A2(n_323), .B1(n_667), .B2(n_739), .C(n_740), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g1525 ( .A1(n_151), .A2(n_323), .B1(n_1526), .B2(n_1527), .Y(n_1525) );
INVx1_ASAP7_75t_L g2045 ( .A(n_152), .Y(n_2045) );
INVx1_ASAP7_75t_L g1546 ( .A(n_153), .Y(n_1546) );
XNOR2xp5_ASAP7_75t_L g1675 ( .A(n_154), .B(n_1676), .Y(n_1675) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_155), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1196 ( .A1(n_156), .A2(n_191), .B1(n_691), .B2(n_693), .C(n_889), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_156), .A2(n_191), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
INVx1_ASAP7_75t_L g1098 ( .A(n_157), .Y(n_1098) );
INVx1_ASAP7_75t_L g1024 ( .A(n_158), .Y(n_1024) );
AOI22xp5_ASAP7_75t_SL g1780 ( .A1(n_159), .A2(n_178), .B1(n_1727), .B2(n_1735), .Y(n_1780) );
CKINVDCx5p33_ASAP7_75t_R g1140 ( .A(n_160), .Y(n_1140) );
INVx1_ASAP7_75t_L g1423 ( .A(n_161), .Y(n_1423) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_161), .A2(n_310), .B1(n_1442), .B2(n_1444), .Y(n_1441) );
INVxp67_ASAP7_75t_L g1191 ( .A(n_162), .Y(n_1191) );
INVxp33_ASAP7_75t_SL g1511 ( .A(n_163), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_163), .A2(n_306), .B1(n_550), .B2(n_1527), .Y(n_1529) );
INVx1_ASAP7_75t_L g1731 ( .A(n_164), .Y(n_1731) );
INVx1_ASAP7_75t_L g1313 ( .A(n_165), .Y(n_1313) );
AOI221xp5_ASAP7_75t_L g1314 ( .A1(n_166), .A2(n_231), .B1(n_1085), .B2(n_1315), .C(n_1316), .Y(n_1314) );
INVxp67_ASAP7_75t_SL g1336 ( .A(n_166), .Y(n_1336) );
INVx1_ASAP7_75t_L g1619 ( .A(n_167), .Y(n_1619) );
INVx1_ASAP7_75t_L g1564 ( .A(n_168), .Y(n_1564) );
CKINVDCx16_ASAP7_75t_R g1773 ( .A(n_169), .Y(n_1773) );
INVx1_ASAP7_75t_L g1647 ( .A(n_170), .Y(n_1647) );
INVxp67_ASAP7_75t_L g1692 ( .A(n_171), .Y(n_1692) );
AOI22xp33_ASAP7_75t_L g1710 ( .A1(n_171), .A2(n_211), .B1(n_656), .B2(n_744), .Y(n_1710) );
INVx1_ASAP7_75t_L g1989 ( .A(n_173), .Y(n_1989) );
AOI221xp5_ASAP7_75t_L g2013 ( .A1(n_173), .A2(n_222), .B1(n_496), .B2(n_740), .C(n_2014), .Y(n_2013) );
INVx1_ASAP7_75t_L g1732 ( .A(n_174), .Y(n_1732) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_174), .B(n_1730), .Y(n_1737) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_175), .A2(n_260), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_175), .A2(n_260), .B1(n_897), .B2(n_1042), .C(n_1043), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g1650 ( .A1(n_176), .A2(n_204), .B1(n_791), .B2(n_797), .Y(n_1650) );
INVxp67_ASAP7_75t_SL g1667 ( .A(n_176), .Y(n_1667) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_177), .A2(n_232), .B1(n_480), .B2(n_483), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_177), .A2(n_326), .B1(n_529), .B2(n_532), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_179), .A2(n_455), .B(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g572 ( .A(n_179), .Y(n_572) );
INVx1_ASAP7_75t_L g1981 ( .A(n_180), .Y(n_1981) );
AOI21xp33_ASAP7_75t_L g2011 ( .A1(n_180), .A2(n_658), .B(n_727), .Y(n_2011) );
INVx1_ASAP7_75t_L g1698 ( .A(n_181), .Y(n_1698) );
INVx2_ASAP7_75t_L g395 ( .A(n_182), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g2037 ( .A(n_183), .Y(n_2037) );
INVx1_ASAP7_75t_L g1982 ( .A(n_184), .Y(n_1982) );
AOI22xp33_ASAP7_75t_L g2010 ( .A1(n_184), .A2(n_237), .B1(n_442), .B2(n_660), .Y(n_2010) );
OAI22x1_ASAP7_75t_SL g1397 ( .A1(n_185), .A2(n_1398), .B1(n_1484), .B2(n_1485), .Y(n_1397) );
INVx1_ASAP7_75t_L g1484 ( .A(n_185), .Y(n_1484) );
INVx1_ASAP7_75t_L g421 ( .A(n_186), .Y(n_421) );
BUFx3_ASAP7_75t_L g438 ( .A(n_186), .Y(n_438) );
INVx1_ASAP7_75t_L g1640 ( .A(n_188), .Y(n_1640) );
INVxp33_ASAP7_75t_L g588 ( .A(n_190), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_190), .A2(n_238), .B1(n_663), .B2(n_664), .C(n_665), .Y(n_662) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_192), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g1597 ( .A(n_194), .Y(n_1597) );
AOI22xp33_ASAP7_75t_L g2060 ( .A1(n_195), .A2(n_337), .B1(n_1107), .B2(n_1390), .Y(n_2060) );
AOI22xp33_ASAP7_75t_L g2075 ( .A1(n_195), .A2(n_337), .B1(n_791), .B2(n_805), .Y(n_2075) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_197), .Y(n_1372) );
INVx1_ASAP7_75t_L g1061 ( .A(n_198), .Y(n_1061) );
OAI22xp33_ASAP7_75t_R g1309 ( .A1(n_199), .A2(n_369), .B1(n_734), .B2(n_931), .Y(n_1309) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_199), .A2(n_369), .B1(n_599), .B2(n_691), .C(n_692), .Y(n_1328) );
OAI221xp5_ASAP7_75t_SL g955 ( .A1(n_200), .A2(n_361), .B1(n_670), .B2(n_734), .C(n_956), .Y(n_955) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_200), .A2(n_361), .B1(n_596), .B2(n_691), .C(n_988), .Y(n_987) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_201), .Y(n_884) );
INVx1_ASAP7_75t_L g1320 ( .A(n_202), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1192 ( .A(n_203), .Y(n_1192) );
INVxp67_ASAP7_75t_SL g1670 ( .A(n_204), .Y(n_1670) );
INVx1_ASAP7_75t_L g1023 ( .A(n_205), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1138 ( .A(n_206), .Y(n_1138) );
CKINVDCx5p33_ASAP7_75t_R g1658 ( .A(n_207), .Y(n_1658) );
INVxp33_ASAP7_75t_SL g1539 ( .A(n_208), .Y(n_1539) );
AOI221xp5_ASAP7_75t_L g1565 ( .A1(n_208), .A2(n_267), .B1(n_927), .B2(n_1566), .C(n_1568), .Y(n_1565) );
INVxp67_ASAP7_75t_SL g1337 ( .A(n_209), .Y(n_1337) );
INVxp33_ASAP7_75t_L g1688 ( .A(n_211), .Y(n_1688) );
INVx1_ASAP7_75t_L g977 ( .A(n_212), .Y(n_977) );
AOI221xp5_ASAP7_75t_L g1369 ( .A1(n_213), .A2(n_328), .B1(n_458), .B2(n_480), .C(n_652), .Y(n_1369) );
INVxp33_ASAP7_75t_SL g1379 ( .A(n_213), .Y(n_1379) );
INVx1_ASAP7_75t_L g417 ( .A(n_214), .Y(n_417) );
INVx1_ASAP7_75t_L g460 ( .A(n_214), .Y(n_460) );
INVxp33_ASAP7_75t_L g1418 ( .A(n_215), .Y(n_1418) );
INVx1_ASAP7_75t_L g1021 ( .A(n_217), .Y(n_1021) );
INVxp33_ASAP7_75t_SL g585 ( .A(n_218), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_218), .A2(n_226), .B1(n_667), .B2(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g2041 ( .A(n_219), .Y(n_2041) );
OAI221xp5_ASAP7_75t_L g2056 ( .A1(n_219), .A2(n_248), .B1(n_844), .B2(n_2057), .C(n_2059), .Y(n_2056) );
CKINVDCx20_ASAP7_75t_R g1831 ( .A(n_221), .Y(n_1831) );
INVx1_ASAP7_75t_L g1991 ( .A(n_222), .Y(n_1991) );
INVx1_ASAP7_75t_L g1363 ( .A(n_223), .Y(n_1363) );
OAI221xp5_ASAP7_75t_L g1380 ( .A1(n_223), .A2(n_262), .B1(n_591), .B2(n_988), .C(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g624 ( .A(n_224), .Y(n_624) );
INVxp33_ASAP7_75t_SL g589 ( .A(n_226), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_227), .Y(n_1089) );
INVx1_ASAP7_75t_L g1550 ( .A(n_228), .Y(n_1550) );
AOI221xp5_ASAP7_75t_L g1595 ( .A1(n_229), .A2(n_331), .B1(n_805), .B2(n_1085), .C(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1627 ( .A(n_229), .Y(n_1627) );
AOI22xp33_ASAP7_75t_SL g1654 ( .A1(n_230), .A2(n_301), .B1(n_724), .B2(n_797), .Y(n_1654) );
OAI211xp5_ASAP7_75t_SL g1660 ( .A1(n_230), .A2(n_824), .B(n_1661), .C(n_1664), .Y(n_1660) );
INVxp67_ASAP7_75t_SL g1332 ( .A(n_231), .Y(n_1332) );
INVx1_ASAP7_75t_L g578 ( .A(n_233), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g1997 ( .A(n_234), .Y(n_1997) );
XNOR2x1_ASAP7_75t_L g877 ( .A(n_235), .B(n_878), .Y(n_877) );
CKINVDCx14_ASAP7_75t_R g1756 ( .A(n_236), .Y(n_1756) );
INVx1_ASAP7_75t_L g1977 ( .A(n_237), .Y(n_1977) );
INVxp33_ASAP7_75t_L g586 ( .A(n_238), .Y(n_586) );
INVx1_ASAP7_75t_L g996 ( .A(n_240), .Y(n_996) );
INVx1_ASAP7_75t_L g882 ( .A(n_241), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_242), .A2(n_252), .B1(n_470), .B2(n_805), .Y(n_1254) );
INVx1_ASAP7_75t_L g1267 ( .A(n_242), .Y(n_1267) );
INVx1_ASAP7_75t_L g1281 ( .A(n_243), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_244), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_244), .A2(n_261), .B1(n_442), .B2(n_1234), .C(n_1235), .Y(n_1233) );
INVx1_ASAP7_75t_L g1307 ( .A(n_245), .Y(n_1307) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_246), .A2(n_330), .B1(n_797), .B2(n_800), .Y(n_799) );
OAI221xp5_ASAP7_75t_L g845 ( .A1(n_246), .A2(n_846), .B1(n_848), .B2(n_858), .C(n_866), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_247), .A2(n_319), .B1(n_973), .B2(n_974), .Y(n_972) );
INVx1_ASAP7_75t_L g993 ( .A(n_247), .Y(n_993) );
INVx1_ASAP7_75t_L g2042 ( .A(n_248), .Y(n_2042) );
INVx1_ASAP7_75t_L g1298 ( .A(n_249), .Y(n_1298) );
INVx1_ASAP7_75t_L g1111 ( .A(n_250), .Y(n_1111) );
INVxp67_ASAP7_75t_L g1691 ( .A(n_251), .Y(n_1691) );
AOI221xp5_ASAP7_75t_L g1708 ( .A1(n_251), .A2(n_368), .B1(n_652), .B2(n_653), .C(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1272 ( .A(n_252), .Y(n_1272) );
INVx1_ASAP7_75t_L g678 ( .A(n_253), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g1241 ( .A(n_254), .B(n_1242), .Y(n_1241) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_255), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_256), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_257), .A2(n_313), .B1(n_973), .B2(n_1357), .Y(n_1356) );
INVxp67_ASAP7_75t_L g1384 ( .A(n_257), .Y(n_1384) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_258), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_258), .A2(n_300), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g712 ( .A(n_259), .Y(n_712) );
INVxp33_ASAP7_75t_L g1203 ( .A(n_261), .Y(n_1203) );
INVx1_ASAP7_75t_L g1364 ( .A(n_262), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_263), .A2(n_273), .B1(n_442), .B2(n_660), .Y(n_960) );
INVxp33_ASAP7_75t_L g985 ( .A(n_263), .Y(n_985) );
INVxp67_ASAP7_75t_SL g1556 ( .A(n_264), .Y(n_1556) );
INVx1_ASAP7_75t_L g1360 ( .A(n_266), .Y(n_1360) );
INVxp33_ASAP7_75t_SL g1542 ( .A(n_267), .Y(n_1542) );
CKINVDCx20_ASAP7_75t_R g1770 ( .A(n_268), .Y(n_1770) );
BUFx3_ASAP7_75t_L g420 ( .A(n_269), .Y(n_420) );
INVx1_ASAP7_75t_L g444 ( .A(n_269), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_270), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1593 ( .A(n_271), .Y(n_1593) );
AO221x2_ASAP7_75t_L g1828 ( .A1(n_272), .A2(n_346), .B1(n_1795), .B2(n_1829), .C(n_1830), .Y(n_1828) );
INVxp33_ASAP7_75t_L g981 ( .A(n_273), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g1747 ( .A1(n_274), .A2(n_275), .B1(n_1739), .B2(n_1743), .Y(n_1747) );
INVx1_ASAP7_75t_L g1007 ( .A(n_275), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_276), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_276), .B(n_352), .Y(n_502) );
INVx1_ASAP7_75t_L g562 ( .A(n_276), .Y(n_562) );
AND2x2_ASAP7_75t_L g568 ( .A(n_276), .B(n_561), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_277), .Y(n_905) );
INVx1_ASAP7_75t_L g709 ( .A(n_278), .Y(n_709) );
INVx1_ASAP7_75t_L g1102 ( .A(n_279), .Y(n_1102) );
AOI21xp5_ASAP7_75t_L g1503 ( .A1(n_280), .A2(n_1504), .B(n_1505), .Y(n_1503) );
INVx1_ASAP7_75t_L g1518 ( .A(n_280), .Y(n_1518) );
OAI332xp33_ASAP7_75t_L g1125 ( .A1(n_281), .A2(n_556), .A3(n_603), .B1(n_1126), .B2(n_1129), .B3(n_1133), .C1(n_1139), .C2(n_1142), .Y(n_1125) );
INVx1_ASAP7_75t_L g1168 ( .A(n_281), .Y(n_1168) );
INVx1_ASAP7_75t_L g706 ( .A(n_282), .Y(n_706) );
INVx1_ASAP7_75t_L g1575 ( .A(n_283), .Y(n_1575) );
OR2x2_ASAP7_75t_L g416 ( .A(n_284), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g428 ( .A(n_284), .Y(n_428) );
INVx1_ASAP7_75t_L g564 ( .A(n_285), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_287), .Y(n_1128) );
INVx1_ASAP7_75t_L g1213 ( .A(n_288), .Y(n_1213) );
INVx1_ASAP7_75t_L g1371 ( .A(n_289), .Y(n_1371) );
CKINVDCx16_ASAP7_75t_R g1012 ( .A(n_290), .Y(n_1012) );
INVx1_ASAP7_75t_L g629 ( .A(n_291), .Y(n_629) );
INVxp33_ASAP7_75t_SL g1684 ( .A(n_292), .Y(n_1684) );
INVx1_ASAP7_75t_L g497 ( .A(n_293), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_294), .A2(n_305), .B1(n_791), .B2(n_793), .Y(n_790) );
INVxp67_ASAP7_75t_L g852 ( .A(n_294), .Y(n_852) );
INVx1_ASAP7_75t_L g892 ( .A(n_296), .Y(n_892) );
INVx1_ASAP7_75t_L g1354 ( .A(n_297), .Y(n_1354) );
INVx1_ASAP7_75t_L g2068 ( .A(n_298), .Y(n_2068) );
AOI22xp33_ASAP7_75t_L g2078 ( .A1(n_298), .A2(n_327), .B1(n_791), .B2(n_1301), .Y(n_2078) );
INVx1_ASAP7_75t_L g963 ( .A(n_299), .Y(n_963) );
INVxp33_ASAP7_75t_SL g700 ( .A(n_300), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g1665 ( .A1(n_301), .A2(n_846), .B1(n_866), .B2(n_1666), .C(n_1669), .Y(n_1665) );
INVxp67_ASAP7_75t_L g1452 ( .A(n_302), .Y(n_1452) );
INVx1_ASAP7_75t_L g1414 ( .A(n_303), .Y(n_1414) );
AOI22xp5_ASAP7_75t_SL g1763 ( .A1(n_304), .A2(n_308), .B1(n_1743), .B2(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1972 ( .A(n_304), .Y(n_1972) );
AOI22xp33_ASAP7_75t_L g2026 ( .A1(n_304), .A2(n_2027), .B1(n_2030), .B2(n_2079), .Y(n_2026) );
INVxp67_ASAP7_75t_L g849 ( .A(n_305), .Y(n_849) );
INVxp67_ASAP7_75t_SL g1507 ( .A(n_306), .Y(n_1507) );
AOI221xp5_ASAP7_75t_L g1500 ( .A1(n_307), .A2(n_317), .B1(n_667), .B2(n_744), .C(n_1501), .Y(n_1500) );
INVxp33_ASAP7_75t_L g1516 ( .A(n_307), .Y(n_1516) );
INVx1_ASAP7_75t_L g1366 ( .A(n_309), .Y(n_1366) );
INVx1_ASAP7_75t_L g1428 ( .A(n_310), .Y(n_1428) );
CKINVDCx5p33_ASAP7_75t_R g1295 ( .A(n_312), .Y(n_1295) );
INVxp67_ASAP7_75t_L g1391 ( .A(n_313), .Y(n_1391) );
INVx1_ASAP7_75t_L g776 ( .A(n_314), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_315), .A2(n_333), .B1(n_729), .B2(n_1318), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1475 ( .A1(n_315), .A2(n_333), .B1(n_1476), .B2(n_1478), .Y(n_1475) );
INVxp33_ASAP7_75t_SL g688 ( .A(n_316), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g1592 ( .A(n_318), .Y(n_1592) );
INVx1_ASAP7_75t_L g1000 ( .A(n_319), .Y(n_1000) );
INVx1_ASAP7_75t_L g2074 ( .A(n_320), .Y(n_2074) );
CKINVDCx5p33_ASAP7_75t_R g2001 ( .A(n_321), .Y(n_2001) );
INVxp67_ASAP7_75t_L g1435 ( .A(n_322), .Y(n_1435) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_325), .A2(n_363), .B1(n_668), .B2(n_1146), .Y(n_1259) );
INVx1_ASAP7_75t_L g1284 ( .A(n_325), .Y(n_1284) );
INVx1_ASAP7_75t_L g2067 ( .A(n_327), .Y(n_2067) );
INVxp33_ASAP7_75t_SL g1377 ( .A(n_328), .Y(n_1377) );
OAI211xp5_ASAP7_75t_SL g823 ( .A1(n_330), .A2(n_824), .B(n_829), .C(n_840), .Y(n_823) );
INVx1_ASAP7_75t_L g1629 ( .A(n_331), .Y(n_1629) );
INVx1_ASAP7_75t_L g1220 ( .A(n_332), .Y(n_1220) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_334), .Y(n_703) );
INVx1_ASAP7_75t_L g490 ( .A(n_335), .Y(n_490) );
INVx1_ASAP7_75t_L g957 ( .A(n_336), .Y(n_957) );
INVx1_ASAP7_75t_L g580 ( .A(n_338), .Y(n_580) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_339), .B(n_383), .Y(n_1734) );
AND3x2_ASAP7_75t_L g1740 ( .A(n_339), .B(n_383), .C(n_1731), .Y(n_1740) );
INVx2_ASAP7_75t_L g396 ( .A(n_341), .Y(n_396) );
XNOR2x2_ASAP7_75t_L g1535 ( .A(n_342), .B(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g413 ( .A(n_343), .Y(n_413) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_344), .Y(n_860) );
INVx1_ASAP7_75t_L g1540 ( .A(n_345), .Y(n_1540) );
CKINVDCx5p33_ASAP7_75t_R g1127 ( .A(n_347), .Y(n_1127) );
INVx1_ASAP7_75t_L g1305 ( .A(n_348), .Y(n_1305) );
INVx1_ASAP7_75t_L g632 ( .A(n_349), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g1609 ( .A(n_350), .Y(n_1609) );
OAI221xp5_ASAP7_75t_L g1983 ( .A1(n_351), .A2(n_355), .B1(n_591), .B2(n_599), .C(n_1381), .Y(n_1983) );
OAI221xp5_ASAP7_75t_L g2007 ( .A1(n_351), .A2(n_355), .B1(n_433), .B2(n_2008), .C(n_2009), .Y(n_2007) );
INVx1_ASAP7_75t_L g398 ( .A(n_352), .Y(n_398) );
INVx2_ASAP7_75t_L g561 ( .A(n_352), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1608 ( .A(n_353), .Y(n_1608) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_354), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g1580 ( .A1(n_356), .A2(n_370), .B1(n_441), .B2(n_1071), .Y(n_1580) );
INVxp67_ASAP7_75t_SL g1671 ( .A(n_357), .Y(n_1671) );
INVxp67_ASAP7_75t_SL g1498 ( .A(n_358), .Y(n_1498) );
INVx1_ASAP7_75t_L g630 ( .A(n_359), .Y(n_630) );
INVxp67_ASAP7_75t_SL g1531 ( .A(n_360), .Y(n_1531) );
INVx1_ASAP7_75t_L g1278 ( .A(n_363), .Y(n_1278) );
INVx1_ASAP7_75t_L g1617 ( .A(n_364), .Y(n_1617) );
INVx1_ASAP7_75t_L g1712 ( .A(n_365), .Y(n_1712) );
CKINVDCx5p33_ASAP7_75t_R g1495 ( .A(n_366), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g1248 ( .A(n_367), .Y(n_1248) );
INVxp33_ASAP7_75t_L g1689 ( .A(n_368), .Y(n_1689) );
INVxp67_ASAP7_75t_SL g1555 ( .A(n_370), .Y(n_1555) );
INVx1_ASAP7_75t_L g2044 ( .A(n_371), .Y(n_2044) );
AOI21xp5_ASAP7_75t_L g2054 ( .A1(n_371), .A2(n_838), .B(n_2055), .Y(n_2054) );
INVx1_ASAP7_75t_L g976 ( .A(n_372), .Y(n_976) );
INVx1_ASAP7_75t_L g637 ( .A(n_373), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_374), .Y(n_453) );
INVx1_ASAP7_75t_L g513 ( .A(n_375), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_399), .B(n_1718), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_386), .Y(n_380) );
AND2x4_ASAP7_75t_L g2025 ( .A(n_381), .B(n_387), .Y(n_2025) );
NOR2xp33_ASAP7_75t_SL g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_SL g2029 ( .A(n_382), .Y(n_2029) );
NAND2xp5_ASAP7_75t_L g2084 ( .A(n_382), .B(n_384), .Y(n_2084) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g2028 ( .A(n_384), .B(n_2029), .Y(n_2028) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_392), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g1458 ( .A(n_389), .B(n_505), .Y(n_1458) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g527 ( .A(n_390), .B(n_398), .Y(n_527) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g604 ( .A(n_391), .B(n_605), .Y(n_604) );
INVx8_ASAP7_75t_L g1454 ( .A(n_392), .Y(n_1454) );
OR2x6_ASAP7_75t_L g392 ( .A(n_393), .B(n_397), .Y(n_392) );
OR2x2_ASAP7_75t_L g500 ( .A(n_393), .B(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_393), .Y(n_609) );
INVx2_ASAP7_75t_SL g697 ( .A(n_393), .Y(n_697) );
INVx2_ASAP7_75t_SL g862 ( .A(n_393), .Y(n_862) );
INVx1_ASAP7_75t_L g992 ( .A(n_393), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_393), .A2(n_635), .B1(n_1081), .B2(n_1111), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1202 ( .A(n_393), .Y(n_1202) );
OR2x6_ASAP7_75t_L g1457 ( .A(n_393), .B(n_1447), .Y(n_1457) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g517 ( .A(n_395), .Y(n_517) );
INVx1_ASAP7_75t_L g522 ( .A(n_395), .Y(n_522) );
AND2x2_ASAP7_75t_L g531 ( .A(n_395), .B(n_396), .Y(n_531) );
INVx2_ASAP7_75t_L g538 ( .A(n_395), .Y(n_538) );
AND2x4_ASAP7_75t_L g544 ( .A(n_395), .B(n_523), .Y(n_544) );
INVx1_ASAP7_75t_L g511 ( .A(n_396), .Y(n_511) );
INVx2_ASAP7_75t_L g523 ( .A(n_396), .Y(n_523) );
INVx1_ASAP7_75t_L g540 ( .A(n_396), .Y(n_540) );
INVx1_ASAP7_75t_L g614 ( .A(n_396), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_396), .B(n_538), .Y(n_620) );
AND2x4_ASAP7_75t_L g1443 ( .A(n_397), .B(n_511), .Y(n_1443) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_398), .B(n_516), .Y(n_1444) );
OAI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_1487), .B(n_1715), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_1181), .Y(n_400) );
INVx2_ASAP7_75t_L g1488 ( .A(n_401), .Y(n_1488) );
AOI33xp33_ASAP7_75t_L g1715 ( .A1(n_401), .A2(n_1181), .A3(n_1182), .B1(n_1716), .B2(n_1717), .B3(n_2086), .Y(n_1715) );
INVx1_ASAP7_75t_L g1716 ( .A(n_401), .Y(n_1716) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_875), .B1(n_1178), .B2(n_1179), .Y(n_402) );
INVx1_ASAP7_75t_L g1178 ( .A(n_403), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_676), .B1(n_873), .B2(n_874), .Y(n_403) );
INVx1_ASAP7_75t_L g873 ( .A(n_404), .Y(n_873) );
XOR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_579), .Y(n_404) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_578), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_507), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B1(n_497), .B2(n_498), .Y(n_407) );
INVx2_ASAP7_75t_L g944 ( .A(n_408), .Y(n_944) );
OAI31xp33_ASAP7_75t_SL g1588 ( .A1(n_408), .A2(n_1589), .A3(n_1595), .B(n_1599), .Y(n_1588) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g643 ( .A(n_409), .Y(n_643) );
AND2x4_ASAP7_75t_L g1399 ( .A(n_409), .B(n_1400), .Y(n_1399) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g526 ( .A(n_410), .Y(n_526) );
OR2x6_ASAP7_75t_L g603 ( .A(n_410), .B(n_604), .Y(n_603) );
NAND3xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_461), .C(n_489), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B(n_422), .C(n_439), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_414), .A2(n_630), .B1(n_662), .B2(n_666), .C(n_669), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_414), .A2(n_491), .B1(n_709), .B2(n_711), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g943 ( .A1(n_414), .A2(n_491), .B1(n_909), .B2(n_911), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_414), .A2(n_491), .B1(n_976), .B2(n_977), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g1238 ( .A1(n_414), .A2(n_491), .B1(n_1215), .B2(n_1220), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_414), .A2(n_1250), .B1(n_1251), .B2(n_1254), .C(n_1255), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_414), .A2(n_491), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_414), .A2(n_491), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_414), .A2(n_491), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
AOI221xp5_ASAP7_75t_L g1701 ( .A1(n_414), .A2(n_1695), .B1(n_1702), .B2(n_1705), .C(n_1706), .Y(n_1701) );
AOI22xp33_ASAP7_75t_L g2018 ( .A1(n_414), .A2(n_491), .B1(n_1998), .B2(n_2001), .Y(n_2018) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx2_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
OR2x2_ASAP7_75t_L g492 ( .A(n_416), .B(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g759 ( .A(n_416), .B(n_558), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_SL g1144 ( .A1(n_416), .A2(n_1145), .B(n_1147), .C(n_1149), .Y(n_1144) );
INVx1_ASAP7_75t_L g426 ( .A(n_417), .Y(n_426) );
INVx1_ASAP7_75t_L g668 ( .A(n_418), .Y(n_668) );
INVx2_ASAP7_75t_L g1019 ( .A(n_418), .Y(n_1019) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g446 ( .A(n_419), .Y(n_446) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_419), .Y(n_485) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_419), .Y(n_660) );
INVx1_ASAP7_75t_L g758 ( .A(n_419), .Y(n_758) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx2_ASAP7_75t_L g432 ( .A(n_420), .Y(n_432) );
AND2x2_ASAP7_75t_L g466 ( .A(n_420), .B(n_438), .Y(n_466) );
INVx1_ASAP7_75t_L g451 ( .A(n_421), .Y(n_451) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g733 ( .A(n_424), .Y(n_733) );
INVx2_ASAP7_75t_SL g931 ( .A(n_424), .Y(n_931) );
AOI222xp33_ASAP7_75t_L g1015 ( .A1(n_424), .A2(n_467), .B1(n_735), .B2(n_1016), .C1(n_1023), .C2(n_1024), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_424), .A2(n_735), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_424), .A2(n_735), .B1(n_1575), .B2(n_1576), .Y(n_1574) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_429), .Y(n_424) );
AND2x2_ASAP7_75t_L g434 ( .A(n_425), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g488 ( .A(n_425), .Y(n_488) );
AND2x2_ASAP7_75t_L g506 ( .A(n_425), .B(n_457), .Y(n_506) );
AND2x4_ASAP7_75t_L g671 ( .A(n_425), .B(n_429), .Y(n_671) );
AND2x4_ASAP7_75t_L g673 ( .A(n_425), .B(n_435), .Y(n_673) );
AND2x2_ASAP7_75t_L g735 ( .A(n_425), .B(n_435), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g781 ( .A(n_425), .B(n_557), .Y(n_781) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_425), .Y(n_1079) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AND2x4_ASAP7_75t_L g459 ( .A(n_427), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g478 ( .A(n_428), .B(n_460), .Y(n_478) );
INVx1_ASAP7_75t_L g1407 ( .A(n_428), .Y(n_1407) );
INVx1_ASAP7_75t_L g1412 ( .A(n_428), .Y(n_1412) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_428), .Y(n_1417) );
INVxp67_ASAP7_75t_L g1076 ( .A(n_429), .Y(n_1076) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g779 ( .A(n_430), .Y(n_779) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g1427 ( .A(n_431), .Y(n_1427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g457 ( .A(n_432), .B(n_437), .Y(n_457) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g785 ( .A(n_435), .Y(n_785) );
INVx1_ASAP7_75t_L g1077 ( .A(n_435), .Y(n_1077) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x6_ASAP7_75t_L g1429 ( .A(n_436), .B(n_1412), .Y(n_1429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g443 ( .A(n_438), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g1567 ( .A(n_442), .Y(n_1567) );
BUFx3_ASAP7_75t_L g1656 ( .A(n_442), .Y(n_1656) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_443), .Y(n_472) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_443), .Y(n_496) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_443), .Y(n_649) );
BUFx2_ASAP7_75t_L g667 ( .A(n_443), .Y(n_667) );
BUFx2_ASAP7_75t_L g738 ( .A(n_443), .Y(n_738) );
INVx2_ASAP7_75t_SL g773 ( .A(n_443), .Y(n_773) );
BUFx3_ASAP7_75t_L g792 ( .A(n_443), .Y(n_792) );
AND2x6_ASAP7_75t_L g1410 ( .A(n_443), .B(n_1411), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1465 ( .A(n_443), .Y(n_1465) );
HB1xp67_ASAP7_75t_L g1709 ( .A(n_443), .Y(n_1709) );
INVx1_ASAP7_75t_L g452 ( .A(n_444), .Y(n_452) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g1031 ( .A(n_446), .Y(n_1031) );
INVx1_ASAP7_75t_L g1318 ( .A(n_446), .Y(n_1318) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_453), .B(n_454), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g1563 ( .A1(n_448), .A2(n_471), .B1(n_971), .B2(n_1549), .C(n_1564), .Y(n_1563) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g938 ( .A(n_449), .Y(n_938) );
INVx1_ASAP7_75t_L g1591 ( .A(n_449), .Y(n_1591) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g763 ( .A(n_450), .Y(n_763) );
BUFx4f_ASAP7_75t_L g959 ( .A(n_450), .Y(n_959) );
INVx1_ASAP7_75t_L g1158 ( .A(n_450), .Y(n_1158) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
OR2x2_ASAP7_75t_L g493 ( .A(n_451), .B(n_452), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_453), .A2(n_564), .B1(n_565), .B2(n_569), .Y(n_563) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_455), .Y(n_925) );
BUFx3_ASAP7_75t_L g973 ( .A(n_455), .Y(n_973) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
INVx2_ASAP7_75t_SL g658 ( .A(n_456), .Y(n_658) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_456), .Y(n_726) );
INVx1_ASAP7_75t_L g796 ( .A(n_456), .Y(n_796) );
INVx1_ASAP7_75t_L g801 ( .A(n_456), .Y(n_801) );
INVx2_ASAP7_75t_L g1408 ( .A(n_456), .Y(n_1408) );
INVx6_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g663 ( .A(n_457), .Y(n_663) );
INVx2_ASAP7_75t_L g768 ( .A(n_457), .Y(n_768) );
AND2x4_ASAP7_75t_L g1415 ( .A(n_457), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1308 ( .A(n_458), .Y(n_1308) );
BUFx2_ASAP7_75t_L g1505 ( .A(n_458), .Y(n_1505) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g665 ( .A(n_459), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_459), .Y(n_727) );
AND2x4_ASAP7_75t_L g807 ( .A(n_459), .B(n_505), .Y(n_807) );
INVx2_ASAP7_75t_SL g942 ( .A(n_459), .Y(n_942) );
HB1xp67_ASAP7_75t_L g1571 ( .A(n_459), .Y(n_1571) );
INVx1_ASAP7_75t_L g1400 ( .A(n_460), .Y(n_1400) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_468), .B1(n_469), .B2(n_479), .C(n_486), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_462), .A2(n_486), .B1(n_637), .B2(n_651), .C(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g1260 ( .A(n_463), .Y(n_1260) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g746 ( .A(n_464), .Y(n_746) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_464), .Y(n_928) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_464), .A2(n_1221), .B1(n_1233), .B2(n_1236), .C(n_1237), .Y(n_1232) );
INVx1_ASAP7_75t_L g1312 ( .A(n_464), .Y(n_1312) );
INVx1_ASAP7_75t_L g1353 ( .A(n_464), .Y(n_1353) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
BUFx3_ASAP7_75t_L g652 ( .A(n_465), .Y(n_652) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_465), .Y(n_798) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_465), .Y(n_1028) );
BUFx4f_ASAP7_75t_L g1227 ( .A(n_465), .Y(n_1227) );
AND2x4_ASAP7_75t_L g1237 ( .A(n_465), .B(n_1079), .Y(n_1237) );
INVx1_ASAP7_75t_L g1704 ( .A(n_465), .Y(n_1704) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_466), .Y(n_476) );
AND2x4_ASAP7_75t_L g495 ( .A(n_467), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g648 ( .A(n_467), .B(n_649), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g1067 ( .A1(n_467), .A2(n_1068), .B(n_1070), .Y(n_1067) );
OAI21xp5_ASAP7_75t_L g1577 ( .A1(n_467), .A2(n_1578), .B(n_1580), .Y(n_1577) );
OAI21xp33_ASAP7_75t_L g1602 ( .A1(n_467), .A2(n_1603), .B(n_1605), .Y(n_1602) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OAI221xp5_ASAP7_75t_L g1590 ( .A1(n_471), .A2(n_1591), .B1(n_1592), .B2(n_1593), .C(n_1594), .Y(n_1590) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g1160 ( .A(n_472), .Y(n_1160) );
A2O1A1Ixp33_ASAP7_75t_SL g1600 ( .A1(n_473), .A2(n_1074), .B(n_1078), .C(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_L g486 ( .A(n_475), .B(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_475), .Y(n_664) );
INVx1_ASAP7_75t_L g921 ( .A(n_475), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_475), .A2(n_649), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
INVx1_ASAP7_75t_L g2015 ( .A(n_475), .Y(n_2015) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g723 ( .A(n_476), .Y(n_723) );
INVx1_ASAP7_75t_L g969 ( .A(n_476), .Y(n_969) );
BUFx6f_ASAP7_75t_L g1234 ( .A(n_476), .Y(n_1234) );
AND2x4_ASAP7_75t_L g1431 ( .A(n_476), .B(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g971 ( .A(n_477), .Y(n_971) );
BUFx2_ASAP7_75t_L g1316 ( .A(n_477), .Y(n_1316) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g654 ( .A(n_478), .Y(n_654) );
INVx2_ASAP7_75t_L g789 ( .A(n_478), .Y(n_789) );
INVx1_ASAP7_75t_L g1235 ( .A(n_478), .Y(n_1235) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_482), .Y(n_743) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g744 ( .A(n_484), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_484), .A2(n_1162), .B1(n_1163), .B2(n_1164), .Y(n_1161) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_485), .Y(n_927) );
BUFx6f_ASAP7_75t_L g974 ( .A(n_485), .Y(n_974) );
AND2x6_ASAP7_75t_L g1419 ( .A(n_485), .B(n_1406), .Y(n_1419) );
INVx1_ASAP7_75t_L g1467 ( .A(n_485), .Y(n_1467) );
INVx1_ASAP7_75t_L g1653 ( .A(n_485), .Y(n_1653) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_486), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_486), .A2(n_913), .B1(n_919), .B2(n_924), .C(n_928), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g962 ( .A1(n_486), .A2(n_928), .B1(n_963), .B2(n_964), .C(n_972), .Y(n_962) );
AOI21xp33_ASAP7_75t_L g1025 ( .A1(n_486), .A2(n_1026), .B(n_1029), .Y(n_1025) );
INVx1_ASAP7_75t_L g1149 ( .A(n_486), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1310 ( .A1(n_486), .A2(n_1311), .B1(n_1313), .B2(n_1314), .C(n_1317), .Y(n_1310) );
AOI221xp5_ASAP7_75t_L g1351 ( .A1(n_486), .A2(n_1352), .B1(n_1354), .B2(n_1355), .C(n_1356), .Y(n_1351) );
AOI221xp5_ASAP7_75t_L g1707 ( .A1(n_486), .A2(n_1352), .B1(n_1698), .B2(n_1708), .C(n_1710), .Y(n_1707) );
AOI221xp5_ASAP7_75t_L g2012 ( .A1(n_486), .A2(n_928), .B1(n_2002), .B2(n_2013), .C(n_2016), .Y(n_2012) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g932 ( .A(n_488), .B(n_785), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_494), .B2(n_495), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_491), .A2(n_629), .B1(n_632), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_491), .A2(n_648), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1711 ( .A1(n_491), .A2(n_495), .B1(n_1694), .B2(n_1697), .Y(n_1711) );
INVx6_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g940 ( .A(n_493), .Y(n_940) );
BUFx2_ASAP7_75t_L g1306 ( .A(n_493), .Y(n_1306) );
INVx1_ASAP7_75t_L g1570 ( .A(n_493), .Y(n_1570) );
INVx1_ASAP7_75t_L g731 ( .A(n_495), .Y(n_731) );
AOI211xp5_ASAP7_75t_L g929 ( .A1(n_495), .A2(n_905), .B(n_930), .C(n_933), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g953 ( .A1(n_495), .A2(n_954), .B(n_955), .Y(n_953) );
HB1xp67_ASAP7_75t_L g1299 ( .A(n_495), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_495), .B(n_1371), .Y(n_1370) );
AOI21xp5_ASAP7_75t_L g2006 ( .A1(n_495), .A2(n_1997), .B(n_2007), .Y(n_2006) );
INVx2_ASAP7_75t_SL g804 ( .A(n_496), .Y(n_804) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_496), .Y(n_1030) );
AOI21xp33_ASAP7_75t_SL g950 ( .A1(n_498), .A2(n_951), .B(n_952), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_498), .A2(n_1349), .B1(n_1350), .B2(n_1372), .Y(n_1348) );
AOI21xp33_ASAP7_75t_L g2003 ( .A1(n_498), .A2(n_2004), .B(n_2005), .Y(n_2003) );
INVx5_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g675 ( .A(n_499), .Y(n_675) );
INVx1_ASAP7_75t_L g915 ( .A(n_499), .Y(n_915) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_499), .Y(n_1239) );
INVx2_ASAP7_75t_L g1263 ( .A(n_499), .Y(n_1263) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx2_ASAP7_75t_L g1062 ( .A(n_500), .Y(n_1062) );
INVx3_ASAP7_75t_L g512 ( .A(n_501), .Y(n_512) );
INVx1_ASAP7_75t_L g820 ( .A(n_502), .Y(n_820) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x6_ASAP7_75t_L g814 ( .A(n_504), .B(n_815), .Y(n_814) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g1036 ( .A(n_506), .Y(n_1036) );
AND4x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_524), .C(n_563), .D(n_571), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_513), .B1(n_514), .B2(n_518), .C(n_519), .Y(n_508) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1023), .C(n_1024), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1113 ( .A1(n_509), .A2(n_519), .B(n_1114), .Y(n_1113) );
AOI221xp5_ASAP7_75t_L g1530 ( .A1(n_509), .A2(n_514), .B1(n_519), .B2(n_1531), .C(n_1532), .Y(n_1530) );
INVx1_ASAP7_75t_L g1585 ( .A(n_509), .Y(n_1585) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
AND2x2_ASAP7_75t_L g842 ( .A(n_510), .B(n_818), .Y(n_842) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g595 ( .A(n_511), .Y(n_595) );
AND2x4_ASAP7_75t_L g514 ( .A(n_512), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g519 ( .A(n_512), .B(n_520), .Y(n_519) );
NAND2x1_ASAP7_75t_SL g593 ( .A(n_512), .B(n_594), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_512), .B(n_597), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_512), .B(n_570), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_514), .A2(n_1062), .B1(n_1073), .B2(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1583 ( .A(n_514), .Y(n_1583) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g613 ( .A(n_517), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_517), .B(n_614), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g1581 ( .A1(n_519), .A2(n_1575), .B1(n_1576), .B2(n_1582), .C(n_1584), .Y(n_1581) );
AOI221xp5_ASAP7_75t_L g1630 ( .A1(n_519), .A2(n_1582), .B1(n_1584), .B2(n_1608), .C(n_1609), .Y(n_1630) );
INVx1_ASAP7_75t_L g1437 ( .A(n_520), .Y(n_1437) );
HB1xp67_ASAP7_75t_L g1527 ( .A(n_520), .Y(n_1527) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_521), .Y(n_534) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_521), .Y(n_554) );
BUFx3_ASAP7_75t_L g570 ( .A(n_521), .Y(n_570) );
BUFx3_ASAP7_75t_L g828 ( .A(n_521), .Y(n_828) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_521), .B(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1474 ( .A(n_521), .Y(n_1474) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
AOI33xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_528), .A3(n_535), .B1(n_545), .B2(n_549), .B3(n_555), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g1053 ( .A1(n_525), .A2(n_1037), .B1(n_1054), .B2(n_1062), .Y(n_1053) );
AOI322xp5_ASAP7_75t_L g1105 ( .A1(n_525), .A2(n_555), .A3(n_1089), .B1(n_1106), .B2(n_1108), .C1(n_1109), .C2(n_1112), .Y(n_1105) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
OR2x6_ASAP7_75t_L g788 ( .A(n_526), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g816 ( .A(n_526), .Y(n_816) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_526), .Y(n_1171) );
AND2x4_ASAP7_75t_L g1470 ( .A(n_526), .B(n_527), .Y(n_1470) );
INVx1_ASAP7_75t_L g865 ( .A(n_527), .Y(n_865) );
INVx1_ASAP7_75t_L g837 ( .A(n_529), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_529), .A2(n_1044), .B1(n_1045), .B2(n_1046), .Y(n_1043) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g847 ( .A(n_530), .B(n_568), .Y(n_847) );
BUFx2_ASAP7_75t_L g1472 ( .A(n_530), .Y(n_1472) );
INVx3_ASAP7_75t_L g1553 ( .A(n_530), .Y(n_1553) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g1046 ( .A(n_533), .Y(n_1046) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g1526 ( .A(n_536), .Y(n_1526) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_537), .Y(n_577) );
AND2x2_ASAP7_75t_L g870 ( .A(n_537), .B(n_568), .Y(n_870) );
INVx1_ASAP7_75t_L g1049 ( .A(n_537), .Y(n_1049) );
INVx1_ASAP7_75t_L g1056 ( .A(n_537), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g1107 ( .A(n_537), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1446 ( .A(n_537), .B(n_1447), .Y(n_1446) );
BUFx6f_ASAP7_75t_L g1477 ( .A(n_537), .Y(n_1477) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g704 ( .A(n_541), .Y(n_704) );
BUFx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g566 ( .A(n_542), .B(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g548 ( .A(n_543), .Y(n_548) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_543), .Y(n_908) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_544), .Y(n_623) );
INVx1_ASAP7_75t_L g857 ( .A(n_544), .Y(n_857) );
INVx1_ASAP7_75t_L g1451 ( .A(n_544), .Y(n_1451) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_547), .A2(n_1248), .B1(n_1250), .B2(n_1282), .Y(n_1287) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g901 ( .A(n_548), .Y(n_901) );
INVx2_ASAP7_75t_L g1003 ( .A(n_548), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_548), .B(n_567), .Y(n_1103) );
INVx2_ASAP7_75t_L g1137 ( .A(n_548), .Y(n_1137) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g574 ( .A(n_552), .Y(n_574) );
INVx2_ASAP7_75t_SL g821 ( .A(n_552), .Y(n_821) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_554), .B(n_567), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_555), .A2(n_567), .B1(n_1041), .B2(n_1047), .Y(n_1040) );
INVx1_ASAP7_75t_L g1222 ( .A(n_555), .Y(n_1222) );
INVx2_ASAP7_75t_L g1395 ( .A(n_555), .Y(n_1395) );
AOI33xp33_ASAP7_75t_L g1468 ( .A1(n_555), .A2(n_1469), .A3(n_1471), .B1(n_1475), .B2(n_1482), .B3(n_1483), .Y(n_1468) );
INVx6_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx5_ASAP7_75t_L g639 ( .A(n_556), .Y(n_639) );
OR2x6_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g567 ( .A(n_558), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g839 ( .A(n_559), .Y(n_839) );
NAND2x1p5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g1440 ( .A(n_560), .Y(n_1440) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g605 ( .A(n_561), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_565), .A2(n_569), .B1(n_585), .B2(n_586), .Y(n_584) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_566), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
BUFx2_ASAP7_75t_L g883 ( .A(n_566), .Y(n_883) );
BUFx2_ASAP7_75t_L g982 ( .A(n_566), .Y(n_982) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_566), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_566), .A2(n_689), .B1(n_1305), .B2(n_1327), .Y(n_1326) );
BUFx2_ASAP7_75t_L g1376 ( .A(n_566), .Y(n_1376) );
BUFx2_ASAP7_75t_L g1517 ( .A(n_566), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1626 ( .A1(n_566), .A2(n_569), .B1(n_1597), .B2(n_1627), .Y(n_1626) );
BUFx2_ASAP7_75t_L g1978 ( .A(n_566), .Y(n_1978) );
AND2x6_ASAP7_75t_L g569 ( .A(n_567), .B(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g573 ( .A(n_567), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g576 ( .A(n_567), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g685 ( .A(n_567), .B(n_577), .Y(n_685) );
AND2x2_ASAP7_75t_L g986 ( .A(n_567), .B(n_577), .Y(n_986) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_567), .B(n_577), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_567), .B(n_821), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_567), .B(n_577), .Y(n_1543) );
INVx2_ASAP7_75t_L g827 ( .A(n_568), .Y(n_827) );
BUFx2_ASAP7_75t_L g689 ( .A(n_569), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_569), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_569), .A2(n_957), .B1(n_981), .B2(n_982), .Y(n_980) );
INVx1_ASAP7_75t_SL g1120 ( .A(n_569), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_569), .A2(n_1267), .B1(n_1268), .B2(n_1269), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_569), .A2(n_1368), .B1(n_1376), .B2(n_1377), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_569), .A2(n_883), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
AOI22xp33_ASAP7_75t_L g1679 ( .A1(n_569), .A2(n_982), .B1(n_1680), .B2(n_1681), .Y(n_1679) );
AOI22xp33_ASAP7_75t_L g1976 ( .A1(n_569), .A2(n_1977), .B1(n_1978), .B2(n_1979), .Y(n_1976) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_575), .B2(n_576), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_573), .A2(n_576), .B1(n_588), .B2(n_589), .Y(n_587) );
BUFx2_ASAP7_75t_L g683 ( .A(n_573), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_573), .A2(n_685), .B1(n_886), .B2(n_887), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_573), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_573), .A2(n_685), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_573), .A2(n_986), .B1(n_1366), .B2(n_1379), .Y(n_1378) );
AOI21xp5_ASAP7_75t_L g1545 ( .A1(n_573), .A2(n_1546), .B(n_1547), .Y(n_1545) );
AOI22xp33_ASAP7_75t_L g1682 ( .A1(n_573), .A2(n_685), .B1(n_1683), .B2(n_1684), .Y(n_1682) );
AOI22xp33_ASAP7_75t_L g1980 ( .A1(n_573), .A2(n_1543), .B1(n_1981), .B2(n_1982), .Y(n_1980) );
XNOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_640), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .C(n_601), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g691 ( .A(n_592), .Y(n_691) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g1274 ( .A(n_593), .Y(n_1274) );
NAND2x1p5_ASAP7_75t_L g2057 ( .A(n_594), .B(n_2058), .Y(n_2057) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx4f_ASAP7_75t_L g693 ( .A(n_596), .Y(n_693) );
BUFx4f_ASAP7_75t_L g1381 ( .A(n_596), .Y(n_1381) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x6_ASAP7_75t_L g844 ( .A(n_598), .B(n_819), .Y(n_844) );
BUFx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx3_ASAP7_75t_L g889 ( .A(n_600), .Y(n_889) );
BUFx2_ASAP7_75t_L g988 ( .A(n_600), .Y(n_988) );
OAI33xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_606), .A3(n_616), .B1(n_625), .B2(n_631), .B3(n_638), .Y(n_601) );
OAI33xp33_ASAP7_75t_L g1686 ( .A1(n_602), .A2(n_638), .A3(n_1687), .B1(n_1690), .B2(n_1693), .B3(n_1696), .Y(n_1686) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI33xp33_ASAP7_75t_L g694 ( .A1(n_603), .A2(n_695), .A3(n_701), .B1(n_705), .B2(n_710), .B3(n_713), .Y(n_694) );
OAI33xp33_ASAP7_75t_L g890 ( .A1(n_603), .A2(n_638), .A3(n_891), .B1(n_895), .B2(n_902), .B3(n_910), .Y(n_890) );
OAI33xp33_ASAP7_75t_L g989 ( .A1(n_603), .A2(n_638), .A3(n_990), .B1(n_997), .B2(n_1001), .B3(n_1004), .Y(n_989) );
OAI33xp33_ASAP7_75t_L g1197 ( .A1(n_603), .A2(n_1198), .A3(n_1205), .B1(n_1212), .B2(n_1219), .B3(n_1222), .Y(n_1197) );
OAI33xp33_ASAP7_75t_L g1275 ( .A1(n_603), .A2(n_638), .A3(n_1276), .B1(n_1280), .B2(n_1287), .B3(n_1288), .Y(n_1275) );
OAI33xp33_ASAP7_75t_L g1329 ( .A1(n_603), .A2(n_1222), .A3(n_1330), .B1(n_1333), .B2(n_1338), .B3(n_1339), .Y(n_1329) );
OAI33xp33_ASAP7_75t_L g1382 ( .A1(n_603), .A2(n_1383), .A3(n_1387), .B1(n_1392), .B2(n_1393), .B3(n_1395), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_603), .A2(n_638), .B1(n_1548), .B2(n_1554), .Y(n_1547) );
OAI33xp33_ASAP7_75t_L g1611 ( .A1(n_603), .A2(n_1395), .A3(n_1612), .B1(n_1616), .B2(n_1618), .B3(n_1622), .Y(n_1611) );
INVx1_ASAP7_75t_L g1986 ( .A(n_603), .Y(n_1986) );
INVx1_ASAP7_75t_L g1447 ( .A(n_605), .Y(n_1447) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_610), .B1(n_611), .B2(n_615), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_607), .A2(n_632), .B1(n_633), .B2(n_637), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g1687 ( .A1(n_607), .A2(n_611), .B1(n_1688), .B2(n_1689), .Y(n_1687) );
OAI22xp33_ASAP7_75t_L g1696 ( .A1(n_607), .A2(n_611), .B1(n_1697), .B2(n_1698), .Y(n_1696) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g1006 ( .A(n_609), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_609), .A2(n_612), .B1(n_1022), .B2(n_1052), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_609), .A2(n_612), .B1(n_1060), .B2(n_1061), .Y(n_1059) );
OAI22xp5_ASAP7_75t_SL g1139 ( .A1(n_609), .A2(n_633), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
BUFx2_ASAP7_75t_L g2000 ( .A(n_609), .Y(n_2000) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_611), .A2(n_963), .B1(n_976), .B2(n_1005), .Y(n_1004) );
BUFx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g867 ( .A(n_613), .Y(n_867) );
BUFx2_ASAP7_75t_L g995 ( .A(n_613), .Y(n_995) );
INVx2_ASAP7_75t_L g1204 ( .A(n_613), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_621), .B1(n_622), .B2(n_624), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g1690 ( .A1(n_617), .A2(n_1042), .B1(n_1691), .B2(n_1692), .Y(n_1690) );
BUFx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_618), .A2(n_998), .B1(n_999), .B2(n_1000), .Y(n_997) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g1208 ( .A(n_619), .Y(n_1208) );
HB1xp67_ASAP7_75t_L g1335 ( .A(n_619), .Y(n_1335) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g628 ( .A(n_620), .Y(n_628) );
BUFx2_ASAP7_75t_L g904 ( .A(n_620), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_622), .A2(n_626), .B1(n_629), .B2(n_630), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_622), .A2(n_832), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVx2_ASAP7_75t_L g1524 ( .A(n_622), .Y(n_1524) );
INVx4_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g708 ( .A(n_623), .Y(n_708) );
INVx2_ASAP7_75t_SL g834 ( .A(n_623), .Y(n_834) );
INVx2_ASAP7_75t_SL g1042 ( .A(n_623), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_623), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_626), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_626), .A2(n_706), .B1(n_707), .B2(n_709), .Y(n_705) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g1283 ( .A(n_627), .Y(n_1283) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g833 ( .A(n_628), .Y(n_833) );
OAI22xp5_ASAP7_75t_SL g1219 ( .A1(n_633), .A2(n_861), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
OAI22xp33_ASAP7_75t_L g1288 ( .A1(n_633), .A2(n_1247), .B1(n_1261), .B2(n_1277), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1330 ( .A1(n_633), .A2(n_861), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
OAI22xp33_ASAP7_75t_L g1339 ( .A1(n_633), .A2(n_834), .B1(n_1313), .B2(n_1321), .Y(n_1339) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g912 ( .A(n_634), .Y(n_912) );
INVx1_ASAP7_75t_L g1385 ( .A(n_634), .Y(n_1385) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx3_ASAP7_75t_L g699 ( .A(n_635), .Y(n_699) );
BUFx3_ASAP7_75t_L g1394 ( .A(n_635), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g714 ( .A(n_638), .Y(n_714) );
OAI33xp33_ASAP7_75t_L g1984 ( .A1(n_638), .A2(n_1985), .A3(n_1987), .B1(n_1990), .B2(n_1996), .B3(n_1999), .Y(n_1984) );
CKINVDCx8_ASAP7_75t_R g638 ( .A(n_639), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B1(n_674), .B2(n_675), .Y(n_640) );
INVx1_ASAP7_75t_SL g749 ( .A(n_641), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g1699 ( .A1(n_641), .A2(n_1263), .B1(n_1700), .B2(n_1712), .Y(n_1699) );
INVx5_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI31xp33_ASAP7_75t_L g1659 ( .A1(n_642), .A2(n_1660), .A3(n_1665), .B(n_1672), .Y(n_1659) );
AOI221x1_ASAP7_75t_SL g2033 ( .A1(n_642), .A2(n_1399), .B1(n_2034), .B2(n_2046), .C(n_2069), .Y(n_2033) );
BUFx8_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
OAI31xp33_ASAP7_75t_L g822 ( .A1(n_643), .A2(n_823), .A3(n_845), .B(n_868), .Y(n_822) );
INVx2_ASAP7_75t_L g1244 ( .A(n_643), .Y(n_1244) );
AOI31xp33_ASAP7_75t_L g1296 ( .A1(n_643), .A2(n_1297), .A3(n_1310), .B(n_1319), .Y(n_1296) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_650), .C(n_661), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_648), .A2(n_1213), .B1(n_1226), .B2(n_1228), .C(n_1229), .Y(n_1225) );
BUFx2_ASAP7_75t_L g729 ( .A(n_649), .Y(n_729) );
INVx1_ASAP7_75t_L g935 ( .A(n_649), .Y(n_935) );
INVx1_ASAP7_75t_L g966 ( .A(n_649), .Y(n_966) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g740 ( .A(n_654), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_654), .A2(n_1127), .B1(n_1132), .B2(n_1157), .C(n_1159), .Y(n_1156) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g1155 ( .A(n_659), .Y(n_1155) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx3_ASAP7_75t_L g805 ( .A(n_660), .Y(n_805) );
INVx1_ASAP7_75t_L g1358 ( .A(n_660), .Y(n_1358) );
INVx1_ASAP7_75t_L g1604 ( .A(n_660), .Y(n_1604) );
A2O1A1Ixp33_ASAP7_75t_L g1573 ( .A1(n_663), .A2(n_664), .B(n_1078), .C(n_1544), .Y(n_1573) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_664), .Y(n_739) );
INVx1_ASAP7_75t_L g1169 ( .A(n_665), .Y(n_1169) );
INVx1_ASAP7_75t_L g1579 ( .A(n_668), .Y(n_1579) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx4_ASAP7_75t_L g1230 ( .A(n_671), .Y(n_1230) );
INVx1_ASAP7_75t_SL g2008 ( .A(n_671), .Y(n_2008) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g1231 ( .A(n_673), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1606 ( .A1(n_673), .A2(n_1607), .B1(n_1608), .B2(n_1609), .Y(n_1606) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_675), .A2(n_716), .B(n_717), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g1494 ( .A1(n_675), .A2(n_1495), .B(n_1496), .Y(n_1494) );
INVx1_ASAP7_75t_L g874 ( .A(n_676), .Y(n_874) );
XOR2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_750), .Y(n_676) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_715), .Y(n_679) );
NOR3xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_690), .C(n_694), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_683), .A2(n_685), .B1(n_1307), .B2(n_1325), .Y(n_1324) );
AOI21xp5_ASAP7_75t_L g1610 ( .A1(n_683), .A2(n_1598), .B(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_689), .A2(n_1516), .B1(n_1517), .B2(n_1518), .Y(n_1515) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_696), .A2(n_699), .B1(n_711), .B2(n_712), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g1987 ( .A1(n_696), .A2(n_994), .B1(n_1988), .B2(n_1989), .Y(n_1987) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx3_ASAP7_75t_L g859 ( .A(n_699), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_699), .A2(n_1130), .B1(n_1131), .B2(n_1132), .Y(n_1129) );
AOI221xp5_ASAP7_75t_SL g718 ( .A1(n_706), .A2(n_719), .B1(n_728), .B2(n_730), .C(n_732), .Y(n_718) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g999 ( .A(n_708), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_712), .A2(n_737), .B1(n_741), .B2(n_745), .C(n_747), .Y(n_736) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI33xp33_ASAP7_75t_L g1520 ( .A1(n_714), .A2(n_1521), .A3(n_1523), .B1(n_1525), .B2(n_1528), .B3(n_1529), .Y(n_1520) );
AOI31xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_736), .A3(n_748), .B(n_749), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g2039 ( .A1(n_720), .A2(n_1424), .B1(n_1429), .B2(n_2040), .C1(n_2041), .C2(n_2042), .Y(n_2039) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g1074 ( .A(n_726), .Y(n_1074) );
INVx4_ASAP7_75t_L g1146 ( .A(n_726), .Y(n_1146) );
AOI211xp5_ASAP7_75t_SL g1497 ( .A1(n_730), .A2(n_1498), .B(n_1499), .C(n_1500), .Y(n_1497) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g1506 ( .A1(n_745), .A2(n_747), .B1(n_1507), .B2(n_1508), .C(n_1509), .Y(n_1506) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
AOI31xp33_ASAP7_75t_L g1496 ( .A1(n_749), .A2(n_1497), .A3(n_1506), .B(n_1510), .Y(n_1496) );
AND3x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_812), .C(n_822), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_774), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_764), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_760), .B2(n_761), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_755), .A2(n_770), .B1(n_830), .B2(n_834), .C(n_835), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1638 ( .A1(n_756), .A2(n_771), .B1(n_1639), .B2(n_1640), .Y(n_1638) );
CKINVDCx6p67_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
OR2x6_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx2_ASAP7_75t_L g793 ( .A(n_758), .Y(n_793) );
OR2x6_ASAP7_75t_L g762 ( .A(n_759), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g769 ( .A(n_759), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1641 ( .A1(n_761), .A2(n_766), .B1(n_1642), .B2(n_1643), .Y(n_1641) );
CKINVDCx6p67_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
BUFx3_ASAP7_75t_L g1082 ( .A(n_763), .Y(n_1082) );
INVx1_ASAP7_75t_L g1091 ( .A(n_763), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_770), .B2(n_771), .Y(n_764) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .Y(n_766) );
INVx2_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g1252 ( .A(n_768), .Y(n_1252) );
INVx1_ASAP7_75t_L g2017 ( .A(n_768), .Y(n_2017) );
AND2x2_ASAP7_75t_L g771 ( .A(n_769), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_773), .Y(n_1085) );
INVx1_ASAP7_75t_L g1258 ( .A(n_773), .Y(n_1258) );
NAND3xp33_ASAP7_75t_SL g774 ( .A(n_775), .B(n_786), .C(n_808), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_782), .B2(n_783), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_776), .A2(n_782), .B1(n_841), .B2(n_843), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1645 ( .A1(n_777), .A2(n_783), .B1(n_1646), .B2(n_1647), .Y(n_1645) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2x1p5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx2_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
OR2x6_ASAP7_75t_L g784 ( .A(n_781), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g811 ( .A(n_781), .Y(n_811) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AOI33xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_790), .A3(n_794), .B1(n_799), .B2(n_802), .B3(n_806), .Y(n_786) );
AOI33xp33_ASAP7_75t_L g1460 ( .A1(n_787), .A2(n_806), .A3(n_1461), .B1(n_1462), .B2(n_1463), .B3(n_1464), .Y(n_1460) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g1649 ( .A(n_788), .Y(n_1649) );
INVx2_ASAP7_75t_L g2071 ( .A(n_788), .Y(n_2071) );
INVx1_ASAP7_75t_L g1087 ( .A(n_789), .Y(n_1087) );
BUFx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_SL g923 ( .A(n_792), .Y(n_923) );
BUFx2_ASAP7_75t_L g936 ( .A(n_793), .Y(n_936) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g1562 ( .A(n_796), .Y(n_1562) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_798), .B(n_811), .Y(n_810) );
BUFx2_ASAP7_75t_SL g1148 ( .A(n_798), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_798), .Y(n_1422) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx4f_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI33xp33_ASAP7_75t_L g1648 ( .A1(n_807), .A2(n_1649), .A3(n_1650), .B1(n_1651), .B2(n_1654), .B3(n_1655), .Y(n_1648) );
INVx4_ASAP7_75t_L g2076 ( .A(n_807), .Y(n_2076) );
NAND3xp33_ASAP7_75t_SL g1644 ( .A(n_808), .B(n_1645), .C(n_1648), .Y(n_1644) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_814), .B(n_1658), .Y(n_1657) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx2_ASAP7_75t_L g1038 ( .A(n_816), .Y(n_1038) );
AOI211xp5_ASAP7_75t_L g1065 ( .A1(n_816), .A2(n_1066), .B(n_1094), .C(n_1104), .Y(n_1065) );
INVx1_ASAP7_75t_L g2063 ( .A(n_817), .Y(n_2063) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_821), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g866 ( .A(n_819), .B(n_867), .Y(n_866) );
OR2x6_ASAP7_75t_L g2049 ( .A(n_819), .B(n_867), .Y(n_2049) );
INVx1_ASAP7_75t_L g2058 ( .A(n_819), .Y(n_2058) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx8_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI222xp33_ASAP7_75t_L g2062 ( .A1(n_825), .A2(n_847), .B1(n_2037), .B2(n_2063), .C1(n_2064), .C2(n_2065), .Y(n_2062) );
AND2x4_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .Y(n_825) );
AND2x4_ASAP7_75t_L g872 ( .A(n_826), .B(n_856), .Y(n_872) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
BUFx6f_ASAP7_75t_L g1558 ( .A(n_828), .Y(n_1558) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_830), .A2(n_1388), .B1(n_1389), .B2(n_1391), .Y(n_1387) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_830), .A2(n_1361), .B1(n_1371), .B2(n_1389), .Y(n_1392) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_832), .A2(n_954), .B1(n_977), .B2(n_1002), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1693 ( .A1(n_832), .A2(n_1002), .B1(n_1694), .B2(n_1695), .Y(n_1693) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_SL g851 ( .A(n_833), .Y(n_851) );
INVx2_ASAP7_75t_L g897 ( .A(n_833), .Y(n_897) );
INVx2_ASAP7_75t_L g1214 ( .A(n_833), .Y(n_1214) );
OAI22xp5_ASAP7_75t_L g1333 ( .A1(n_834), .A2(n_1334), .B1(n_1336), .B2(n_1337), .Y(n_1333) );
OAI221xp5_ASAP7_75t_L g1554 ( .A1(n_834), .A2(n_851), .B1(n_1555), .B2(n_1556), .C(n_1557), .Y(n_1554) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1664 ( .A1(n_841), .A2(n_843), .B1(n_1646), .B2(n_1647), .Y(n_1664) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
CKINVDCx11_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
CKINVDCx6p67_ASAP7_75t_R g846 ( .A(n_847), .Y(n_846) );
OAI22xp5_ASAP7_75t_SL g848 ( .A1(n_849), .A2(n_850), .B1(n_852), .B2(n_853), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_850), .A2(n_861), .B1(n_1298), .B2(n_1320), .Y(n_1338) );
BUFx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g1618 ( .A1(n_851), .A2(n_1619), .B1(n_1620), .B2(n_1621), .Y(n_1618) );
OAI22xp5_ASAP7_75t_L g1669 ( .A1(n_853), .A2(n_1334), .B1(n_1670), .B2(n_1671), .Y(n_1669) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g1218 ( .A(n_857), .Y(n_1218) );
OAI221xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_861), .B2(n_863), .C(n_864), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_859), .A2(n_892), .B1(n_893), .B2(n_894), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g1666 ( .A1(n_859), .A2(n_861), .B1(n_864), .B2(n_1667), .C(n_1668), .Y(n_1666) );
BUFx2_ASAP7_75t_L g893 ( .A(n_861), .Y(n_893) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g1615 ( .A(n_867), .Y(n_1615) );
INVx3_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g2066 ( .A1(n_870), .A2(n_872), .B1(n_2067), .B2(n_2068), .Y(n_2066) );
INVx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_945), .B1(n_1175), .B2(n_1177), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_877), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_877), .A2(n_945), .B1(n_946), .B2(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g878 ( .A(n_879), .B(n_914), .Y(n_878) );
NOR3xp33_ASAP7_75t_SL g879 ( .A(n_880), .B(n_888), .C(n_890), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_885), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_884), .A2(n_886), .B1(n_938), .B2(n_939), .C(n_941), .Y(n_937) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_893), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_893), .A2(n_1354), .B1(n_1360), .B2(n_1394), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_895) );
OAI221xp5_ASAP7_75t_L g1661 ( .A1(n_897), .A2(n_1058), .B1(n_1639), .B2(n_1640), .C(n_1662), .Y(n_1661) );
INVx2_ASAP7_75t_SL g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g1050 ( .A(n_901), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_905), .B1(n_906), .B2(n_909), .Y(n_902) );
BUFx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g1136 ( .A(n_904), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g1548 ( .A1(n_906), .A2(n_1135), .B1(n_1549), .B2(n_1550), .C(n_1551), .Y(n_1548) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx3_ASAP7_75t_L g1390 ( .A(n_908), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g1616 ( .A1(n_908), .A2(n_1207), .B1(n_1593), .B2(n_1617), .Y(n_1616) );
INVx2_ASAP7_75t_SL g1995 ( .A(n_908), .Y(n_1995) );
INVx2_ASAP7_75t_L g2051 ( .A(n_908), .Y(n_2051) );
OAI22xp33_ASAP7_75t_L g1622 ( .A1(n_912), .A2(n_1131), .B1(n_1623), .B2(n_1624), .Y(n_1622) );
AOI21xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B(n_917), .Y(n_914) );
AOI31xp33_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_929), .A3(n_943), .B(n_944), .Y(n_917) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_922), .A2(n_1134), .B1(n_1141), .B2(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_936), .A2(n_1138), .B1(n_1140), .B2(n_1146), .Y(n_1145) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx2_ASAP7_75t_L g1069 ( .A(n_940), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_940), .Y(n_1154) );
INVx2_ASAP7_75t_L g1167 ( .A(n_940), .Y(n_1167) );
OAI221xp5_ASAP7_75t_L g1596 ( .A1(n_941), .A2(n_1071), .B1(n_1569), .B2(n_1597), .C(n_1598), .Y(n_1596) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
AOI31xp33_ASAP7_75t_L g952 ( .A1(n_944), .A2(n_953), .A3(n_962), .B(n_975), .Y(n_952) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx2_ASAP7_75t_L g1176 ( .A(n_946), .Y(n_1176) );
XNOR2x1_ASAP7_75t_L g946 ( .A(n_947), .B(n_1008), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
XNOR2x1_ASAP7_75t_L g948 ( .A(n_949), .B(n_1007), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_978), .Y(n_949) );
OAI211xp5_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_958), .B(n_960), .C(n_961), .Y(n_956) );
OAI221xp5_ASAP7_75t_L g1568 ( .A1(n_958), .A2(n_1540), .B1(n_1546), .B2(n_1569), .C(n_1571), .Y(n_1568) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_959), .Y(n_1071) );
INVx1_ASAP7_75t_L g1304 ( .A(n_959), .Y(n_1304) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
NOR3xp33_ASAP7_75t_SL g978 ( .A(n_979), .B(n_987), .C(n_989), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_983), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g1628 ( .A1(n_986), .A2(n_1062), .B1(n_1601), .B2(n_1629), .Y(n_1628) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_993), .B1(n_994), .B2(n_996), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx2_ASAP7_75t_L g1131 ( .A(n_992), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1276 ( .A1(n_994), .A2(n_1277), .B1(n_1278), .B2(n_1279), .Y(n_1276) );
OAI22xp33_ASAP7_75t_L g1999 ( .A1(n_994), .A2(n_2000), .B1(n_2001), .B2(n_2002), .Y(n_1999) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1996 ( .A1(n_999), .A2(n_1992), .B1(n_1997), .B2(n_1998), .Y(n_1996) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1003), .Y(n_1286) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
OAI22x1_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1115), .B2(n_1174), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
XNOR2x1_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1064), .Y(n_1010) );
XNOR2x1_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1013), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1039), .Y(n_1013) );
AOI31xp33_ASAP7_75t_SL g1014 ( .A1(n_1015), .A2(n_1025), .A3(n_1032), .B(n_1038), .Y(n_1014) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1019), .Y(n_1302) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1028), .Y(n_1253) );
INVxp67_ASAP7_75t_L g1163 ( .A(n_1030), .Y(n_1163) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1031), .Y(n_1367) );
AOI22xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1034), .B1(n_1035), .B2(n_1037), .Y(n_1032) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1038), .Y(n_1349) );
NAND3xp33_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1053), .C(n_1063), .Y(n_1039) );
INVx2_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g1541 ( .A1(n_1062), .A2(n_1542), .B1(n_1543), .B2(n_1544), .Y(n_1541) );
NAND4xp25_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1072), .C(n_1080), .D(n_1088), .Y(n_1066) );
OAI211xp5_ASAP7_75t_L g2009 ( .A1(n_1071), .A2(n_1979), .B(n_2010), .C(n_2011), .Y(n_2009) );
A2O1A1Ixp33_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B(n_1075), .C(n_1078), .Y(n_1072) );
BUFx3_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OAI211xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B(n_1083), .C(n_1084), .Y(n_1080) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
OAI211xp5_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1090), .B(n_1092), .C(n_1093), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g2072 ( .A1(n_1090), .A2(n_1167), .B1(n_2073), .B2(n_2074), .C(n_2075), .Y(n_2072) );
OAI221xp5_ASAP7_75t_L g2077 ( .A1(n_1090), .A2(n_1153), .B1(n_2064), .B2(n_2065), .C(n_2078), .Y(n_2077) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1096), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_1096), .A2(n_1101), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
AOI22xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1101), .B1(n_1102), .B2(n_1103), .Y(n_1099) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1101), .Y(n_1142) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1103), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_1103), .A2(n_1112), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1113), .Y(n_1104) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1115), .Y(n_1174) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1116), .Y(n_1172) );
NAND3xp33_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1123), .C(n_1143), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1121), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1125), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_1128), .A2(n_1130), .B1(n_1153), .B2(n_1155), .Y(n_1152) );
OAI22xp33_ASAP7_75t_L g1383 ( .A1(n_1131), .A2(n_1384), .B1(n_1385), .B2(n_1386), .Y(n_1383) );
OAI22xp33_ASAP7_75t_L g1612 ( .A1(n_1131), .A2(n_1592), .B1(n_1613), .B2(n_1614), .Y(n_1612) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1135), .B1(n_1137), .B2(n_1138), .Y(n_1133) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1137), .Y(n_1211) );
OAI31xp33_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1150), .A3(n_1151), .B(n_1170), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_1152), .A2(n_1156), .B1(n_1161), .B2(n_1165), .Y(n_1151) );
OAI21xp5_ASAP7_75t_SL g1501 ( .A1(n_1153), .A2(n_1502), .B(n_1503), .Y(n_1501) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_1157), .A2(n_1166), .B1(n_1167), .B2(n_1168), .C(n_1169), .Y(n_1165) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1157), .Y(n_1504) );
BUFx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI221xp5_ASAP7_75t_L g1365 ( .A1(n_1163), .A2(n_1366), .B1(n_1367), .B2(n_1368), .C(n_1369), .Y(n_1365) );
AOI22xp5_ASAP7_75t_L g1223 ( .A1(n_1170), .A2(n_1224), .B1(n_1239), .B2(n_1240), .Y(n_1223) );
OAI31xp33_ASAP7_75t_SL g1559 ( .A1(n_1170), .A2(n_1560), .A3(n_1565), .B(n_1572), .Y(n_1559) );
INVx2_ASAP7_75t_L g2019 ( .A(n_1170), .Y(n_2019) );
CKINVDCx8_ASAP7_75t_R g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1177), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
OAI21xp5_ASAP7_75t_L g1487 ( .A1(n_1182), .A2(n_1488), .B(n_1489), .Y(n_1487) );
XOR2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1289), .Y(n_1182) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
XNOR2xp5_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1241), .Y(n_1184) );
XNOR2x1_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1223), .Y(n_1187) );
NOR3xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1196), .C(n_1197), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1193), .Y(n_1189) );
OAI22xp33_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1200), .B1(n_1203), .B2(n_1204), .Y(n_1198) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
INVx2_ASAP7_75t_SL g1277 ( .A(n_1201), .Y(n_1277) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_1202), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1207), .B1(n_1209), .B2(n_1210), .Y(n_1205) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
OAI22xp5_ASAP7_75t_SL g1212 ( .A1(n_1213), .A2(n_1214), .B1(n_1215), .B2(n_1216), .Y(n_1212) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1232), .C(n_1238), .Y(n_1224) );
BUFx2_ASAP7_75t_L g1315 ( .A(n_1227), .Y(n_1315) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1230), .Y(n_1607) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1235), .Y(n_1594) );
AOI221xp5_ASAP7_75t_L g1256 ( .A1(n_1237), .A2(n_1257), .B1(n_1259), .B2(n_1260), .C(n_1261), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1264), .Y(n_1242) );
AOI22xp5_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1245), .B1(n_1262), .B2(n_1263), .Y(n_1243) );
NAND3xp33_ASAP7_75t_SL g1245 ( .A(n_1246), .B(n_1249), .C(n_1256), .Y(n_1245) );
AOI21xp5_ASAP7_75t_L g1294 ( .A1(n_1263), .A2(n_1295), .B(n_1296), .Y(n_1294) );
NOR3xp33_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1273), .C(n_1275), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1270), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1282), .B1(n_1284), .B2(n_1285), .Y(n_1280) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx2_ASAP7_75t_L g1992 ( .A(n_1283), .Y(n_1992) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1291), .B1(n_1341), .B2(n_1342), .Y(n_1289) );
INVx2_ASAP7_75t_SL g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1322), .Y(n_1293) );
AOI211xp5_ASAP7_75t_L g1297 ( .A1(n_1298), .A2(n_1299), .B(n_1300), .C(n_1309), .Y(n_1297) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
OAI221xp5_ASAP7_75t_L g1303 ( .A1(n_1304), .A2(n_1305), .B1(n_1306), .B2(n_1307), .C(n_1308), .Y(n_1303) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
NOR3xp33_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1328), .C(n_1329), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1326), .Y(n_1323) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1344), .B1(n_1396), .B2(n_1486), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
XNOR2x1_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1347), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1373), .Y(n_1347) );
NAND5xp2_ASAP7_75t_SL g1350 ( .A(n_1351), .B(n_1359), .C(n_1362), .D(n_1365), .E(n_1370), .Y(n_1350) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
NOR3xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1380), .C(n_1382), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1378), .Y(n_1374) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1390), .Y(n_1620) );
INVxp67_ASAP7_75t_SL g1396 ( .A(n_1397), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g1486 ( .A(n_1397), .Y(n_1486) );
INVx2_ASAP7_75t_L g1485 ( .A(n_1398), .Y(n_1485) );
AO211x2_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1401), .B(n_1433), .C(n_1459), .Y(n_1398) );
NAND4xp25_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1413), .C(n_1420), .D(n_1430), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .B1(n_1409), .B2(n_1410), .Y(n_1402) );
HB1xp67_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g2043 ( .A1(n_1405), .A2(n_1410), .B1(n_2044), .B2(n_2045), .Y(n_2043) );
AND2x4_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1408), .Y(n_1405) );
INVx1_ASAP7_75t_SL g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1411), .Y(n_1432) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_1414), .A2(n_1415), .B1(n_1418), .B2(n_1419), .Y(n_1413) );
AOI22xp33_ASAP7_75t_SL g1453 ( .A1(n_1414), .A2(n_1454), .B1(n_1455), .B2(n_1456), .Y(n_1453) );
AOI22xp33_ASAP7_75t_L g2036 ( .A1(n_1415), .A2(n_1419), .B1(n_2037), .B2(n_2038), .Y(n_2036) );
AND2x4_ASAP7_75t_L g1425 ( .A(n_1416), .B(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
AOI222xp33_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1422), .B1(n_1423), .B2(n_1424), .C1(n_1428), .C2(n_1429), .Y(n_1420) );
BUFx4f_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
BUFx2_ASAP7_75t_L g2035 ( .A(n_1430), .Y(n_2035) );
INVx5_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
AOI31xp33_ASAP7_75t_L g1433 ( .A1(n_1434), .A2(n_1445), .A3(n_1453), .B(n_1458), .Y(n_1433) );
AOI211xp5_ASAP7_75t_L g1434 ( .A1(n_1435), .A2(n_1436), .B(n_1438), .C(n_1441), .Y(n_1434) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
AOI22xp33_ASAP7_75t_SL g1445 ( .A1(n_1446), .A2(n_1448), .B1(n_1449), .B2(n_1452), .Y(n_1445) );
AND2x4_ASAP7_75t_L g1449 ( .A(n_1447), .B(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g1481 ( .A(n_1451), .Y(n_1481) );
INVx4_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1468), .Y(n_1459) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
BUFx3_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1470), .Y(n_1522) );
INVx2_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
BUFx3_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1489), .Y(n_1717) );
OAI22xp5_ASAP7_75t_L g1489 ( .A1(n_1490), .A2(n_1632), .B1(n_1633), .B2(n_1714), .Y(n_1489) );
INVx2_ASAP7_75t_L g1714 ( .A(n_1490), .Y(n_1714) );
AO22x2_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1533), .B1(n_1534), .B2(n_1631), .Y(n_1490) );
INVx2_ASAP7_75t_SL g1631 ( .A(n_1491), .Y(n_1631) );
XNOR2x1_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g1774 ( .A1(n_1492), .A2(n_1775), .B1(n_1776), .B2(n_1777), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1513), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1519), .Y(n_1513) );
NAND2xp5_ASAP7_75t_SL g1519 ( .A(n_1520), .B(n_1530), .Y(n_1519) );
INVx2_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVx2_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
XOR2x2_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1586), .Y(n_1534) );
NAND4xp25_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1545), .C(n_1559), .D(n_1581), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1541), .Y(n_1537) );
INVx2_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx2_ASAP7_75t_SL g1663 ( .A(n_1553), .Y(n_1663) );
INVx2_ASAP7_75t_L g2055 ( .A(n_1553), .Y(n_2055) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx2_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
NAND3xp33_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1574), .C(n_1577), .Y(n_1572) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
NAND4xp25_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1610), .C(n_1625), .D(n_1630), .Y(n_1587) );
NAND3xp33_ASAP7_75t_SL g1599 ( .A(n_1600), .B(n_1602), .C(n_1606), .Y(n_1599) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g2053 ( .A(n_1615), .Y(n_2053) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1628), .Y(n_1625) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
OAI22xp5_ASAP7_75t_L g1633 ( .A1(n_1634), .A2(n_1673), .B1(n_1674), .B2(n_1713), .Y(n_1633) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1634), .Y(n_1713) );
NAND3xp33_ASAP7_75t_L g1635 ( .A(n_1636), .B(n_1657), .C(n_1659), .Y(n_1635) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1644), .Y(n_1636) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1638), .B(n_1641), .Y(n_1637) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
HB1xp67_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1699), .Y(n_1676) );
NOR3xp33_ASAP7_75t_SL g1677 ( .A(n_1678), .B(n_1685), .C(n_1686), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1679), .B(n_1682), .Y(n_1678) );
NAND3xp33_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1707), .C(n_1711), .Y(n_1700) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
OAI221xp5_ASAP7_75t_L g1718 ( .A1(n_1719), .A2(n_1968), .B1(n_1969), .B2(n_2020), .C(n_2026), .Y(n_1718) );
O2A1O1Ixp33_ASAP7_75t_L g1719 ( .A1(n_1720), .A2(n_1850), .B(n_1886), .C(n_1936), .Y(n_1719) );
NAND5xp2_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1807), .C(n_1835), .D(n_1844), .E(n_1848), .Y(n_1720) );
AOI221xp5_ASAP7_75t_L g1721 ( .A1(n_1722), .A2(n_1758), .B1(n_1782), .B2(n_1789), .C(n_1796), .Y(n_1721) );
INVxp67_ASAP7_75t_SL g1722 ( .A(n_1723), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1748), .Y(n_1723) );
AOI221xp5_ASAP7_75t_L g1937 ( .A1(n_1724), .A2(n_1765), .B1(n_1871), .B2(n_1938), .C(n_1939), .Y(n_1937) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1725), .B(n_1744), .Y(n_1724) );
INVx2_ASAP7_75t_L g1751 ( .A(n_1725), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1725), .B(n_1788), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1802 ( .A(n_1725), .B(n_1752), .Y(n_1802) );
OR2x2_ASAP7_75t_L g1838 ( .A(n_1725), .B(n_1752), .Y(n_1838) );
NOR2xp33_ASAP7_75t_L g1892 ( .A(n_1725), .B(n_1744), .Y(n_1892) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1738), .Y(n_1725) );
AND2x4_ASAP7_75t_L g1727 ( .A(n_1728), .B(n_1733), .Y(n_1727) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
OR2x2_ASAP7_75t_L g1755 ( .A(n_1729), .B(n_1734), .Y(n_1755) );
NAND2xp5_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1732), .Y(n_1729) );
HB1xp67_ASAP7_75t_L g2082 ( .A(n_1730), .Y(n_2082) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1732), .Y(n_1742) );
AND2x4_ASAP7_75t_L g1735 ( .A(n_1733), .B(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
OR2x2_ASAP7_75t_L g1757 ( .A(n_1734), .B(n_1737), .Y(n_1757) );
BUFx2_ASAP7_75t_L g1793 ( .A(n_1735), .Y(n_1793) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1740), .B(n_1741), .Y(n_1739) );
AND2x4_ASAP7_75t_L g1743 ( .A(n_1740), .B(n_1742), .Y(n_1743) );
AND2x4_ASAP7_75t_L g1764 ( .A(n_1740), .B(n_1741), .Y(n_1764) );
HB1xp67_ASAP7_75t_L g2083 ( .A(n_1741), .Y(n_2083) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx2_ASAP7_75t_L g1777 ( .A(n_1743), .Y(n_1777) );
OR2x2_ASAP7_75t_L g1801 ( .A(n_1744), .B(n_1761), .Y(n_1801) );
OR2x2_ASAP7_75t_L g1811 ( .A(n_1744), .B(n_1812), .Y(n_1811) );
NAND2xp5_ASAP7_75t_L g1813 ( .A(n_1744), .B(n_1751), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1826 ( .A(n_1744), .B(n_1787), .Y(n_1826) );
AND2x2_ASAP7_75t_L g1898 ( .A(n_1744), .B(n_1899), .Y(n_1898) );
OAI322xp33_ASAP7_75t_L g1908 ( .A1(n_1744), .A2(n_1894), .A3(n_1909), .B1(n_1910), .B2(n_1911), .C1(n_1912), .C2(n_1914), .Y(n_1908) );
AND2x2_ASAP7_75t_L g1913 ( .A(n_1744), .B(n_1788), .Y(n_1913) );
BUFx3_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
INVxp67_ASAP7_75t_L g1749 ( .A(n_1745), .Y(n_1749) );
BUFx2_ASAP7_75t_L g1818 ( .A(n_1745), .Y(n_1818) );
OR2x2_ASAP7_75t_L g1855 ( .A(n_1745), .B(n_1752), .Y(n_1855) );
AND2x2_ASAP7_75t_L g1864 ( .A(n_1745), .B(n_1865), .Y(n_1864) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1746), .B(n_1747), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1847 ( .A(n_1748), .B(n_1823), .Y(n_1847) );
NAND2xp5_ASAP7_75t_L g1872 ( .A(n_1748), .B(n_1761), .Y(n_1872) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1749), .B(n_1750), .Y(n_1748) );
NAND2xp5_ASAP7_75t_L g1786 ( .A(n_1749), .B(n_1787), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1836 ( .A(n_1749), .B(n_1837), .Y(n_1836) );
AND2x2_ASAP7_75t_L g1950 ( .A(n_1749), .B(n_1870), .Y(n_1950) );
AND2x2_ASAP7_75t_L g1964 ( .A(n_1749), .B(n_1865), .Y(n_1964) );
AND2x2_ASAP7_75t_L g1804 ( .A(n_1750), .B(n_1760), .Y(n_1804) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1750), .Y(n_1879) );
AND2x2_ASAP7_75t_L g1903 ( .A(n_1750), .B(n_1818), .Y(n_1903) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1751), .B(n_1752), .Y(n_1750) );
INVx2_ASAP7_75t_SL g1788 ( .A(n_1752), .Y(n_1788) );
OAI22xp5_ASAP7_75t_L g1753 ( .A1(n_1754), .A2(n_1755), .B1(n_1756), .B2(n_1757), .Y(n_1753) );
BUFx6f_ASAP7_75t_L g1769 ( .A(n_1755), .Y(n_1769) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1757), .Y(n_1772) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1765), .Y(n_1759) );
NOR2xp33_ASAP7_75t_L g1837 ( .A(n_1760), .B(n_1838), .Y(n_1837) );
AND2x2_ASAP7_75t_L g1878 ( .A(n_1760), .B(n_1865), .Y(n_1878) );
AND2x2_ASAP7_75t_L g1899 ( .A(n_1760), .B(n_1802), .Y(n_1899) );
NOR2xp33_ASAP7_75t_L g1952 ( .A(n_1760), .B(n_1825), .Y(n_1952) );
INVx2_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
BUFx2_ASAP7_75t_L g1785 ( .A(n_1761), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1817 ( .A(n_1761), .B(n_1818), .Y(n_1817) );
INVx2_ASAP7_75t_L g1824 ( .A(n_1761), .Y(n_1824) );
AND2x2_ASAP7_75t_L g1870 ( .A(n_1761), .B(n_1802), .Y(n_1870) );
NAND2xp5_ASAP7_75t_L g1909 ( .A(n_1761), .B(n_1843), .Y(n_1909) );
NAND2xp5_ASAP7_75t_L g1922 ( .A(n_1761), .B(n_1766), .Y(n_1922) );
AND2x2_ASAP7_75t_L g1931 ( .A(n_1761), .B(n_1846), .Y(n_1931) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1763), .Y(n_1761) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1764), .Y(n_1775) );
BUFx3_ASAP7_75t_L g1829 ( .A(n_1764), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1839 ( .A(n_1765), .B(n_1840), .Y(n_1839) );
INVx1_ASAP7_75t_L g1926 ( .A(n_1765), .Y(n_1926) );
AND2x4_ASAP7_75t_L g1765 ( .A(n_1766), .B(n_1778), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1766), .B(n_1779), .Y(n_1798) );
HB1xp67_ASAP7_75t_L g1815 ( .A(n_1766), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1823 ( .A(n_1766), .B(n_1824), .Y(n_1823) );
INVx2_ASAP7_75t_SL g1861 ( .A(n_1766), .Y(n_1861) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1766), .Y(n_1881) );
NAND2xp5_ASAP7_75t_L g1907 ( .A(n_1766), .B(n_1840), .Y(n_1907) );
NOR2xp33_ASAP7_75t_L g1918 ( .A(n_1766), .B(n_1824), .Y(n_1918) );
CKINVDCx5p33_ASAP7_75t_R g1766 ( .A(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1843 ( .A(n_1767), .B(n_1778), .Y(n_1843) );
AND2x2_ASAP7_75t_L g1928 ( .A(n_1767), .B(n_1779), .Y(n_1928) );
OR2x2_ASAP7_75t_L g1767 ( .A(n_1768), .B(n_1774), .Y(n_1767) );
OAI22xp5_ASAP7_75t_L g1768 ( .A1(n_1769), .A2(n_1770), .B1(n_1771), .B2(n_1773), .Y(n_1768) );
BUFx3_ASAP7_75t_L g1832 ( .A(n_1769), .Y(n_1832) );
HB1xp67_ASAP7_75t_L g1834 ( .A(n_1771), .Y(n_1834) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVx2_ASAP7_75t_L g1795 ( .A(n_1777), .Y(n_1795) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1778), .B(n_1791), .Y(n_1806) );
OR2x2_ASAP7_75t_L g1820 ( .A(n_1778), .B(n_1821), .Y(n_1820) );
AOI22xp5_ASAP7_75t_L g1852 ( .A1(n_1778), .A2(n_1853), .B1(n_1854), .B2(n_1856), .Y(n_1852) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1778), .Y(n_1867) );
NAND3xp33_ASAP7_75t_L g1917 ( .A(n_1778), .B(n_1865), .C(n_1918), .Y(n_1917) );
NOR2xp33_ASAP7_75t_L g1921 ( .A(n_1778), .B(n_1922), .Y(n_1921) );
INVx3_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1789 ( .A(n_1779), .B(n_1790), .Y(n_1789) );
OR2x2_ASAP7_75t_L g1862 ( .A(n_1779), .B(n_1791), .Y(n_1862) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1780), .B(n_1781), .Y(n_1779) );
AOI211xp5_ASAP7_75t_L g1941 ( .A1(n_1782), .A2(n_1798), .B(n_1942), .C(n_1953), .Y(n_1941) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
OR2x2_ASAP7_75t_L g1783 ( .A(n_1784), .B(n_1786), .Y(n_1783) );
NAND2xp5_ASAP7_75t_L g1809 ( .A(n_1784), .B(n_1789), .Y(n_1809) );
NAND2xp5_ASAP7_75t_L g1891 ( .A(n_1784), .B(n_1892), .Y(n_1891) );
NAND2xp5_ASAP7_75t_L g1902 ( .A(n_1784), .B(n_1903), .Y(n_1902) );
OAI21xp33_ASAP7_75t_L g1965 ( .A1(n_1784), .A2(n_1879), .B(n_1966), .Y(n_1965) );
INVx2_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
NAND2xp5_ASAP7_75t_L g1934 ( .A(n_1785), .B(n_1787), .Y(n_1934) );
NAND2xp5_ASAP7_75t_L g1946 ( .A(n_1785), .B(n_1867), .Y(n_1946) );
INVx1_ASAP7_75t_L g1925 ( .A(n_1787), .Y(n_1925) );
NOR2x1_ASAP7_75t_L g1961 ( .A(n_1788), .B(n_1818), .Y(n_1961) );
NAND2xp5_ASAP7_75t_L g1880 ( .A(n_1789), .B(n_1881), .Y(n_1880) );
AOI22xp5_ASAP7_75t_L g1897 ( .A1(n_1789), .A2(n_1847), .B1(n_1867), .B2(n_1898), .Y(n_1897) );
AOI322xp5_ASAP7_75t_L g1962 ( .A1(n_1789), .A2(n_1854), .A3(n_1889), .B1(n_1963), .B2(n_1964), .C1(n_1965), .C2(n_1967), .Y(n_1962) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1790), .Y(n_1840) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1790), .Y(n_1851) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1791), .Y(n_1821) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1791), .Y(n_1846) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_1792), .B(n_1794), .Y(n_1791) );
OAI22xp5_ASAP7_75t_L g1796 ( .A1(n_1797), .A2(n_1799), .B1(n_1803), .B2(n_1805), .Y(n_1796) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
NAND2xp5_ASAP7_75t_L g1799 ( .A(n_1800), .B(n_1802), .Y(n_1799) );
OAI211xp5_ASAP7_75t_SL g1956 ( .A1(n_1800), .A2(n_1899), .B(n_1957), .C(n_1960), .Y(n_1956) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
OR2x2_ASAP7_75t_L g1905 ( .A(n_1801), .B(n_1838), .Y(n_1905) );
OR2x2_ASAP7_75t_L g1924 ( .A(n_1801), .B(n_1925), .Y(n_1924) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1802), .Y(n_1812) );
NAND2xp5_ASAP7_75t_L g1816 ( .A(n_1802), .B(n_1817), .Y(n_1816) );
AND2x2_ASAP7_75t_L g1856 ( .A(n_1802), .B(n_1818), .Y(n_1856) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
OAI21xp33_ASAP7_75t_L g1951 ( .A1(n_1804), .A2(n_1839), .B(n_1952), .Y(n_1951) );
NAND2xp5_ASAP7_75t_L g1863 ( .A(n_1805), .B(n_1864), .Y(n_1863) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
AOI221xp5_ASAP7_75t_L g1887 ( .A1(n_1806), .A2(n_1888), .B1(n_1889), .B2(n_1890), .C(n_1893), .Y(n_1887) );
NAND2xp5_ASAP7_75t_L g1911 ( .A(n_1806), .B(n_1881), .Y(n_1911) );
AOI211xp5_ASAP7_75t_SL g1807 ( .A1(n_1808), .A2(n_1810), .B(n_1814), .C(n_1819), .Y(n_1807) );
INVxp67_ASAP7_75t_SL g1808 ( .A(n_1809), .Y(n_1808) );
NAND2xp5_ASAP7_75t_L g1810 ( .A(n_1811), .B(n_1813), .Y(n_1810) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1811), .Y(n_1888) );
NOR2xp33_ASAP7_75t_L g1841 ( .A(n_1813), .B(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1944 ( .A(n_1813), .Y(n_1944) );
NOR2xp33_ASAP7_75t_L g1814 ( .A(n_1815), .B(n_1816), .Y(n_1814) );
A2O1A1Ixp33_ASAP7_75t_L g1954 ( .A1(n_1815), .A2(n_1870), .B(n_1904), .C(n_1955), .Y(n_1954) );
NAND2xp5_ASAP7_75t_L g1868 ( .A(n_1816), .B(n_1869), .Y(n_1868) );
AND2x2_ASAP7_75t_L g1948 ( .A(n_1817), .B(n_1865), .Y(n_1948) );
AOI321xp33_ASAP7_75t_L g1929 ( .A1(n_1818), .A2(n_1930), .A3(n_1931), .B1(n_1932), .B2(n_1933), .C(n_1935), .Y(n_1929) );
A2O1A1Ixp33_ASAP7_75t_L g1819 ( .A1(n_1820), .A2(n_1822), .B(n_1825), .C(n_1827), .Y(n_1819) );
INVx1_ASAP7_75t_L g1955 ( .A(n_1820), .Y(n_1955) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
NAND2xp5_ASAP7_75t_L g1842 ( .A(n_1824), .B(n_1843), .Y(n_1842) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
INVx3_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
INVx3_ASAP7_75t_L g1935 ( .A(n_1828), .Y(n_1935) );
CKINVDCx5p33_ASAP7_75t_R g1968 ( .A(n_1829), .Y(n_1968) );
OAI22xp33_ASAP7_75t_L g1830 ( .A1(n_1831), .A2(n_1832), .B1(n_1833), .B2(n_1834), .Y(n_1830) );
AOI21xp5_ASAP7_75t_L g1835 ( .A1(n_1836), .A2(n_1839), .B(n_1841), .Y(n_1835) );
INVx1_ASAP7_75t_L g1914 ( .A(n_1837), .Y(n_1914) );
NOR2xp33_ASAP7_75t_L g1849 ( .A(n_1838), .B(n_1842), .Y(n_1849) );
INVx1_ASAP7_75t_L g1865 ( .A(n_1838), .Y(n_1865) );
AND2x2_ASAP7_75t_L g1895 ( .A(n_1840), .B(n_1881), .Y(n_1895) );
INVx2_ASAP7_75t_L g1910 ( .A(n_1840), .Y(n_1910) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1842), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1889 ( .A(n_1843), .B(n_1846), .Y(n_1889) );
NAND2xp5_ASAP7_75t_L g1844 ( .A(n_1845), .B(n_1847), .Y(n_1844) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
NAND2xp5_ASAP7_75t_L g1875 ( .A(n_1846), .B(n_1876), .Y(n_1875) );
INVxp67_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
OAI211xp5_ASAP7_75t_L g1850 ( .A1(n_1851), .A2(n_1852), .B(n_1857), .C(n_1882), .Y(n_1850) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1851), .Y(n_1873) );
OAI211xp5_ASAP7_75t_SL g1936 ( .A1(n_1851), .A2(n_1937), .B(n_1941), .C(n_1962), .Y(n_1936) );
INVx1_ASAP7_75t_L g1959 ( .A(n_1851), .Y(n_1959) );
NAND2xp5_ASAP7_75t_L g1920 ( .A(n_1854), .B(n_1921), .Y(n_1920) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
INVx1_ASAP7_75t_L g1940 ( .A(n_1856), .Y(n_1940) );
AOI221xp5_ASAP7_75t_L g1857 ( .A1(n_1858), .A2(n_1870), .B1(n_1871), .B2(n_1873), .C(n_1874), .Y(n_1857) );
NAND3xp33_ASAP7_75t_L g1858 ( .A(n_1859), .B(n_1863), .C(n_1866), .Y(n_1858) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
NOR2xp33_ASAP7_75t_L g1860 ( .A(n_1861), .B(n_1862), .Y(n_1860) );
INVx2_ASAP7_75t_L g1869 ( .A(n_1861), .Y(n_1869) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1861), .Y(n_1876) );
AND2x2_ASAP7_75t_L g1947 ( .A(n_1861), .B(n_1948), .Y(n_1947) );
INVxp67_ASAP7_75t_L g1884 ( .A(n_1863), .Y(n_1884) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1864), .Y(n_1896) );
INVxp67_ASAP7_75t_L g1883 ( .A(n_1866), .Y(n_1883) );
NAND2xp5_ASAP7_75t_L g1866 ( .A(n_1867), .B(n_1868), .Y(n_1866) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
OAI22xp5_ASAP7_75t_L g1874 ( .A1(n_1875), .A2(n_1877), .B1(n_1879), .B2(n_1880), .Y(n_1874) );
INVx1_ASAP7_75t_L g1932 ( .A(n_1875), .Y(n_1932) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1878), .Y(n_1877) );
NAND2xp5_ASAP7_75t_L g1930 ( .A(n_1879), .B(n_1925), .Y(n_1930) );
INVx1_ASAP7_75t_L g1967 ( .A(n_1880), .Y(n_1967) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1881), .Y(n_1885) );
OAI21xp5_ASAP7_75t_L g1882 ( .A1(n_1883), .A2(n_1884), .B(n_1885), .Y(n_1882) );
NAND5xp2_ASAP7_75t_L g1886 ( .A(n_1887), .B(n_1897), .C(n_1900), .D(n_1915), .E(n_1929), .Y(n_1886) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
NOR2xp33_ASAP7_75t_L g1893 ( .A(n_1894), .B(n_1896), .Y(n_1893) );
INVx1_ASAP7_75t_L g1894 ( .A(n_1895), .Y(n_1894) );
O2A1O1Ixp33_ASAP7_75t_L g1900 ( .A1(n_1901), .A2(n_1904), .B(n_1906), .C(n_1908), .Y(n_1900) );
INVx1_ASAP7_75t_L g1901 ( .A(n_1902), .Y(n_1901) );
INVx1_ASAP7_75t_L g1966 ( .A(n_1903), .Y(n_1966) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
OAI22xp33_ASAP7_75t_L g1923 ( .A1(n_1905), .A2(n_1924), .B1(n_1926), .B2(n_1927), .Y(n_1923) );
INVx1_ASAP7_75t_L g1906 ( .A(n_1907), .Y(n_1906) );
INVx1_ASAP7_75t_L g1938 ( .A(n_1909), .Y(n_1938) );
OAI221xp5_ASAP7_75t_L g1942 ( .A1(n_1910), .A2(n_1911), .B1(n_1943), .B2(n_1949), .C(n_1951), .Y(n_1942) );
INVx1_ASAP7_75t_L g1912 ( .A(n_1913), .Y(n_1912) );
NOR3xp33_ASAP7_75t_SL g1915 ( .A(n_1916), .B(n_1919), .C(n_1923), .Y(n_1915) );
INVxp67_ASAP7_75t_L g1916 ( .A(n_1917), .Y(n_1916) );
INVxp67_ASAP7_75t_SL g1919 ( .A(n_1920), .Y(n_1919) );
INVx1_ASAP7_75t_L g1963 ( .A(n_1922), .Y(n_1963) );
NOR2xp33_ASAP7_75t_L g1939 ( .A(n_1926), .B(n_1940), .Y(n_1939) );
OR2x2_ASAP7_75t_L g1958 ( .A(n_1927), .B(n_1959), .Y(n_1958) );
CKINVDCx5p33_ASAP7_75t_R g1927 ( .A(n_1928), .Y(n_1927) );
INVx1_ASAP7_75t_L g1933 ( .A(n_1934), .Y(n_1933) );
AOI21xp33_ASAP7_75t_L g1943 ( .A1(n_1944), .A2(n_1945), .B(n_1947), .Y(n_1943) );
INVx1_ASAP7_75t_L g1945 ( .A(n_1946), .Y(n_1945) );
INVx1_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
NAND2xp5_ASAP7_75t_SL g1953 ( .A(n_1954), .B(n_1956), .Y(n_1953) );
INVx1_ASAP7_75t_L g1957 ( .A(n_1958), .Y(n_1957) );
INVx1_ASAP7_75t_L g1960 ( .A(n_1961), .Y(n_1960) );
INVx1_ASAP7_75t_L g1969 ( .A(n_1970), .Y(n_1969) );
HB1xp67_ASAP7_75t_L g1970 ( .A(n_1971), .Y(n_1970) );
XNOR2x1_ASAP7_75t_L g1971 ( .A(n_1972), .B(n_1973), .Y(n_1971) );
AND2x2_ASAP7_75t_L g1973 ( .A(n_1974), .B(n_2003), .Y(n_1973) );
NOR3xp33_ASAP7_75t_SL g1974 ( .A(n_1975), .B(n_1983), .C(n_1984), .Y(n_1974) );
NAND2xp5_ASAP7_75t_L g1975 ( .A(n_1976), .B(n_1980), .Y(n_1975) );
INVx1_ASAP7_75t_L g1985 ( .A(n_1986), .Y(n_1985) );
OAI22xp5_ASAP7_75t_L g1990 ( .A1(n_1991), .A2(n_1992), .B1(n_1993), .B2(n_1994), .Y(n_1990) );
INVx1_ASAP7_75t_L g1994 ( .A(n_1995), .Y(n_1994) );
AOI31xp33_ASAP7_75t_L g2005 ( .A1(n_2006), .A2(n_2012), .A3(n_2018), .B(n_2019), .Y(n_2005) );
INVx1_ASAP7_75t_L g2014 ( .A(n_2015), .Y(n_2014) );
INVx1_ASAP7_75t_SL g2020 ( .A(n_2021), .Y(n_2020) );
INVx1_ASAP7_75t_L g2021 ( .A(n_2022), .Y(n_2021) );
INVx1_ASAP7_75t_L g2022 ( .A(n_2023), .Y(n_2022) );
INVx1_ASAP7_75t_L g2023 ( .A(n_2024), .Y(n_2023) );
INVx1_ASAP7_75t_L g2024 ( .A(n_2025), .Y(n_2024) );
BUFx2_ASAP7_75t_L g2027 ( .A(n_2028), .Y(n_2027) );
A2O1A1Ixp33_ASAP7_75t_L g2080 ( .A1(n_2029), .A2(n_2081), .B(n_2083), .C(n_2084), .Y(n_2080) );
INVxp33_ASAP7_75t_L g2030 ( .A(n_2031), .Y(n_2030) );
HB1xp67_ASAP7_75t_SL g2032 ( .A(n_2033), .Y(n_2032) );
NAND4xp25_ASAP7_75t_L g2034 ( .A(n_2035), .B(n_2036), .C(n_2039), .D(n_2043), .Y(n_2034) );
OAI21xp5_ASAP7_75t_SL g2052 ( .A1(n_2040), .A2(n_2053), .B(n_2054), .Y(n_2052) );
NAND3xp33_ASAP7_75t_L g2046 ( .A(n_2047), .B(n_2062), .C(n_2066), .Y(n_2046) );
NOR3xp33_ASAP7_75t_SL g2047 ( .A(n_2048), .B(n_2050), .C(n_2056), .Y(n_2047) );
INVx2_ASAP7_75t_L g2048 ( .A(n_2049), .Y(n_2048) );
NAND2xp5_ASAP7_75t_L g2059 ( .A(n_2060), .B(n_2061), .Y(n_2059) );
OAI22xp5_ASAP7_75t_L g2069 ( .A1(n_2070), .A2(n_2072), .B1(n_2076), .B2(n_2077), .Y(n_2069) );
INVx1_ASAP7_75t_L g2070 ( .A(n_2071), .Y(n_2070) );
HB1xp67_ASAP7_75t_L g2079 ( .A(n_2080), .Y(n_2079) );
INVx1_ASAP7_75t_L g2081 ( .A(n_2082), .Y(n_2081) );
endmodule