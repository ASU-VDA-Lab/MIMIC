module fake_jpeg_23457_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_1),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_26),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_26),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_18),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_18),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_27),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_21),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_23),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_44),
.B(n_19),
.C(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_88),
.B(n_101),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_48),
.B1(n_47),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_56),
.B1(n_25),
.B2(n_31),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_36),
.B1(n_33),
.B2(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_93),
.B1(n_98),
.B2(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_36),
.B1(n_33),
.B2(n_47),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_23),
.B1(n_28),
.B2(n_30),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_27),
.B1(n_34),
.B2(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_35),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_28),
.B1(n_30),
.B2(n_19),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_28),
.B1(n_20),
.B2(n_22),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_31),
.B1(n_25),
.B2(n_35),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_44),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_25),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_25),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_56),
.A3(n_65),
.B1(n_62),
.B2(n_74),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_149),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_131),
.Y(n_163)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_52),
.CON(n_123),
.SN(n_123)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_118),
.B(n_103),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_22),
.B(n_29),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_125),
.A2(n_106),
.B(n_31),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_150),
.B1(n_92),
.B2(n_114),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_2),
.Y(n_132)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_94),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_151),
.Y(n_170)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_130),
.B1(n_101),
.B2(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_62),
.C(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_162),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_104),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_157),
.A2(n_160),
.B(n_161),
.Y(n_214)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_105),
.B(n_107),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_164),
.A2(n_6),
.B(n_7),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_166),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_177),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_169),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_184),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_90),
.B1(n_118),
.B2(n_96),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_90),
.B1(n_96),
.B2(n_100),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_100),
.B1(n_114),
.B2(n_86),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_124),
.A2(n_84),
.B1(n_86),
.B2(n_109),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_84),
.B1(n_70),
.B2(n_64),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_119),
.B1(n_140),
.B2(n_128),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_61),
.B1(n_62),
.B2(n_35),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_179),
.A2(n_186),
.B1(n_151),
.B2(n_147),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_136),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_119),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_116),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_126),
.A2(n_61),
.B1(n_31),
.B2(n_116),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_137),
.C(n_146),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_8),
.C(n_9),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_188),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_133),
.Y(n_190)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_203),
.B(n_217),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_194),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_204),
.B1(n_182),
.B2(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_129),
.B(n_5),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_216),
.B(n_10),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_6),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_154),
.B1(n_165),
.B2(n_181),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_172),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_161),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_8),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_160),
.C(n_154),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_203),
.C(n_200),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_199),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_235),
.C(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_226),
.B(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_155),
.B1(n_160),
.B2(n_186),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_228),
.B1(n_191),
.B2(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_156),
.B1(n_162),
.B2(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_209),
.B1(n_205),
.B2(n_198),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_192),
.B(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_16),
.C(n_11),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_15),
.B(n_12),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_250),
.B1(n_221),
.B2(n_239),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_217),
.C(n_193),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_214),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_263),
.B(n_253),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_262),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_188),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_255),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_233),
.B1(n_228),
.B2(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_197),
.B1(n_201),
.B2(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_195),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_191),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_204),
.B(n_243),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_201),
.C(n_190),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_234),
.C(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_195),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_236),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_219),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_271),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_237),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_220),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_277),
.C(n_279),
.Y(n_290)
);

XOR2x1_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_231),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_254),
.B1(n_256),
.B2(n_248),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_254),
.B1(n_229),
.B2(n_252),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_280),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_234),
.C(n_221),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_244),
.B1(n_246),
.B2(n_218),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_212),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_272),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_218),
.B(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_274),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_285),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_278),
.B(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_289),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_280),
.B(n_270),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_194),
.C(n_12),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_294),
.C(n_279),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_11),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_12),
.C(n_13),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_282),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_268),
.C(n_269),
.Y(n_301)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_265),
.B1(n_14),
.B2(n_15),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_14),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_292),
.B1(n_284),
.B2(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_291),
.B1(n_294),
.B2(n_290),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_313),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_300),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_293),
.B1(n_296),
.B2(n_306),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_304),
.Y(n_317)
);

AOI31xp33_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_312),
.A3(n_307),
.B(n_302),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_307),
.C(n_320),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_315),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_323),
.C(n_319),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_299),
.Y(n_329)
);


endmodule