module real_aes_10246_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_22;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_8;
wire n_10;
OAI221xp5_ASAP7_75t_L g15 ( .A1(n_0), .A2(n_5), .B1(n_16), .B2(n_17), .C(n_22), .Y(n_15) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
AOI32xp33_ASAP7_75t_L g7 ( .A1(n_2), .A2(n_8), .A3(n_9), .B1(n_13), .B2(n_15), .Y(n_7) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
INVx2_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
BUFx2_ASAP7_75t_L g21 ( .A(n_6), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_9), .B(n_12), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_SL g16 ( .A(n_17), .Y(n_16) );
INVx5_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
BUFx8_ASAP7_75t_SL g18 ( .A(n_19), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
endmodule