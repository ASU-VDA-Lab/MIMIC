module real_jpeg_30254_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_586, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;
input n_586;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_323;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_0),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_1),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_1),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_1),
.B(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_1),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_1),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_2),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_2),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_2),
.B(n_300),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g320 ( 
.A(n_2),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_2),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

NAND2x1_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_46),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_3),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_3),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_3),
.B(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

NAND2x1_ASAP7_75t_L g373 ( 
.A(n_3),
.B(n_374),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_14),
.B1(n_19),
.B2(n_21),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_5),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_6),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_6),
.B(n_184),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_6),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_6),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_6),
.B(n_441),
.Y(n_440)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_6),
.B(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_7),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_8),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_8),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_8),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_8),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_8),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_8),
.B(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_10),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_11),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_12),
.B(n_43),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_12),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_12),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_12),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_12),
.B(n_166),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_12),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_12),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_12),
.B(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_13),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_15),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_16),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_16),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_16),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_16),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_16),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_16),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_16),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_17),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_17),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_17),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_17),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g451 ( 
.A(n_17),
.B(n_452),
.Y(n_451)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_451),
.B(n_474),
.C(n_569),
.D(n_584),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_466),
.Y(n_23)
);

NAND3xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_247),
.C(n_366),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_192),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_138),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_27),
.B(n_138),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_75),
.C(n_117),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_28),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_49),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_29),
.B(n_56),
.C(n_73),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_39),
.C(n_44),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_30),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_31),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_31),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_31),
.B(n_160),
.C(n_165),
.Y(n_241)
);

AO22x1_ASAP7_75t_SL g266 ( 
.A1(n_31),
.A2(n_35),
.B1(n_36),
.B2(n_163),
.Y(n_266)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_33),
.Y(n_212)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_33),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_34),
.B(n_387),
.C(n_447),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_34),
.A2(n_35),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_34),
.B(n_86),
.C(n_451),
.Y(n_519)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22x1_ASAP7_75t_L g386 ( 
.A1(n_35),
.A2(n_36),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_255)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_48),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B1(n_73),
.B2(n_74),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B(n_55),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_54),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_53),
.Y(n_148)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_53),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_55),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_55),
.B(n_149),
.C(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

XNOR2x1_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_58),
.B(n_68),
.C(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_62),
.Y(n_220)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_62),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_64),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_64),
.B(n_373),
.C(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_66),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_66),
.Y(n_265)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_66),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_67),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_70),
.B(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_75),
.B(n_118),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_92),
.C(n_107),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_76),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_86),
.C(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_81),
.A2(n_86),
.B1(n_449),
.B2(n_455),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_81),
.B(n_492),
.C(n_506),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_81),
.A2(n_86),
.B1(n_506),
.B2(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_91),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_92),
.A2(n_107),
.B1(n_108),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_92),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.C(n_102),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_93),
.B(n_102),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

XNOR2x2_ASAP7_75t_SL g353 ( 
.A(n_98),
.B(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_106),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_106),
.Y(n_407)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_113),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_109),
.A2(n_110),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_110),
.B(n_206),
.C(n_211),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_141),
.C(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_130),
.C(n_134),
.Y(n_172)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g430 ( 
.A(n_129),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_130),
.A2(n_164),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_130),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_130),
.A2(n_492),
.B1(n_513),
.B2(n_514),
.Y(n_512)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_137),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_137),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_168),
.Y(n_138)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_156),
.Y(n_143)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_167),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_162),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_164),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_164),
.A2(n_167),
.B1(n_222),
.B2(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_167),
.B(n_489),
.C(n_492),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_167),
.B(n_518),
.C(n_537),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_190),
.B2(n_191),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_188),
.C(n_227),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_181),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_183),
.A2(n_189),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_186),
.Y(n_385)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_192),
.A2(n_468),
.B(n_469),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_193),
.B(n_196),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_197),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_228),
.B1(n_229),
.B2(n_243),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_226),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_213),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_204),
.B(n_213),
.C(n_246),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_205),
.B(n_482),
.Y(n_525)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_206),
.B(n_481),
.C(n_484),
.Y(n_480)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_258),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_210),
.A2(n_211),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_211),
.B(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_211),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_226),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

XOR2x2_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_221),
.Y(n_214)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_218),
.Y(n_379)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_220),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_221),
.B(n_222),
.C(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_222),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_222),
.A2(n_408),
.B1(n_414),
.B2(n_537),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_222),
.B(n_408),
.C(n_506),
.Y(n_584)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_224),
.Y(n_388)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_227),
.B(n_517),
.C(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_242),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

HB1xp67_ASAP7_75t_SL g393 ( 
.A(n_231),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_232),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_241),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_238),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_239),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_240),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_241),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_242),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_243),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_269),
.B(n_365),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_267),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_249),
.B(n_267),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_250),
.B(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_256),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_266),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_257),
.B(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_261),
.A2(n_262),
.B1(n_266),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_266),
.Y(n_357)
);

AOI21x1_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_359),
.B(n_364),
.Y(n_269)
);

OAI21x1_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_347),
.B(n_358),
.Y(n_270)
);

AOI21x1_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_317),
.B(n_346),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_291),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_273),
.B(n_291),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_285),
.C(n_288),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_274),
.A2(n_275),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_288),
.B1(n_289),
.B2(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_297),
.B1(n_315),
.B2(n_316),
.Y(n_291)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_296),
.C(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_306),
.C(n_310),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_328),
.B(n_345),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_324),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_334),
.B(n_344),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_331),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_350),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_353),
.C(n_355),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_SL g364 ( 
.A(n_360),
.B(n_363),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_366),
.A2(n_467),
.B(n_470),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_418),
.B1(n_457),
.B2(n_462),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_367),
.B(n_418),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_367),
.B(n_418),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_390),
.C(n_395),
.Y(n_367)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_368),
.B(n_391),
.Y(n_465)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_377),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_378),
.C(n_380),
.Y(n_436)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_387),
.Y(n_389)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_389),
.Y(n_489)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.C(n_394),
.Y(n_391)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_395)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_396),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_415),
.C(n_420),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.C(n_400),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_402),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_408),
.B1(n_412),
.B2(n_414),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_406),
.Y(n_413)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_408),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_408),
.A2(n_414),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_412),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_412),
.Y(n_435)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_428),
.C(n_431),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_419),
.B(n_566),
.C(n_568),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_437),
.B2(n_456),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_436),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_433),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_425),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_431),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_433),
.B(n_551),
.C(n_552),
.Y(n_550)
);

INVxp33_ASAP7_75t_SL g551 ( 
.A(n_436),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_437),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_448),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_446),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_439),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_440),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_440),
.A2(n_518),
.B1(n_536),
.B2(n_538),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_522),
.C(n_523),
.Y(n_521)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_449),
.Y(n_455)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_463),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.C(n_461),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_472),
.B(n_473),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_543),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_475),
.A2(n_570),
.B(n_573),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_527),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_476),
.B(n_527),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_511),
.C(n_520),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_478),
.B(n_559),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_479),
.A2(n_493),
.B1(n_509),
.B2(n_510),
.Y(n_478)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_488),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_480),
.B(n_488),
.C(n_509),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_505),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_495),
.A2(n_501),
.B1(n_503),
.B2(n_504),
.Y(n_494)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_501),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_501),
.B(n_503),
.C(n_541),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_505),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_506),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_506),
.A2(n_515),
.B1(n_580),
.B2(n_581),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_511),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_516),
.C(n_519),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_516),
.B(n_519),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_520),
.B(n_558),
.Y(n_557)
);

MAJx2_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.C(n_526),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_521),
.B(n_548),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_526),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_539),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_528),
.B(n_540),
.C(n_542),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_535),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_530),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_532),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_532),
.B(n_533),
.C(n_535),
.Y(n_583)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_536),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_542),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_560),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_544),
.A2(n_571),
.B(n_572),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_557),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_545),
.B(n_557),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_546),
.A2(n_549),
.B1(n_550),
.B2(n_555),
.Y(n_545)
);

INVxp33_ASAP7_75t_SL g546 ( 
.A(n_547),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_556),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_553),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_550),
.A2(n_562),
.B1(n_563),
.B2(n_564),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_550),
.Y(n_562)
);

OAI33xp33_ASAP7_75t_L g571 ( 
.A1(n_550),
.A2(n_562),
.A3(n_563),
.B1(n_564),
.B2(n_565),
.B3(n_586),
.Y(n_571)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_553),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_556),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_565),
.Y(n_560)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_563),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_575),
.C(n_582),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_576),
.B(n_577),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_583),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_582),
.Y(n_578)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);


endmodule