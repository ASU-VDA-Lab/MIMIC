module fake_jpeg_19128_n_235 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_19),
.B1(n_21),
.B2(n_13),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_20),
.B1(n_24),
.B2(n_14),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_20),
.B1(n_24),
.B2(n_14),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_30),
.B1(n_29),
.B2(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_32),
.B1(n_30),
.B2(n_46),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_61),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_22),
.B1(n_14),
.B2(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_74),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_55),
.B(n_48),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_27),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_18),
.B(n_25),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_58),
.B(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_83),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_52),
.B1(n_61),
.B2(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_83),
.B1(n_80),
.B2(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_65),
.B1(n_54),
.B2(n_36),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_94),
.B1(n_71),
.B2(n_72),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_18),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_54),
.B1(n_59),
.B2(n_41),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_77),
.Y(n_117)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_76),
.C(n_81),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_87),
.C(n_27),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_108),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_81),
.B(n_82),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_117),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_119),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_107),
.B1(n_109),
.B2(n_117),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_88),
.B1(n_97),
.B2(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_63),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_125),
.B1(n_133),
.B2(n_60),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_127),
.C(n_28),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_89),
.B1(n_84),
.B2(n_73),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_40),
.C(n_42),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_69),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_91),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_119),
.B(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_18),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_89),
.B1(n_84),
.B2(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_91),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_105),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_91),
.B(n_69),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_142),
.B(n_150),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_106),
.B(n_103),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_157),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_109),
.B(n_110),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_154),
.B(n_158),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_132),
.B(n_134),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_21),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_118),
.B(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_68),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_159),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_138),
.B1(n_40),
.B2(n_42),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_64),
.B(n_0),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_15),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_138),
.B1(n_127),
.B2(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_138),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_152),
.B1(n_142),
.B2(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_138),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_40),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_157),
.C(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_186),
.C(n_169),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_141),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_179),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_154),
.A3(n_140),
.B1(n_21),
.B2(n_19),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_165),
.B(n_10),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_57),
.C(n_27),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_17),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_168),
.B1(n_163),
.B2(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_191),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_164),
.B(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_195),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_198),
.Y(n_207)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_173),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_57),
.B(n_1),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_192),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_191),
.B(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_185),
.B1(n_186),
.B2(n_57),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_204),
.B1(n_202),
.B2(n_207),
.Y(n_215)
);

OAI21x1_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_9),
.B(n_2),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_208),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_15),
.C(n_28),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_15),
.C(n_28),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_195),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_11),
.B(n_5),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_10),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_10),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_223),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_8),
.B(n_4),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_15),
.C(n_25),
.Y(n_223)
);

AOI221xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_213),
.B(n_214),
.C(n_25),
.D(n_23),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

AOI321xp33_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_225),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_11),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_230),
.A2(n_229),
.B1(n_228),
.B2(n_6),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_232),
.A2(n_231),
.B(n_0),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_32),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_15),
.B(n_23),
.Y(n_235)
);


endmodule