module fake_jpeg_15637_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_41),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_26),
.B(n_29),
.C(n_25),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_47),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_14),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_24),
.B1(n_48),
.B2(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_48),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_5),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_32),
.C(n_35),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_19),
.B1(n_17),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_53),
.B1(n_58),
.B2(n_23),
.Y(n_74)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_24),
.B1(n_17),
.B2(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_13),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_44),
.B1(n_47),
.B2(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_65),
.B(n_13),
.Y(n_69)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_68),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_53),
.B(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_9),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_63),
.B1(n_64),
.B2(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_50),
.C(n_65),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_72),
.B(n_77),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_87),
.Y(n_89)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_94),
.C(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_88),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_79),
.C(n_83),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.C(n_88),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_81),
.C(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_94),
.B1(n_92),
.B2(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_12),
.B1(n_15),
.B2(n_46),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_102),
.B(n_15),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_11),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_91),
.B(n_66),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_106),
.B(n_107),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_11),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_109),
.Y(n_111)
);


endmodule