module fake_jpeg_734_n_490 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_490);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_490;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_53),
.B(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_64),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_68),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_76),
.Y(n_102)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_86),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_95),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_27),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_30),
.B1(n_47),
.B2(n_46),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_100),
.A2(n_119),
.B1(n_129),
.B2(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_43),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_106),
.B(n_110),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_43),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_53),
.A2(n_45),
.B1(n_47),
.B2(n_46),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_19),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_132),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_55),
.A2(n_30),
.B1(n_47),
.B2(n_46),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_19),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_136),
.B(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_36),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_53),
.A2(n_42),
.B1(n_33),
.B2(n_24),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_148),
.Y(n_159)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_50),
.Y(n_145)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_59),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_65),
.A2(n_42),
.B1(n_33),
.B2(n_24),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_38),
.B1(n_44),
.B2(n_42),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_27),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_54),
.A2(n_48),
.B1(n_44),
.B2(n_38),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_44),
.B1(n_48),
.B2(n_38),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_158),
.Y(n_212)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_70),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_167),
.Y(n_218)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

NAND2x1_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_59),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_165),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_101),
.B(n_91),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_166),
.B(n_169),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_78),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_85),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_58),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_170),
.B(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_172),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_96),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_174),
.A2(n_192),
.B1(n_18),
.B2(n_35),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_117),
.B(n_52),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_175),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_102),
.B(n_88),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_191),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_48),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_182),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_146),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_89),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_107),
.B(n_115),
.Y(n_182)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_120),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_82),
.B1(n_93),
.B2(n_92),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_195),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_207),
.B(n_63),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_97),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_198),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_49),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_204),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_109),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_140),
.B(n_74),
.Y(n_202)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_205),
.Y(n_250)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_135),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_208),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_72),
.B1(n_84),
.B2(n_77),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_118),
.B(n_90),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_18),
.C(n_28),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_100),
.B(n_129),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_214),
.A2(n_222),
.B(n_3),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_153),
.B1(n_152),
.B2(n_105),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_229),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_156),
.A2(n_153),
.B1(n_152),
.B2(n_105),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_167),
.A2(n_141),
.B(n_119),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_118),
.B1(n_147),
.B2(n_134),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_224),
.A2(n_228),
.B1(n_233),
.B2(n_186),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_178),
.B1(n_192),
.B2(n_174),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_57),
.B1(n_67),
.B2(n_75),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_160),
.C(n_185),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_251),
.C(n_165),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_147),
.B1(n_134),
.B2(n_144),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_182),
.A2(n_144),
.B1(n_18),
.B2(n_34),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_239),
.A2(n_242),
.B1(n_245),
.B2(n_172),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_18),
.B1(n_35),
.B2(n_28),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_159),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_155),
.A2(n_18),
.B(n_35),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_180),
.B(n_163),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_210),
.B1(n_175),
.B2(n_168),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_259),
.A2(n_263),
.B1(n_266),
.B2(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_175),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_273),
.C(n_294),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_261),
.B(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_212),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_265),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_177),
.B1(n_181),
.B2(n_187),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_232),
.B(n_200),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_264),
.B(n_267),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_195),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_238),
.A2(n_181),
.B1(n_190),
.B2(n_196),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_269),
.A2(n_301),
.B(n_221),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_208),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_209),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_274),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_204),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_276),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_189),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_161),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_218),
.A2(n_164),
.B1(n_161),
.B2(n_203),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_184),
.B1(n_188),
.B2(n_157),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_289),
.B1(n_299),
.B2(n_244),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_223),
.B(n_179),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_281),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_193),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_245),
.A2(n_193),
.B1(n_179),
.B2(n_205),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_284),
.A2(n_285),
.B1(n_229),
.B2(n_244),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_214),
.A2(n_193),
.B1(n_179),
.B2(n_18),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_220),
.B1(n_216),
.B2(n_217),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_225),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_290),
.Y(n_310)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_225),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_221),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_300),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_226),
.A2(n_197),
.B1(n_16),
.B2(n_28),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_293),
.B1(n_242),
.B2(n_247),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_226),
.A2(n_16),
.B1(n_28),
.B2(n_4),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_2),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_2),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_267),
.C(n_294),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_252),
.B(n_3),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_298),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_225),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_239),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_246),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_3),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_247),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_308),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

XOR2x2_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_254),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_312),
.A2(n_322),
.B(n_296),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_315),
.A2(n_326),
.B1(n_333),
.B2(n_337),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_316),
.A2(n_329),
.B1(n_338),
.B2(n_334),
.Y(n_370)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_256),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_341),
.C(n_297),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_325),
.A2(n_334),
.B1(n_291),
.B2(n_285),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_282),
.A2(n_250),
.B1(n_211),
.B2(n_248),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_272),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_282),
.A2(n_250),
.B1(n_211),
.B2(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_259),
.A2(n_255),
.B1(n_213),
.B2(n_240),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_301),
.A2(n_213),
.B1(n_255),
.B2(n_221),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_338),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_269),
.A2(n_234),
.B(n_215),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_336),
.A2(n_280),
.B(n_287),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_240),
.B1(n_230),
.B2(n_237),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_264),
.B(n_249),
.Y(n_341)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_265),
.B(n_276),
.C(n_298),
.D(n_290),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_342),
.A2(n_344),
.B(n_356),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_330),
.C(n_328),
.Y(n_375)
);

NOR3xp33_ASAP7_75t_SL g348 ( 
.A(n_304),
.B(n_297),
.C(n_302),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_349),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_310),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_350),
.A2(n_355),
.B1(n_365),
.B2(n_370),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_273),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_357),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_362),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_263),
.B1(n_286),
.B2(n_284),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_300),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_317),
.B(n_295),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_358),
.B(n_327),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g359 ( 
.A1(n_320),
.A2(n_266),
.A3(n_299),
.B1(n_249),
.B2(n_230),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_361),
.B(n_366),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_246),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_322),
.A2(n_336),
.B(n_321),
.Y(n_361)
);

XNOR2x2_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_243),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_234),
.Y(n_363)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_363),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_3),
.Y(n_364)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_305),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_365)
);

OAI32xp33_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_321),
.B(n_7),
.Y(n_368)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_323),
.A2(n_7),
.B(n_9),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_369),
.A2(n_361),
.B(n_344),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_326),
.A2(n_15),
.B1(n_10),
.B2(n_11),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_372),
.A2(n_318),
.B1(n_337),
.B2(n_314),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_325),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_313),
.B1(n_333),
.B2(n_340),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_393),
.C(n_397),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_353),
.B(n_341),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_384),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_324),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_346),
.B(n_327),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_387),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_349),
.B(n_339),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_386),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_309),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_398),
.Y(n_404)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_323),
.B1(n_306),
.B2(n_340),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_392),
.A2(n_345),
.B1(n_355),
.B2(n_354),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_323),
.C(n_11),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_10),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_396),
.Y(n_423)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_11),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_14),
.C(n_357),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_399),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_408),
.B1(n_418),
.B2(n_381),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_354),
.Y(n_405)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_350),
.C(n_356),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_409),
.C(n_419),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_391),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_348),
.C(n_370),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_411),
.A2(n_392),
.B1(n_400),
.B2(n_390),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_388),
.A2(n_342),
.B(n_351),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_351),
.Y(n_414)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_383),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_415),
.B(n_416),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_358),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_378),
.A2(n_373),
.B1(n_342),
.B2(n_365),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_371),
.C(n_363),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_371),
.C(n_360),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_420),
.B(n_396),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_382),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_424),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_380),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_432),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_426),
.A2(n_434),
.B1(n_411),
.B2(n_412),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_431),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_417),
.A2(n_400),
.B1(n_394),
.B2(n_397),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_368),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_433),
.Y(n_453)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_422),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_422),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_403),
.A2(n_378),
.B1(n_387),
.B2(n_389),
.Y(n_434)
);

BUFx12_ASAP7_75t_L g435 ( 
.A(n_413),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_388),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_420),
.C(n_407),
.Y(n_447)
);

AO221x1_ASAP7_75t_L g439 ( 
.A1(n_418),
.A2(n_372),
.B1(n_398),
.B2(n_359),
.C(n_393),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_439),
.B(n_442),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_449),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_440),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_402),
.C(n_410),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_401),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_450),
.B(n_451),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_402),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_409),
.Y(n_452)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_453),
.B(n_441),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_461),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_454),
.A2(n_428),
.B(n_424),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_464),
.B(n_443),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_460),
.B(n_468),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

XOR2x2_ASAP7_75t_SL g462 ( 
.A(n_443),
.B(n_436),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_447),
.Y(n_474)
);

NOR2x1_ASAP7_75t_SL g463 ( 
.A(n_448),
.B(n_440),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_449),
.Y(n_476)
);

NOR4xp25_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_428),
.C(n_441),
.D(n_414),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_426),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_476),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_467),
.A2(n_444),
.B(n_433),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_471),
.A2(n_473),
.B(n_476),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_465),
.A2(n_413),
.B(n_431),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_458),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_456),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_475),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_457),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_478),
.A2(n_481),
.B1(n_477),
.B2(n_472),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_432),
.Y(n_484)
);

AOI21xp33_ASAP7_75t_L g485 ( 
.A1(n_482),
.A2(n_478),
.B(n_404),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_483),
.B(n_484),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_485),
.Y(n_487)
);

OAI321xp33_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_486),
.A3(n_404),
.B1(n_435),
.B2(n_364),
.C(n_484),
.Y(n_488)
);

AOI322xp5_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_435),
.A3(n_366),
.B1(n_369),
.B2(n_423),
.C1(n_410),
.C2(n_14),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_423),
.Y(n_490)
);


endmodule