module fake_jpeg_16727_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx12f_ASAP7_75t_SL g67 ( 
.A(n_43),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_84),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_51),
.C(n_44),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_60),
.C(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_53),
.B1(n_48),
.B2(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_65),
.B1(n_64),
.B2(n_62),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_49),
.B(n_47),
.C(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_85),
.B1(n_79),
.B2(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_92),
.B1(n_98),
.B2(n_97),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_78),
.B(n_7),
.Y(n_107)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_77),
.B1(n_93),
.B2(n_9),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_6),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_105),
.CI(n_18),
.CON(n_111),
.SN(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_12),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.C(n_108),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_17),
.C(n_22),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_23),
.C(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_26),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_28),
.B(n_31),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_32),
.B(n_34),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_36),
.B(n_38),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_39),
.Y(n_123)
);


endmodule