module fake_jpeg_16962_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_3),
.B(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_7),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_43),
.B1(n_49),
.B2(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_74),
.B1(n_1),
.B2(n_7),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_77),
.B1(n_39),
.B2(n_14),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_56),
.B1(n_50),
.B2(n_53),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx10_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_53),
.B1(n_58),
.B2(n_48),
.Y(n_77)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_51),
.B1(n_40),
.B2(n_41),
.Y(n_86)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_47),
.A3(n_44),
.B1(n_55),
.B2(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_94),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_93),
.C(n_16),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_9),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_47),
.C(n_10),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_26),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_95),
.B1(n_83),
.B2(n_28),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_90),
.B(n_86),
.C(n_95),
.D(n_83),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_97),
.C(n_32),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_97),
.B1(n_30),
.B2(n_31),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_27),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_118),
.Y(n_121)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_113),
.B1(n_105),
.B2(n_116),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_119),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_122),
.B(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_112),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_29),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_33),
.B(n_34),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_35),
.Y(n_133)
);


endmodule