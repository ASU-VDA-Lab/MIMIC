module fake_jpeg_20667_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx8_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_0),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_13),
.B(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_13),
.B1(n_15),
.B2(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_19),
.B(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_37),
.B1(n_24),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_18),
.B1(n_10),
.B2(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_1),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_22),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_54),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_32),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_41),
.B(n_39),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_60),
.B(n_59),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_39),
.C(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_55),
.Y(n_63)
);

AOI221xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_8),
.B1(n_16),
.B2(n_17),
.C(n_7),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_53),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_48),
.B1(n_53),
.B2(n_8),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_16),
.C(n_17),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_66),
.B(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_71),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_62),
.B(n_64),
.Y(n_71)
);

OAI31xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_69),
.A3(n_5),
.B(n_6),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_2),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_40),
.C2(n_49),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_74),
.B(n_73),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_2),
.B(n_5),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_2),
.Y(n_78)
);


endmodule