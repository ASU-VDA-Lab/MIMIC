module fake_jpeg_27632_n_87 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_87);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_11),
.A2(n_20),
.B1(n_19),
.B2(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_20),
.B1(n_11),
.B2(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_13),
.B1(n_21),
.B2(n_15),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_1),
.B(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_34),
.B1(n_21),
.B2(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_3),
.B(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

A2O1A1O1Ixp25_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_32),
.B(n_33),
.C(n_22),
.D(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_18),
.B1(n_14),
.B2(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_53),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_43),
.B1(n_45),
.B2(n_42),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_40),
.B(n_4),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_37),
.C(n_25),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_37),
.C(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_59),
.B1(n_53),
.B2(n_65),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_29),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.C(n_68),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.C(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_74),
.B1(n_29),
.B2(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_65),
.B1(n_62),
.B2(n_57),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_76),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_51),
.C(n_6),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_69),
.B(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_81),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g82 ( 
.A(n_79),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_17),
.C(n_24),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_76),
.B(n_10),
.C(n_17),
.Y(n_84)
);

AOI22x1_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_85),
.B1(n_78),
.B2(n_45),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g87 ( 
.A(n_86),
.Y(n_87)
);


endmodule