module real_aes_18386_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_656;
wire n_316;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_617;
wire n_402;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_604;
wire n_115;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_899;
wire n_365;
wire n_526;
wire n_155;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_0), .Y(n_565) );
AND2x4_ASAP7_75t_L g113 ( .A(n_1), .B(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_2), .A2(n_3), .B1(n_235), .B2(n_236), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_4), .A2(n_21), .B1(n_218), .B2(n_274), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_5), .A2(n_54), .B1(n_164), .B2(n_165), .Y(n_163) );
BUFx3_ASAP7_75t_L g632 ( .A(n_6), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_7), .A2(n_15), .B1(n_200), .B2(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_9), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_10), .A2(n_14), .B1(n_897), .B2(n_898), .Y(n_896) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_10), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_11), .B(n_188), .Y(n_601) );
BUFx2_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
OR2x2_ASAP7_75t_L g135 ( .A(n_12), .B(n_33), .Y(n_135) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_13), .Y(n_156) );
INVx1_ASAP7_75t_L g898 ( .A(n_14), .Y(n_898) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_16), .B(n_155), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_17), .B(n_178), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_18), .A2(n_87), .B1(n_155), .B2(n_274), .Y(n_551) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_19), .A2(n_50), .B(n_170), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_20), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_22), .B(n_218), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_23), .B(n_152), .Y(n_246) );
INVx4_ASAP7_75t_R g187 ( .A(n_24), .Y(n_187) );
INVx1_ASAP7_75t_L g519 ( .A(n_25), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_25), .B(n_142), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_26), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_27), .A2(n_522), .B(n_901), .Y(n_900) );
AO32x1_ASAP7_75t_L g548 ( .A1(n_28), .A2(n_212), .A3(n_213), .B1(n_549), .B2(n_552), .Y(n_548) );
AO32x2_ASAP7_75t_L g640 ( .A1(n_28), .A2(n_212), .A3(n_213), .B1(n_549), .B2(n_552), .Y(n_640) );
INVx1_ASAP7_75t_L g241 ( .A(n_29), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_30), .B(n_218), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_SL g288 ( .A1(n_31), .A2(n_151), .B(n_200), .C(n_289), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_32), .A2(n_47), .B1(n_200), .B2(n_204), .Y(n_275) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_34), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_35), .A2(n_53), .B1(n_189), .B2(n_218), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_36), .A2(n_92), .B1(n_204), .B2(n_274), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_37), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_38), .B(n_574), .Y(n_578) );
INVx1_ASAP7_75t_L g250 ( .A(n_39), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_40), .B(n_200), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_41), .A2(n_69), .B1(n_204), .B2(n_655), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_42), .Y(n_216) );
INVx2_ASAP7_75t_L g124 ( .A(n_43), .Y(n_124) );
INVx1_ASAP7_75t_L g109 ( .A(n_44), .Y(n_109) );
BUFx3_ASAP7_75t_L g532 ( .A(n_44), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_45), .A2(n_66), .B1(n_138), .B2(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_45), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_46), .B(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_48), .A2(n_86), .B1(n_200), .B2(n_204), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_49), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_51), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_52), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_55), .A2(n_79), .B1(n_158), .B2(n_574), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_56), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_57), .A2(n_83), .B1(n_155), .B2(n_274), .Y(n_628) );
INVx1_ASAP7_75t_L g170 ( .A(n_58), .Y(n_170) );
AND2x4_ASAP7_75t_L g173 ( .A(n_59), .B(n_174), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_60), .A2(n_91), .B1(n_204), .B2(n_233), .Y(n_232) );
AO22x1_ASAP7_75t_L g153 ( .A1(n_61), .A2(n_74), .B1(n_154), .B2(n_157), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_62), .B(n_274), .Y(n_600) );
INVx1_ASAP7_75t_L g174 ( .A(n_63), .Y(n_174) );
AND2x2_ASAP7_75t_L g291 ( .A(n_64), .B(n_212), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_65), .B(n_212), .Y(n_606) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_67), .A2(n_161), .B(n_164), .C(n_564), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_68), .B(n_274), .C(n_604), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_70), .B(n_164), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_71), .Y(n_284) );
AND2x2_ASAP7_75t_L g566 ( .A(n_72), .B(n_195), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_73), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_75), .B(n_218), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_76), .A2(n_98), .B1(n_155), .B2(n_158), .Y(n_590) );
INVx2_ASAP7_75t_L g152 ( .A(n_77), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_78), .B(n_219), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_80), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_81), .B(n_212), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_82), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_84), .B(n_168), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_85), .A2(n_894), .B1(n_895), .B2(n_899), .Y(n_893) );
INVx1_ASAP7_75t_L g899 ( .A(n_85), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_88), .B(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_89), .A2(n_102), .B1(n_189), .B2(n_204), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_90), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_93), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g112 ( .A(n_94), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_94), .B(n_133), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_95), .A2(n_104), .B1(n_120), .B2(n_908), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_96), .B(n_178), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_97), .A2(n_164), .B(n_182), .C(n_184), .Y(n_181) );
AND2x2_ASAP7_75t_L g194 ( .A(n_99), .B(n_195), .Y(n_194) );
NAND2xp33_ASAP7_75t_L g222 ( .A(n_100), .B(n_188), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_101), .Y(n_615) );
INVx5_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_115), .Y(n_105) );
OR2x6_ASAP7_75t_L g910 ( .A(n_106), .B(n_115), .Y(n_910) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2x1p5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g133 ( .A(n_109), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g538 ( .A(n_112), .Y(n_538) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_525), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
BUFx8_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g529 ( .A(n_124), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_124), .B(n_905), .Y(n_904) );
OAI21x1_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_136), .B(n_521), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
CKINVDCx8_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_131), .Y(n_524) );
AND2x6_ASAP7_75t_SL g131 ( .A(n_132), .B(n_134), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_134), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2x1_ASAP7_75t_L g907 ( .A(n_135), .B(n_532), .Y(n_907) );
XOR2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_140), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_519), .B(n_520), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI22x1_ASAP7_75t_L g535 ( .A1(n_142), .A2(n_536), .B1(n_539), .B2(n_889), .Y(n_535) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_418), .Y(n_142) );
AND3x1_ASAP7_75t_L g143 ( .A(n_144), .B(n_336), .C(n_395), .Y(n_143) );
AOI221xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_227), .B1(n_255), .B2(n_308), .C(n_311), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_208), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_175), .Y(n_147) );
INVx2_ASAP7_75t_L g266 ( .A(n_148), .Y(n_266) );
AND2x2_ASAP7_75t_L g323 ( .A(n_148), .B(n_265), .Y(n_323) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g416 ( .A(n_149), .B(n_351), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_149), .B(n_197), .Y(n_480) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B(n_159), .C(n_171), .Y(n_150) );
INVx6_ASAP7_75t_L g202 ( .A(n_151), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_222), .B(n_223), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_151), .B(n_153), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_151), .A2(n_287), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_151), .A2(n_600), .B(n_601), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_151), .A2(n_202), .B1(n_628), .B2(n_629), .Y(n_627) );
BUFx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx1_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx1_ASAP7_75t_L g249 ( .A(n_152), .Y(n_249) );
INVxp67_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g580 ( .A(n_155), .Y(n_580) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g158 ( .A(n_156), .Y(n_158) );
INVx1_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
INVx1_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
INVx3_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_156), .Y(n_218) );
INVx1_ASAP7_75t_L g237 ( .A(n_156), .Y(n_237) );
INVx2_ASAP7_75t_L g274 ( .A(n_156), .Y(n_274) );
OAI21xp33_ASAP7_75t_SL g245 ( .A1(n_157), .A2(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_158), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g304 ( .A(n_159), .Y(n_304) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_163), .B(n_167), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_160), .A2(n_252), .B(n_253), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_160), .A2(n_202), .B1(n_273), .B2(n_275), .Y(n_272) );
AOI21x1_ASAP7_75t_L g572 ( .A1(n_160), .A2(n_573), .B(n_575), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_160), .A2(n_202), .B1(n_654), .B2(n_656), .Y(n_653) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_166), .B(n_183), .Y(n_182) );
OAI21xp33_ASAP7_75t_L g171 ( .A1(n_167), .A2(n_168), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g179 ( .A(n_168), .Y(n_179) );
INVx2_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
INVx2_ASAP7_75t_L g205 ( .A(n_168), .Y(n_205) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
INVx1_ASAP7_75t_L g306 ( .A(n_171), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_172), .A2(n_282), .B(n_288), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_172), .A2(n_558), .B(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx10_ASAP7_75t_L g193 ( .A(n_173), .Y(n_193) );
BUFx10_ASAP7_75t_L g226 ( .A(n_173), .Y(n_226) );
INVx1_ASAP7_75t_L g239 ( .A(n_173), .Y(n_239) );
AO31x2_ASAP7_75t_L g652 ( .A1(n_173), .A2(n_586), .A3(n_653), .B(n_657), .Y(n_652) );
INVx2_ASAP7_75t_L g355 ( .A(n_175), .Y(n_355) );
OR2x2_ASAP7_75t_L g444 ( .A(n_175), .B(n_361), .Y(n_444) );
OR2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_197), .Y(n_175) );
INVx1_ASAP7_75t_L g259 ( .A(n_176), .Y(n_259) );
INVx2_ASAP7_75t_L g346 ( .A(n_176), .Y(n_346) );
AND2x2_ASAP7_75t_L g370 ( .A(n_176), .B(n_197), .Y(n_370) );
AND2x4_ASAP7_75t_L g383 ( .A(n_176), .B(n_303), .Y(n_383) );
AND2x2_ASAP7_75t_L g400 ( .A(n_176), .B(n_262), .Y(n_400) );
AND2x2_ASAP7_75t_L g410 ( .A(n_176), .B(n_302), .Y(n_410) );
AND2x2_ASAP7_75t_L g438 ( .A(n_176), .B(n_210), .Y(n_438) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B(n_194), .Y(n_176) );
AOI21x1_ASAP7_75t_L g556 ( .A1(n_177), .A2(n_557), .B(n_566), .Y(n_556) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_185), .B(n_192), .Y(n_180) );
INVx1_ASAP7_75t_L g191 ( .A(n_184), .Y(n_191) );
INVx1_ASAP7_75t_L g562 ( .A(n_184), .Y(n_562) );
INVx1_ASAP7_75t_SL g589 ( .A(n_184), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_186), .B(n_191), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_186) );
INVx2_ASAP7_75t_L g233 ( .A(n_188), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_189), .A2(n_218), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g619 ( .A(n_189), .Y(n_619) );
OAI22x1_ASAP7_75t_L g198 ( .A1(n_191), .A2(n_199), .B1(n_202), .B2(n_203), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_191), .A2(n_202), .B1(n_232), .B2(n_234), .Y(n_231) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_193), .A2(n_198), .A3(n_205), .B(n_206), .Y(n_197) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_196), .B(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_196), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_196), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_196), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
AND2x2_ASAP7_75t_L g307 ( .A(n_197), .B(n_210), .Y(n_307) );
INVx2_ASAP7_75t_L g351 ( .A(n_197), .Y(n_351) );
AND2x2_ASAP7_75t_L g483 ( .A(n_197), .B(n_346), .Y(n_483) );
INVx4_ASAP7_75t_L g201 ( .A(n_200), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_201), .A2(n_216), .B(n_217), .C(n_219), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_202), .A2(n_578), .B(n_579), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_202), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_587) );
INVx2_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_204), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g576 ( .A(n_204), .Y(n_576) );
INVx2_ASAP7_75t_L g597 ( .A(n_205), .Y(n_597) );
AND3x1_ASAP7_75t_L g319 ( .A(n_208), .B(n_259), .C(n_320), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_208), .B(n_323), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_208), .B(n_483), .Y(n_500) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx2_ASAP7_75t_L g404 ( .A(n_209), .Y(n_404) );
AND2x2_ASAP7_75t_L g513 ( .A(n_209), .B(n_295), .Y(n_513) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
AND2x2_ASAP7_75t_L g264 ( .A(n_210), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g352 ( .A(n_210), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
NOR2x1_ASAP7_75t_L g224 ( .A(n_212), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
INVx4_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g254 ( .A(n_213), .B(n_226), .Y(n_254) );
INVx2_ASAP7_75t_SL g570 ( .A(n_213), .Y(n_570) );
BUFx3_ASAP7_75t_L g586 ( .A(n_213), .Y(n_586) );
INVx2_ASAP7_75t_L g612 ( .A(n_213), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_213), .B(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_213), .B(n_658), .Y(n_657) );
OAI21x1_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_221), .B(n_224), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_218), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g655 ( .A(n_218), .Y(n_655) );
INVx2_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_220), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AO31x2_ASAP7_75t_L g271 ( .A1(n_226), .A2(n_272), .A3(n_276), .B(n_277), .Y(n_271) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_226), .A2(n_599), .B(n_602), .Y(n_598) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_226), .A2(n_614), .B(n_617), .Y(n_613) );
AOI31xp67_ASAP7_75t_L g626 ( .A1(n_226), .A2(n_276), .A3(n_627), .B(n_630), .Y(n_626) );
BUFx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g379 ( .A(n_228), .B(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g486 ( .A(n_228), .B(n_376), .Y(n_486) );
AND2x2_ASAP7_75t_L g493 ( .A(n_228), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_242), .Y(n_228) );
INVx1_ASAP7_75t_L g310 ( .A(n_229), .Y(n_310) );
INVx1_ASAP7_75t_L g328 ( .A(n_229), .Y(n_328) );
OR2x2_ASAP7_75t_L g332 ( .A(n_229), .B(n_271), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_229), .B(n_271), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_229), .B(n_297), .Y(n_358) );
INVx1_ASAP7_75t_L g430 ( .A(n_229), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_229), .B(n_279), .Y(n_489) );
AO31x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .A3(n_238), .B(n_240), .Y(n_229) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_230), .A2(n_281), .B(n_291), .Y(n_280) );
O2A1O1Ixp5_ASAP7_75t_L g614 ( .A1(n_236), .A2(n_287), .B(n_615), .C(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_237), .B(n_286), .Y(n_285) );
AO31x2_ASAP7_75t_L g585 ( .A1(n_238), .A2(n_586), .A3(n_587), .B(n_591), .Y(n_585) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_SL g552 ( .A(n_239), .Y(n_552) );
OR2x2_ASAP7_75t_L g327 ( .A(n_242), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_242), .B(n_295), .Y(n_334) );
INVx3_ASAP7_75t_L g342 ( .A(n_242), .Y(n_342) );
NAND2x1p5_ASAP7_75t_SL g367 ( .A(n_242), .B(n_341), .Y(n_367) );
BUFx2_ASAP7_75t_L g389 ( .A(n_242), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_242), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_242), .B(n_430), .Y(n_447) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_251), .B(n_254), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
BUFx4f_ASAP7_75t_L g287 ( .A(n_249), .Y(n_287) );
INVx1_ASAP7_75t_L g604 ( .A(n_249), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_292), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_263), .B(n_267), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g325 ( .A(n_259), .Y(n_325) );
INVx1_ASAP7_75t_L g417 ( .A(n_259), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_260), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g453 ( .A(n_260), .B(n_370), .Y(n_453) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g465 ( .A(n_261), .B(n_383), .Y(n_465) );
BUFx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g369 ( .A(n_262), .B(n_302), .Y(n_369) );
AND2x2_ASAP7_75t_L g409 ( .A(n_262), .B(n_351), .Y(n_409) );
AND2x4_ASAP7_75t_SL g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_264), .B(n_345), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_264), .B(n_383), .Y(n_392) );
AND2x2_ASAP7_75t_L g432 ( .A(n_264), .B(n_425), .Y(n_432) );
INVx1_ASAP7_75t_L g449 ( .A(n_265), .Y(n_449) );
OAI322xp33_ASAP7_75t_L g311 ( .A1(n_266), .A2(n_312), .A3(n_318), .B1(n_321), .B2(n_326), .C1(n_330), .C2(n_335), .Y(n_311) );
AOI32xp33_ASAP7_75t_L g402 ( .A1(n_266), .A2(n_362), .A3(n_403), .B1(n_405), .B2(n_407), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_266), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g490 ( .A(n_266), .B(n_409), .Y(n_490) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g329 ( .A(n_270), .Y(n_329) );
AND2x2_ASAP7_75t_L g393 ( .A(n_270), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g467 ( .A(n_270), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_270), .B(n_429), .Y(n_468) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_279), .Y(n_270) );
INVx2_ASAP7_75t_SL g297 ( .A(n_271), .Y(n_297) );
BUFx2_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_274), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_SL g574 ( .A(n_274), .Y(n_574) );
INVx2_ASAP7_75t_L g341 ( .A(n_279), .Y(n_341) );
OR2x2_ASAP7_75t_L g377 ( .A(n_279), .B(n_297), .Y(n_377) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g295 ( .A(n_280), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B(n_287), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_298), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g494 ( .A(n_294), .Y(n_494) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_295), .B(n_342), .Y(n_357) );
INVxp67_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
OR2x2_ASAP7_75t_L g434 ( .A(n_296), .B(n_341), .Y(n_434) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_307), .Y(n_299) );
AND2x2_ASAP7_75t_L g354 ( .A(n_300), .B(n_355), .Y(n_354) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_300), .B(n_352), .Y(n_517) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g425 ( .A(n_301), .Y(n_425) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g345 ( .A(n_302), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g450 ( .A(n_303), .B(n_346), .Y(n_450) );
AOI21x1_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_306), .Y(n_303) );
INVx2_ASAP7_75t_L g386 ( .A(n_307), .Y(n_386) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g317 ( .A(n_310), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g390 ( .A(n_313), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_313), .B(n_429), .Y(n_498) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_314), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g457 ( .A(n_314), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g366 ( .A(n_317), .B(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_317), .B(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
INVx1_ASAP7_75t_L g458 ( .A(n_327), .Y(n_458) );
INVx1_ASAP7_75t_L g508 ( .A(n_327), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_331), .B(n_381), .Y(n_413) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
OR2x2_ASAP7_75t_L g406 ( .A(n_332), .B(n_367), .Y(n_406) );
OR2x2_ASAP7_75t_L g474 ( .A(n_332), .B(n_381), .Y(n_474) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g422 ( .A(n_334), .B(n_339), .Y(n_422) );
INVx1_ASAP7_75t_L g505 ( .A(n_335), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_371), .Y(n_336) );
OAI321xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .A3(n_347), .B1(n_353), .B2(n_356), .C(n_359), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_338), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
AND2x4_ASAP7_75t_L g429 ( .A(n_342), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g433 ( .A(n_342), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_344), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_348), .A2(n_440), .B(n_443), .C(n_445), .Y(n_439) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g437 ( .A(n_350), .Y(n_437) );
INVx1_ASAP7_75t_L g471 ( .A(n_350), .Y(n_471) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g361 ( .A(n_352), .Y(n_361) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_355), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_356), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_357), .Y(n_461) );
AOI32xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .A3(n_363), .B1(n_365), .B2(n_368), .Y(n_359) );
OR2x2_ASAP7_75t_L g515 ( .A(n_361), .B(n_416), .Y(n_515) );
AND2x2_ASAP7_75t_L g396 ( .A(n_363), .B(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g441 ( .A(n_364), .B(n_442), .Y(n_441) );
NAND2x1_ASAP7_75t_L g507 ( .A(n_364), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AND2x2_ASAP7_75t_L g487 ( .A(n_369), .B(n_483), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_370), .B(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_370), .A2(n_397), .B1(n_493), .B2(n_495), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_378), .B2(n_382), .C(n_384), .Y(n_371) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g428 ( .A(n_376), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g518 ( .A(n_380), .B(n_397), .Y(n_518) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g388 ( .A(n_383), .Y(n_388) );
AND2x2_ASAP7_75t_L g495 ( .A(n_383), .B(n_437), .Y(n_495) );
AOI32xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .A3(n_390), .B1(n_391), .B2(n_393), .Y(n_384) );
NOR2xp33_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g397 ( .A(n_394), .B(n_398), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B(n_401), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_397), .A2(n_412), .B(n_414), .Y(n_411) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_397), .A2(n_511), .B(n_514), .Y(n_510) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_411), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g509 ( .A(n_410), .B(n_471), .Y(n_509) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NOR4xp75_ASAP7_75t_L g418 ( .A(n_419), .B(n_451), .C(n_475), .D(n_501), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_439), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_426), .Y(n_420) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_424), .A2(n_464), .B1(n_466), .B2(n_468), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_431), .B1(n_433), .B2(n_435), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_427), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g442 ( .A(n_429), .Y(n_442) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_436), .A2(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g469 ( .A1(n_444), .A2(n_470), .B(n_472), .Y(n_469) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
OR2x2_ASAP7_75t_L g466 ( .A(n_447), .B(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g462 ( .A(n_448), .Y(n_462) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B(n_459), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_462), .B(n_463), .C(n_469), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g484 ( .A(n_466), .Y(n_484) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2x1_ASAP7_75t_SL g475 ( .A(n_476), .B(n_491), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_481), .B(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_488), .B2(n_490), .Y(n_485) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_493), .A2(n_505), .B1(n_506), .B2(n_509), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_516), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVxp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2xp67_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
OAI21xp5_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_533), .B(n_900), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
BUFx12f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x6_ASAP7_75t_SL g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_892), .B2(n_893), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx12f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
BUFx8_ASAP7_75t_SL g891 ( .A(n_538), .Y(n_891) );
AND2x2_ASAP7_75t_L g906 ( .A(n_538), .B(n_907), .Y(n_906) );
NOR2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_809), .Y(n_539) );
NAND4xp75_ASAP7_75t_L g540 ( .A(n_541), .B(n_688), .C(n_741), .D(n_786), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_645), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_582), .B(n_607), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
AND2x4_ASAP7_75t_L g777 ( .A(n_545), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_545), .B(n_651), .Y(n_805) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_546), .B(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g770 ( .A(n_547), .Y(n_770) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_547), .Y(n_792) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g676 ( .A(n_548), .B(n_652), .Y(n_676) );
INVx1_ASAP7_75t_L g698 ( .A(n_548), .Y(n_698) );
AND2x2_ASAP7_75t_L g732 ( .A(n_548), .B(n_652), .Y(n_732) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_552), .A2(n_572), .B(n_577), .Y(n_571) );
INVxp33_ASAP7_75t_L g727 ( .A(n_553), .Y(n_727) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g839 ( .A(n_554), .B(n_676), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_567), .Y(n_554) );
OR2x2_ASAP7_75t_L g719 ( .A(n_555), .B(n_568), .Y(n_719) );
INVx1_ASAP7_75t_L g752 ( .A(n_555), .Y(n_752) );
INVx1_ASAP7_75t_L g756 ( .A(n_555), .Y(n_756) );
AND2x2_ASAP7_75t_L g872 ( .A(n_555), .B(n_687), .Y(n_872) );
OR2x2_ASAP7_75t_L g878 ( .A(n_555), .B(n_698), .Y(n_878) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g637 ( .A(n_556), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_559), .B(n_562), .Y(n_558) );
AND2x2_ASAP7_75t_L g772 ( .A(n_567), .B(n_722), .Y(n_772) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g638 ( .A(n_568), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g642 ( .A(n_568), .B(n_639), .Y(n_642) );
AND2x2_ASAP7_75t_L g649 ( .A(n_568), .B(n_640), .Y(n_649) );
INVx2_ASAP7_75t_L g673 ( .A(n_568), .Y(n_673) );
INVx1_ASAP7_75t_L g696 ( .A(n_568), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_568), .B(n_652), .Y(n_769) );
AND2x2_ASAP7_75t_L g778 ( .A(n_568), .B(n_636), .Y(n_778) );
INVxp67_ASAP7_75t_L g848 ( .A(n_568), .Y(n_848) );
BUFx2_ASAP7_75t_L g856 ( .A(n_568), .Y(n_856) );
INVx1_ASAP7_75t_L g886 ( .A(n_568), .Y(n_886) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B(n_581), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_576), .A2(n_603), .B(n_605), .Y(n_602) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_593), .Y(n_583) );
OR2x2_ASAP7_75t_L g644 ( .A(n_584), .B(n_610), .Y(n_644) );
AND2x2_ASAP7_75t_L g794 ( .A(n_584), .B(n_678), .Y(n_794) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g623 ( .A(n_585), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g670 ( .A(n_585), .Y(n_670) );
AND2x2_ASAP7_75t_L g693 ( .A(n_585), .B(n_664), .Y(n_693) );
INVx1_ASAP7_75t_L g726 ( .A(n_585), .Y(n_726) );
AND2x2_ASAP7_75t_L g762 ( .A(n_585), .B(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g767 ( .A(n_585), .B(n_624), .Y(n_767) );
AND2x2_ASAP7_75t_L g825 ( .A(n_585), .B(n_667), .Y(n_825) );
OR2x2_ASAP7_75t_L g834 ( .A(n_585), .B(n_611), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_593), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g710 ( .A(n_594), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_594), .B(n_663), .Y(n_751) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g680 ( .A(n_595), .Y(n_680) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g704 ( .A(n_596), .B(n_625), .Y(n_704) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_606), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_597), .A2(n_598), .B(n_606), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_633), .B1(n_641), .B2(n_643), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_609), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_623), .Y(n_609) );
INVx1_ASAP7_75t_L g775 ( .A(n_610), .Y(n_775) );
OR2x2_ASAP7_75t_L g888 ( .A(n_610), .B(n_784), .Y(n_888) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_622), .Y(n_610) );
INVx2_ASAP7_75t_SL g660 ( .A(n_611), .Y(n_660) );
BUFx2_ASAP7_75t_L g701 ( .A(n_611), .Y(n_701) );
AND2x2_ASAP7_75t_L g725 ( .A(n_611), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g763 ( .A(n_611), .Y(n_763) );
OA21x2_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_621), .Y(n_611) );
OA21x2_ASAP7_75t_L g667 ( .A1(n_612), .A2(n_613), .B(n_621), .Y(n_667) );
AND2x2_ASAP7_75t_L g666 ( .A(n_622), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g826 ( .A(n_622), .B(n_664), .Y(n_826) );
INVx1_ASAP7_75t_L g683 ( .A(n_623), .Y(n_683) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g664 ( .A(n_626), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
AND2x2_ASAP7_75t_L g882 ( .A(n_635), .B(n_649), .Y(n_882) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g651 ( .A(n_637), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g686 ( .A(n_637), .Y(n_686) );
INVx1_ASAP7_75t_L g699 ( .A(n_637), .Y(n_699) );
INVx1_ASAP7_75t_L g791 ( .A(n_637), .Y(n_791) );
NAND2x1p5_ASAP7_75t_L g684 ( .A(n_638), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g690 ( .A(n_638), .B(n_651), .Y(n_690) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g722 ( .A(n_640), .B(n_687), .Y(n_722) );
INVx1_ASAP7_75t_L g740 ( .A(n_640), .Y(n_740) );
INVx2_ASAP7_75t_L g835 ( .A(n_641), .Y(n_835) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI321xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_659), .A3(n_661), .B1(n_665), .B2(n_671), .C(n_674), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g671 ( .A(n_651), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g712 ( .A(n_651), .B(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g687 ( .A(n_652), .Y(n_687) );
AND2x2_ASAP7_75t_L g790 ( .A(n_652), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_660), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_662), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g735 ( .A(n_663), .Y(n_735) );
AND2x2_ASAP7_75t_L g797 ( .A(n_663), .B(n_726), .Y(n_797) );
AND2x2_ASAP7_75t_L g817 ( .A(n_663), .B(n_680), .Y(n_817) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g711 ( .A(n_664), .B(n_667), .Y(n_711) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
AND2x2_ASAP7_75t_L g796 ( .A(n_666), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_SL g836 ( .A(n_666), .Y(n_836) );
INVx1_ASAP7_75t_L g681 ( .A(n_667), .Y(n_681) );
OAI32xp33_ASAP7_75t_L g674 ( .A1(n_668), .A2(n_675), .A3(n_677), .B1(n_682), .B2(n_684), .Y(n_674) );
OR2x2_ASAP7_75t_L g708 ( .A(n_668), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g702 ( .A(n_669), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_669), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g869 ( .A(n_669), .B(n_704), .Y(n_869) );
INVx2_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g716 ( .A(n_670), .B(n_680), .Y(n_716) );
OR2x2_ASAP7_75t_L g885 ( .A(n_670), .B(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_672), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g675 ( .A(n_673), .B(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_673), .Y(n_713) );
OR2x2_ASAP7_75t_L g730 ( .A(n_673), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g863 ( .A(n_673), .B(n_790), .Y(n_863) );
INVxp67_ASAP7_75t_SL g877 ( .A(n_673), .Y(n_877) );
INVx2_ASAP7_75t_L g814 ( .A(n_676), .Y(n_814) );
OR2x2_ASAP7_75t_L g855 ( .A(n_676), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g859 ( .A(n_677), .Y(n_859) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g873 ( .A(n_678), .B(n_693), .Y(n_873) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g734 ( .A(n_679), .B(n_735), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx2_ASAP7_75t_L g830 ( .A(n_685), .Y(n_830) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g746 ( .A(n_687), .Y(n_746) );
INVx1_ASAP7_75t_L g782 ( .A(n_687), .Y(n_782) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_705), .Y(n_688) );
AO22x1_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_694), .B2(n_700), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g784 ( .A(n_693), .Y(n_784) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_695), .A2(n_788), .B1(n_793), .B2(n_795), .Y(n_787) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g738 ( .A(n_699), .Y(n_738) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g766 ( .A(n_701), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g803 ( .A(n_701), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_702), .A2(n_808), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g724 ( .A(n_704), .Y(n_724) );
OR2x2_ASAP7_75t_L g849 ( .A(n_704), .B(n_834), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_706), .B(n_728), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_712), .B(n_714), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_707), .A2(n_729), .B1(n_733), .B2(n_736), .Y(n_728) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g759 ( .A(n_709), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx2_ASAP7_75t_L g785 ( .A(n_710), .Y(n_785) );
AND2x2_ASAP7_75t_L g842 ( .A(n_710), .B(n_725), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_711), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g744 ( .A(n_713), .B(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_723), .B2(n_727), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_719), .B(n_731), .Y(n_841) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp33_ASAP7_75t_R g736 ( .A(n_721), .B(n_737), .Y(n_736) );
INVx3_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g754 ( .A(n_722), .B(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g808 ( .A(n_722), .B(n_752), .Y(n_808) );
BUFx2_ASAP7_75t_L g871 ( .A(n_722), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g802 ( .A(n_724), .B(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g846 ( .A(n_724), .B(n_762), .Y(n_846) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_731), .Y(n_801) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g819 ( .A(n_732), .B(n_756), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g867 ( .A(n_738), .Y(n_867) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g862 ( .A(n_740), .Y(n_862) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_764), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_747), .B(n_753), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_743), .A2(n_844), .B(n_852), .Y(n_843) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_752), .Y(n_750) );
AND2x2_ASAP7_75t_L g813 ( .A(n_752), .B(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g816 ( .A(n_762), .B(n_817), .Y(n_816) );
OAI211xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_768), .B(n_771), .C(n_776), .Y(n_764) );
INVxp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI21xp5_ASAP7_75t_SL g852 ( .A1(n_768), .A2(n_849), .B(n_853), .Y(n_852) );
OR2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B(n_783), .C(n_785), .Y(n_776) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_778), .Y(n_851) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g880 ( .A(n_785), .Y(n_880) );
NOR3x1_ASAP7_75t_L g786 ( .A(n_787), .B(n_798), .C(n_806), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_796), .A2(n_800), .B1(n_802), .B2(n_804), .Y(n_799) );
INVx2_ASAP7_75t_L g881 ( .A(n_797), .Y(n_881) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_802), .B(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_802), .A2(n_876), .B1(n_879), .B2(n_882), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_802), .A2(n_819), .B1(n_884), .B2(n_887), .Y(n_883) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND4xp75_ASAP7_75t_L g809 ( .A(n_810), .B(n_843), .C(n_857), .D(n_874), .Y(n_809) );
NOR2xp67_ASAP7_75t_L g810 ( .A(n_811), .B(n_827), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_815), .B1(n_818), .B2(n_820), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g822 ( .A(n_816), .Y(n_822) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AND2x2_ASAP7_75t_L g832 ( .A(n_826), .B(n_833), .Y(n_832) );
OAI321xp33_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_831), .A3(n_835), .B1(n_836), .B2(n_837), .C(n_840), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_830), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_832), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_847), .B1(n_849), .B2(n_850), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_848), .Y(n_847) );
INVxp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_855), .Y(n_868) );
NOR2x1_ASAP7_75t_L g857 ( .A(n_858), .B(n_864), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_863), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_868), .B(n_869), .C(n_870), .Y(n_864) );
INVxp33_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
OAI21xp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B(n_873), .Y(n_870) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_883), .Y(n_874) );
NOR2x1p5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
NOR2xp67_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
INVx3_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx10_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx3_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
INVx4_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
endmodule