module fake_jpeg_30352_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_11),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx9p33_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_66),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_61),
.B1(n_57),
.B2(n_49),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_61),
.B1(n_57),
.B2(n_71),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_53),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_69),
.Y(n_103)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_50),
.B1(n_53),
.B2(n_69),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_104),
.B1(n_111),
.B2(n_5),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_84),
.B1(n_97),
.B2(n_87),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_91),
.B1(n_87),
.B2(n_84),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_62),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_54),
.C(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_115),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_50),
.B1(n_53),
.B2(n_69),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_72),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_73),
.B1(n_50),
.B2(n_67),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_124),
.B(n_23),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_73),
.B1(n_68),
.B2(n_60),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_25),
.B(n_48),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_132),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_13),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_7),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_4),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_26),
.A3(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_6),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_24),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_28),
.CI(n_43),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_151),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_20),
.C(n_40),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_154),
.B1(n_133),
.B2(n_137),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_32),
.C(n_38),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_143),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_132),
.B1(n_138),
.B2(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_155),
.B1(n_153),
.B2(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_15),
.B(n_16),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_167),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_146),
.B(n_145),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_144),
.B1(n_164),
.B2(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_166),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_170),
.B(n_169),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_165),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_159),
.B(n_141),
.C(n_160),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_150),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_17),
.Y(n_177)
);


endmodule