module fake_jpeg_2241_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_38),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_61),
.Y(n_64)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_43),
.B1(n_51),
.B2(n_47),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_47),
.B1(n_48),
.B2(n_39),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_68),
.B1(n_40),
.B2(n_54),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_53),
.B1(n_54),
.B2(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_58),
.B1(n_60),
.B2(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_67),
.B1(n_58),
.B2(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_40),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_102),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_74),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_62),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_51),
.B1(n_62),
.B2(n_48),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_51),
.B1(n_46),
.B2(n_2),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_46),
.B1(n_1),
.B2(n_3),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_0),
.B(n_3),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_110),
.C(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_33),
.C(n_29),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_100),
.B(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_4),
.B(n_5),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_14),
.C(n_15),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_6),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_8),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_118),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_25),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_20),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_97),
.B1(n_101),
.B2(n_92),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_122),
.B1(n_126),
.B2(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_132),
.B1(n_115),
.B2(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_12),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_107),
.B(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_137),
.C(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_105),
.B1(n_114),
.B2(n_112),
.Y(n_137)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_141),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_124),
.C(n_129),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_121),
.C(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_121),
.C(n_140),
.Y(n_145)
);

NAND4xp25_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_142),
.C(n_143),
.D(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_21),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_139),
.C(n_131),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_24),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_22),
.B(n_23),
.Y(n_151)
);


endmodule