module fake_netlist_6_3111_n_1882 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_581, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_393, n_411, n_503, n_152, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1882);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1882;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_699;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_608;
wire n_630;
wire n_792;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_776;
wire n_1823;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_652;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_861;
wire n_857;
wire n_967;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_1260;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1805;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1868;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_176),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_560),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_521),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_517),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_390),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_576),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_459),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_228),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_22),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_206),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_140),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_562),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_289),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_439),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_410),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_351),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_78),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_380),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_220),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_234),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_569),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_66),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_409),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_547),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_166),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_357),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_201),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_233),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_415),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_579),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_342),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_435),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_334),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_114),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_40),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_568),
.Y(n_637)
);

BUFx5_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_102),
.Y(n_639)
);

CKINVDCx14_ASAP7_75t_R g640 ( 
.A(n_252),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_462),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_429),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_571),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_596),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_68),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_495),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_501),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_432),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_419),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_88),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_561),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_111),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_423),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_430),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_331),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_199),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_534),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_103),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_232),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_156),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_154),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_589),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_281),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_590),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_134),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_585),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_163),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_359),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_183),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_408),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

INVx4_ASAP7_75t_R g673 ( 
.A(n_190),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_105),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_145),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_555),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_420),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_424),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_142),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_592),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_32),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_416),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_600),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_15),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_241),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_240),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_481),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_519),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_386),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_177),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_178),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_76),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_51),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_411),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_136),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_54),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_155),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_591),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_421),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_597),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_598),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_180),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

CKINVDCx14_ASAP7_75t_R g705 ( 
.A(n_426),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_230),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_427),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_531),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_532),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_13),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_587),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_273),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_440),
.Y(n_713)
);

CKINVDCx16_ASAP7_75t_R g714 ( 
.A(n_394),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_394),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_515),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_321),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_94),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_109),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_574),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_276),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_187),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_412),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_413),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_397),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_586),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_60),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_40),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_428),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_418),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_233),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_8),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_21),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_565),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_566),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_491),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_463),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_582),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_324),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_205),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_138),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_580),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_142),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_487),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_422),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_488),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_578),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_417),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_131),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_575),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_458),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_493),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_492),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_557),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_490),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_572),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_244),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_476),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_320),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_60),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_121),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_431),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_594),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_553),
.Y(n_764)
);

CKINVDCx14_ASAP7_75t_R g765 ( 
.A(n_356),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_414),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_135),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_464),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_477),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_272),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_513),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_82),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_255),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_244),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_195),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_379),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_282),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_211),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_494),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_550),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_583),
.Y(n_781)
);

HB1xp67_ASAP7_75t_SL g782 ( 
.A(n_588),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_570),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_510),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_101),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_559),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_133),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_226),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_287),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_449),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_162),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_581),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_573),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_516),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_450),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_31),
.Y(n_796)
);

CKINVDCx14_ASAP7_75t_R g797 ( 
.A(n_599),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_115),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_238),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_444),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_99),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_73),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_399),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_287),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_486),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_520),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_593),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_584),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_563),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_558),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_425),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_136),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_95),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_508),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_256),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_344),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_381),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_14),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_489),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_112),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_234),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_556),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_729),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_604),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_651),
.B(n_1),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_725),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_603),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_725),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_601),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_740),
.Y(n_831)
);

CKINVDCx14_ASAP7_75t_R g832 ( 
.A(n_640),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_740),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_740),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_607),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_740),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_608),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_817),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_705),
.B(n_0),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_601),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_753),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_614),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_615),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_726),
.B(n_752),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_642),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_642),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_631),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_642),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_735),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_660),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_703),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_660),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_765),
.B(n_2),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_805),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_809),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_661),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_667),
.B(n_3),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_637),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_613),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_661),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_643),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_661),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_666),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_647),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_714),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_773),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_845),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_856),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_830),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_840),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_844),
.B(n_662),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_842),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_846),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_848),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_850),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_863),
.B(n_793),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_852),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_860),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_862),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_866),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_838),
.B(n_797),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_827),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_839),
.B(n_622),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_824),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_829),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_831),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_833),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_865),
.B(n_701),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_834),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_836),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_825),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_857),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_853),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_835),
.B(n_837),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_832),
.B(n_733),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_843),
.B(n_711),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_SL g898 ( 
.A1(n_859),
.A2(n_632),
.B1(n_658),
.B2(n_623),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_847),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_858),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_828),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_861),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_864),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_851),
.Y(n_904)
);

AND2x6_ASAP7_75t_L g905 ( 
.A(n_826),
.B(n_622),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_823),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_891),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_876),
.B(n_639),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_884),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_885),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_904),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_886),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_896),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_887),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_902),
.Y(n_915)
);

BUFx10_ASAP7_75t_L g916 ( 
.A(n_906),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_890),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_873),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_873),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_875),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_901),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_905),
.B(n_625),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_905),
.B(n_883),
.Y(n_923)
);

INVx4_ASAP7_75t_SL g924 ( 
.A(n_898),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_899),
.B(n_841),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_903),
.Y(n_926)
);

INVx4_ASAP7_75t_SL g927 ( 
.A(n_895),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_892),
.B(n_646),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_869),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_882),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_900),
.B(n_696),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_889),
.Y(n_932)
);

AO22x2_ASAP7_75t_L g933 ( 
.A1(n_888),
.A2(n_707),
.B1(n_728),
.B2(n_706),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_897),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_870),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_893),
.B(n_720),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_872),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_881),
.B(n_720),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_877),
.A2(n_619),
.B1(n_782),
.B2(n_606),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_878),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_874),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_880),
.B(n_854),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_879),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_867),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_868),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_904),
.B(n_730),
.Y(n_946)
);

BUFx4f_ASAP7_75t_L g947 ( 
.A(n_894),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_871),
.B(n_855),
.Y(n_948)
);

OAI221xp5_ASAP7_75t_L g949 ( 
.A1(n_928),
.A2(n_770),
.B1(n_616),
.B2(n_617),
.C(n_609),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_909),
.B(n_910),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_935),
.Y(n_951)
);

AO22x2_ASAP7_75t_L g952 ( 
.A1(n_924),
.A2(n_785),
.B1(n_762),
.B2(n_620),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_921),
.Y(n_953)
);

BUFx8_ASAP7_75t_L g954 ( 
.A(n_911),
.Y(n_954)
);

AO22x2_ASAP7_75t_L g955 ( 
.A1(n_946),
.A2(n_621),
.B1(n_629),
.B2(n_624),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_907),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_940),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_912),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_914),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_917),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_944),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_945),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_941),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_915),
.B(n_602),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_926),
.B(n_605),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_939),
.A2(n_645),
.B1(n_659),
.B2(n_636),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_913),
.B(n_724),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_943),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_937),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_932),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_929),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_922),
.B(n_657),
.Y(n_972)
);

AO22x2_ASAP7_75t_L g973 ( 
.A1(n_936),
.A2(n_679),
.B1(n_684),
.B2(n_671),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_933),
.A2(n_699),
.B1(n_704),
.B2(n_687),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_919),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_934),
.B(n_633),
.Y(n_976)
);

AO22x2_ASAP7_75t_L g977 ( 
.A1(n_938),
.A2(n_669),
.B1(n_674),
.B2(n_665),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_920),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_923),
.B(n_641),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_942),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_908),
.B(n_918),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_931),
.B(n_644),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_948),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_916),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_927),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_925),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_946),
.B(n_741),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_947),
.Y(n_988)
);

AO22x2_ASAP7_75t_L g989 ( 
.A1(n_924),
.A2(n_732),
.B1(n_766),
.B2(n_718),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_935),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_911),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_911),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_935),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_911),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_935),
.Y(n_995)
);

AO22x2_ASAP7_75t_L g996 ( 
.A1(n_924),
.A2(n_682),
.B1(n_685),
.B2(n_675),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_909),
.B(n_672),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_915),
.B(n_676),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_915),
.B(n_689),
.Y(n_999)
);

AO22x2_ASAP7_75t_L g1000 ( 
.A1(n_924),
.A2(n_695),
.B1(n_700),
.B2(n_686),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_930),
.Y(n_1001)
);

BUFx8_ASAP7_75t_L g1002 ( 
.A(n_911),
.Y(n_1002)
);

OR2x2_ASAP7_75t_SL g1003 ( 
.A(n_946),
.B(n_610),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_935),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_935),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_908),
.B(n_804),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_930),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_935),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_935),
.Y(n_1009)
);

AO22x2_ASAP7_75t_L g1010 ( 
.A1(n_924),
.A2(n_760),
.B1(n_767),
.B2(n_757),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_935),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_935),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_969),
.B(n_664),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_951),
.B(n_713),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_991),
.B(n_680),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_992),
.B(n_683),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_957),
.B(n_734),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_983),
.B(n_688),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_958),
.B(n_736),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_950),
.B(n_702),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_SL g1021 ( 
.A(n_985),
.B(n_731),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_959),
.B(n_708),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_960),
.B(n_709),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_990),
.B(n_716),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_993),
.B(n_995),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_SL g1026 ( 
.A(n_956),
.B(n_745),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_970),
.B(n_772),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_984),
.B(n_802),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_987),
.B(n_813),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1004),
.B(n_747),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1005),
.B(n_737),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_1008),
.B(n_750),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1009),
.B(n_738),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1011),
.B(n_776),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_1012),
.B(n_751),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_961),
.B(n_755),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_962),
.B(n_756),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_979),
.B(n_763),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_SL g1039 ( 
.A(n_967),
.B(n_764),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_953),
.B(n_768),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_981),
.B(n_778),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_968),
.B(n_779),
.Y(n_1042)
);

NAND2xp33_ASAP7_75t_SL g1043 ( 
.A(n_974),
.B(n_780),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_971),
.B(n_781),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_SL g1045 ( 
.A(n_982),
.B(n_784),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_963),
.B(n_786),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1001),
.B(n_744),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1007),
.B(n_792),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_997),
.B(n_795),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_972),
.B(n_810),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_977),
.B(n_746),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_976),
.B(n_1006),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_975),
.B(n_814),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_978),
.B(n_611),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_965),
.B(n_758),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_964),
.B(n_783),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_998),
.B(n_742),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1003),
.B(n_612),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_999),
.B(n_807),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_954),
.B(n_807),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_994),
.B(n_807),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1002),
.B(n_819),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_973),
.B(n_754),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_955),
.B(n_769),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_955),
.B(n_771),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_966),
.B(n_790),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_989),
.B(n_794),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_952),
.B(n_618),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_996),
.B(n_800),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_996),
.B(n_806),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1000),
.B(n_808),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1010),
.B(n_822),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_949),
.B(n_638),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_986),
.B(n_638),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_986),
.B(n_638),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_988),
.B(n_626),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_969),
.B(n_627),
.Y(n_1077)
);

NAND2xp33_ASAP7_75t_SL g1078 ( 
.A(n_988),
.B(n_628),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_986),
.B(n_630),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_SL g1080 ( 
.A(n_988),
.B(n_634),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_986),
.B(n_635),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_986),
.B(n_648),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_986),
.B(n_649),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_986),
.B(n_650),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_970),
.B(n_787),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_986),
.B(n_652),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_969),
.B(n_653),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_986),
.B(n_654),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_986),
.B(n_655),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_969),
.B(n_656),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_980),
.B(n_668),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_SL g1092 ( 
.A(n_988),
.B(n_670),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_986),
.B(n_677),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_986),
.B(n_678),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_986),
.B(n_681),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_970),
.B(n_791),
.Y(n_1096)
);

NAND2xp33_ASAP7_75t_SL g1097 ( 
.A(n_988),
.B(n_690),
.Y(n_1097)
);

CKINVDCx8_ASAP7_75t_R g1098 ( 
.A(n_1041),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1091),
.B(n_691),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1074),
.A2(n_803),
.B(n_796),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1095),
.B(n_692),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1075),
.A2(n_694),
.B(n_663),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_1051),
.A2(n_717),
.A3(n_739),
.B(n_719),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1027),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_1025),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_SL g1106 ( 
.A1(n_1063),
.A2(n_798),
.B(n_434),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_SL g1107 ( 
.A(n_1013),
.B(n_433),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1047),
.A2(n_697),
.B(n_693),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1052),
.B(n_436),
.Y(n_1109)
);

AOI221x1_ASAP7_75t_L g1110 ( 
.A1(n_1043),
.A2(n_673),
.B1(n_4),
.B2(n_2),
.C(n_3),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1077),
.B(n_698),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1014),
.A2(n_438),
.B(n_437),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1029),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1020),
.A2(n_442),
.B(n_441),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1027),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1022),
.A2(n_445),
.B(n_443),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1023),
.A2(n_447),
.B(n_446),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1017),
.A2(n_1031),
.B(n_1019),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1087),
.A2(n_712),
.B1(n_715),
.B2(n_710),
.Y(n_1119)
);

OA21x2_ASAP7_75t_L g1120 ( 
.A1(n_1033),
.A2(n_722),
.B(n_721),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1041),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1018),
.B(n_723),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1046),
.A2(n_451),
.B(n_448),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1090),
.B(n_727),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1085),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1085),
.B(n_452),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1058),
.B(n_1068),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1026),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1048),
.A2(n_454),
.B(n_453),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1024),
.A2(n_456),
.B(n_455),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_1096),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_1034),
.Y(n_1132)
);

NOR2x1_ASAP7_75t_SL g1133 ( 
.A(n_1044),
.B(n_457),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1067),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1069),
.B(n_5),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1079),
.A2(n_748),
.B1(n_749),
.B2(n_743),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1066),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1042),
.A2(n_461),
.B(n_460),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1081),
.A2(n_761),
.B(n_759),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1028),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1082),
.B(n_774),
.Y(n_1141)
);

AO32x2_ASAP7_75t_L g1142 ( 
.A1(n_1064),
.A2(n_9),
.A3(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1083),
.B(n_1084),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1065),
.Y(n_1144)
);

INVx3_ASAP7_75t_R g1145 ( 
.A(n_1060),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1030),
.A2(n_1035),
.B(n_1032),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1061),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1036),
.A2(n_466),
.B(n_465),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1070),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1040),
.B(n_775),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1037),
.A2(n_468),
.B(n_467),
.Y(n_1151)
);

AO22x2_ASAP7_75t_L g1152 ( 
.A1(n_1071),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1086),
.B(n_777),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1062),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_L g1155 ( 
.A1(n_1050),
.A2(n_470),
.B(n_471),
.C(n_469),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1054),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1038),
.A2(n_473),
.B(n_472),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1049),
.A2(n_475),
.B(n_474),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1088),
.B(n_788),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1089),
.B(n_789),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1072),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1055),
.B(n_11),
.Y(n_1162)
);

AOI221x1_ASAP7_75t_L g1163 ( 
.A1(n_1045),
.A2(n_1039),
.B1(n_1053),
.B2(n_1021),
.C(n_1076),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1073),
.A2(n_479),
.A3(n_480),
.B(n_478),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_1131),
.B(n_1056),
.Y(n_1165)
);

OA21x2_ASAP7_75t_L g1166 ( 
.A1(n_1118),
.A2(n_1094),
.B(n_1093),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1125),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1113),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1123),
.A2(n_1129),
.B(n_1158),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1137),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1101),
.B(n_1015),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1100),
.A2(n_1059),
.B(n_1057),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1111),
.B(n_1016),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1128),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1138),
.A2(n_1080),
.B(n_1078),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1144),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1135),
.B(n_1092),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1098),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1105),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1110),
.A2(n_1097),
.A3(n_482),
.B(n_483),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1124),
.B(n_799),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_1149),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1143),
.A2(n_485),
.B(n_484),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1122),
.B(n_801),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1146),
.A2(n_812),
.B(n_811),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1112),
.A2(n_497),
.B(n_496),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1155),
.A2(n_1114),
.B(n_1157),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1107),
.A2(n_499),
.A3(n_500),
.B(n_498),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1163),
.A2(n_503),
.A3(n_504),
.B(n_502),
.Y(n_1190)
);

AOI222xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1136),
.A2(n_820),
.B1(n_816),
.B2(n_821),
.C1(n_818),
.C2(n_815),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1133),
.A2(n_506),
.A3(n_507),
.B(n_505),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1104),
.B(n_509),
.Y(n_1193)
);

INVx3_ASAP7_75t_SL g1194 ( 
.A(n_1154),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1115),
.B(n_12),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1161),
.Y(n_1196)
);

INVx5_ASAP7_75t_L g1197 ( 
.A(n_1121),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1103),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1121),
.B(n_511),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1103),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1119),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.C(n_19),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1134),
.B(n_512),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1150),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1160),
.B(n_20),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1140),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_1116),
.A2(n_1130),
.B(n_1117),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1156),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1126),
.B(n_514),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1135),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1120),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1109),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1108),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1139),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1141),
.B(n_23),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1142),
.Y(n_1215)
);

OR3x4_ASAP7_75t_SL g1216 ( 
.A(n_1145),
.B(n_1152),
.C(n_1162),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1152),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1153),
.B(n_26),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1159),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1164),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1148),
.A2(n_522),
.B(n_518),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1151),
.A2(n_525),
.B(n_524),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1125),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1102),
.A2(n_527),
.B(n_526),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1128),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1099),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1226)
);

OAI222xp33_ASAP7_75t_L g1227 ( 
.A1(n_1135),
.A2(n_30),
.B1(n_32),
.B2(n_28),
.C1(n_29),
.C2(n_31),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1147),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1102),
.A2(n_529),
.B(n_528),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1102),
.A2(n_533),
.B(n_530),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1106),
.A2(n_536),
.B(n_535),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1099),
.B(n_33),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1170),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1177),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1197),
.B(n_537),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1196),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1180),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1198),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1200),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1183),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1167),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1217),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1173),
.B(n_34),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1195),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1207),
.Y(n_1245)
);

OR2x6_ASAP7_75t_L g1246 ( 
.A(n_1205),
.B(n_1179),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1193),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1168),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1211),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1223),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1212),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1225),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1169),
.A2(n_539),
.B(n_538),
.Y(n_1253)
);

OAI211xp5_ASAP7_75t_L g1254 ( 
.A1(n_1232),
.A2(n_1226),
.B(n_1201),
.C(n_1213),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1224),
.A2(n_541),
.B(n_540),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1215),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1228),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1203),
.B(n_542),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1228),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1204),
.B(n_35),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1182),
.B(n_36),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1197),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1194),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1166),
.Y(n_1264)
);

OAI221xp5_ASAP7_75t_L g1265 ( 
.A1(n_1185),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1220),
.A2(n_544),
.B(n_543),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1175),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1229),
.A2(n_546),
.B(n_545),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1230),
.A2(n_549),
.B(n_548),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1214),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1202),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1218),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1210),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1181),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1181),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1165),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1208),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1190),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1178),
.B(n_1209),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1219),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1190),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1171),
.B(n_38),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1174),
.B(n_39),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1178),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1252),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_R g1286 ( 
.A(n_1277),
.B(n_1186),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_R g1287 ( 
.A(n_1248),
.B(n_1221),
.Y(n_1287)
);

OR2x6_ASAP7_75t_L g1288 ( 
.A(n_1246),
.B(n_1199),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1280),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1242),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1284),
.B(n_1231),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_R g1292 ( 
.A(n_1245),
.B(n_1222),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_R g1293 ( 
.A(n_1259),
.B(n_1235),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1261),
.B(n_1216),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_R g1295 ( 
.A(n_1263),
.B(n_551),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1233),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_R g1297 ( 
.A(n_1279),
.B(n_1172),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1276),
.B(n_1176),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1234),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1250),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1271),
.B(n_552),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1282),
.B(n_1189),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1257),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1241),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1262),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1246),
.B(n_1267),
.Y(n_1306)
);

XOR2x2_ASAP7_75t_SL g1307 ( 
.A(n_1283),
.B(n_1227),
.Y(n_1307)
);

BUFx2_ASAP7_75t_SL g1308 ( 
.A(n_1247),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1270),
.B(n_1184),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_R g1310 ( 
.A(n_1272),
.B(n_1244),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1260),
.B(n_1189),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_1258),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1311),
.B(n_1251),
.Y(n_1313)
);

AOI222xp33_ASAP7_75t_L g1314 ( 
.A1(n_1294),
.A2(n_1254),
.B1(n_1265),
.B2(n_1191),
.C1(n_1243),
.C2(n_1240),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1290),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1304),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1302),
.B(n_1273),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1300),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1298),
.B(n_1238),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1289),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1296),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1299),
.B(n_1256),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1310),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1298),
.B(n_1237),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1291),
.B(n_1236),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1291),
.B(n_1249),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1309),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1306),
.Y(n_1328)
);

AND2x2_ASAP7_75t_SL g1329 ( 
.A(n_1293),
.B(n_1266),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1308),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1297),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1303),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1305),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1312),
.B(n_1278),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1287),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1285),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1307),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1286),
.A2(n_1275),
.A3(n_1274),
.B(n_1281),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1288),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1295),
.B(n_1239),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1301),
.B(n_1264),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1292),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1315),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1328),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1321),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1339),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1313),
.B(n_1253),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1322),
.Y(n_1348)
);

INVxp67_ASAP7_75t_SL g1349 ( 
.A(n_1327),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1314),
.B(n_1206),
.C(n_1192),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1332),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1323),
.B(n_1255),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1319),
.B(n_1187),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1324),
.Y(n_1354)
);

NAND2xp67_ASAP7_75t_L g1355 ( 
.A(n_1334),
.B(n_41),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1335),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1320),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1342),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1331),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1317),
.B(n_1268),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1341),
.A2(n_1269),
.B(n_1188),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1325),
.Y(n_1362)
);

NAND4xp25_ASAP7_75t_L g1363 ( 
.A(n_1333),
.B(n_43),
.C(n_41),
.D(n_42),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1326),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1330),
.Y(n_1365)
);

INVx3_ASAP7_75t_SL g1366 ( 
.A(n_1336),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1338),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1338),
.Y(n_1368)
);

OAI33xp33_ASAP7_75t_L g1369 ( 
.A1(n_1340),
.A2(n_46),
.A3(n_48),
.B1(n_44),
.B2(n_45),
.B3(n_47),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1318),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1315),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1316),
.Y(n_1372)
);

INVx5_ASAP7_75t_SL g1373 ( 
.A(n_1329),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1316),
.B(n_49),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1315),
.Y(n_1375)
);

AOI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1337),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.C(n_53),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1316),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1315),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1316),
.B(n_54),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1318),
.B(n_55),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1327),
.B(n_55),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1319),
.B(n_56),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1318),
.B(n_57),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1315),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1358),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1356),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1343),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1359),
.B(n_58),
.Y(n_1388)
);

INVxp67_ASAP7_75t_SL g1389 ( 
.A(n_1349),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1371),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1372),
.B(n_59),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1375),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1377),
.B(n_61),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1378),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1354),
.B(n_62),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1370),
.B(n_63),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1384),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1365),
.B(n_1362),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1364),
.B(n_64),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1348),
.B(n_65),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1345),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1373),
.B(n_67),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1366),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_67),
.Y(n_1404)
);

INVx3_ASAP7_75t_SL g1405 ( 
.A(n_1382),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1351),
.B(n_1347),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1352),
.B(n_69),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1368),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1367),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1360),
.B(n_70),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1374),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1379),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1357),
.B(n_71),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1361),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1381),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1353),
.B(n_72),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1353),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1380),
.B(n_74),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1355),
.B(n_74),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1383),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_1350),
.B(n_75),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1363),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1376),
.B(n_76),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1369),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1343),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1344),
.B(n_77),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1343),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1358),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1365),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1346),
.B(n_78),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1343),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1343),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1366),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1343),
.Y(n_1434)
);

OR2x2_ASAP7_75t_SL g1435 ( 
.A(n_1356),
.B(n_79),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1365),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1343),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1343),
.Y(n_1438)
);

NOR2x1_ASAP7_75t_L g1439 ( 
.A(n_1403),
.B(n_80),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1406),
.B(n_81),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1387),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1386),
.B(n_81),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1433),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1428),
.B(n_83),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1417),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1408),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1389),
.B(n_1415),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1424),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1419),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_87),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1422),
.B(n_1430),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1412),
.B(n_1390),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1392),
.B(n_88),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_SL g1454 ( 
.A(n_1405),
.B(n_1402),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1394),
.B(n_89),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1423),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_SL g1457 ( 
.A(n_1404),
.B(n_91),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1426),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1407),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1397),
.B(n_1425),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_L g1461 ( 
.A(n_1391),
.B(n_92),
.Y(n_1461)
);

AO221x2_ASAP7_75t_L g1462 ( 
.A1(n_1420),
.A2(n_96),
.B1(n_98),
.B2(n_95),
.C(n_97),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1388),
.B(n_93),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1416),
.B(n_100),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1427),
.B(n_101),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1396),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1429),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_SL g1469 ( 
.A(n_1393),
.B(n_104),
.Y(n_1469)
);

AO221x2_ASAP7_75t_L g1470 ( 
.A1(n_1400),
.A2(n_106),
.B1(n_108),
.B2(n_105),
.C(n_107),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1410),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1398),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_R g1473 ( 
.A(n_1413),
.B(n_113),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1434),
.B(n_116),
.Y(n_1474)
);

AO221x2_ASAP7_75t_L g1475 ( 
.A1(n_1399),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1437),
.B(n_122),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1438),
.B(n_123),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1395),
.Y(n_1478)
);

INVxp33_ASAP7_75t_SL g1479 ( 
.A(n_1418),
.Y(n_1479)
);

AO221x2_ASAP7_75t_L g1480 ( 
.A1(n_1436),
.A2(n_125),
.B1(n_127),
.B2(n_124),
.C(n_126),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1401),
.B(n_125),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1414),
.A2(n_1409),
.B1(n_129),
.B2(n_128),
.Y(n_1482)
);

NOR2x1_ASAP7_75t_L g1483 ( 
.A(n_1403),
.B(n_129),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1385),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1403),
.B(n_130),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1421),
.A2(n_135),
.B1(n_132),
.B2(n_133),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1386),
.B(n_137),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1385),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1403),
.B(n_139),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1424),
.A2(n_148),
.B(n_151),
.C(n_141),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1406),
.B(n_143),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1403),
.B(n_143),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1403),
.B(n_144),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1405),
.B(n_146),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1385),
.B(n_147),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1386),
.B(n_149),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1386),
.B(n_150),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1385),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1385),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1386),
.B(n_152),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1403),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1403),
.B(n_153),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1441),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1449),
.B(n_157),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1488),
.B(n_157),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1446),
.A2(n_158),
.B(n_159),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1447),
.B(n_158),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1501),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1460),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1498),
.B(n_159),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1472),
.B(n_160),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1445),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1454),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1468),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1484),
.A2(n_161),
.B(n_163),
.Y(n_1515)
);

NAND2xp33_ASAP7_75t_L g1516 ( 
.A(n_1490),
.B(n_164),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1499),
.B(n_164),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1459),
.B(n_165),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1452),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1467),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1451),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1495),
.B(n_167),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1453),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1442),
.B(n_1450),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1440),
.B(n_167),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_168),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1458),
.B(n_1466),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1455),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1443),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1464),
.B(n_169),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1448),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.C(n_173),
.Y(n_1532)
);

NOR2x1_ASAP7_75t_L g1533 ( 
.A(n_1439),
.B(n_1483),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1473),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1465),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1485),
.B(n_171),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1461),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1487),
.B(n_174),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1494),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1474),
.B(n_175),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1457),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1456),
.B(n_179),
.C(n_181),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1477),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1444),
.B(n_182),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1478),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1469),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1482),
.B(n_184),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1479),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1470),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1500),
.B(n_188),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1463),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1475),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1493),
.B(n_189),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1502),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1462),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1480),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1471),
.B(n_191),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1486),
.B(n_192),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1441),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1441),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1488),
.B(n_192),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1501),
.B(n_193),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1441),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1488),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1449),
.B(n_194),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1501),
.B(n_196),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1488),
.B(n_196),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1490),
.A2(n_197),
.B(n_198),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1488),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1488),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1488),
.B(n_199),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1447),
.B(n_200),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1488),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1495),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1458),
.Y(n_1578)
);

INVx3_ASAP7_75t_SL g1579 ( 
.A(n_1443),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1454),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1454),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1488),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1447),
.B(n_202),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1488),
.B(n_203),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1488),
.B(n_204),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1449),
.A2(n_204),
.B(n_207),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1501),
.B(n_207),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1449),
.B(n_208),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1488),
.B(n_209),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1488),
.B(n_210),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1488),
.B(n_210),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1488),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1488),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1488),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1443),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1443),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1488),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1488),
.B(n_212),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1441),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1441),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1488),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1441),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1516),
.A2(n_213),
.B(n_214),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1550),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1513),
.B(n_215),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1503),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1562),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1563),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1537),
.B(n_216),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1521),
.B(n_217),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1533),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1567),
.B(n_217),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1571),
.A2(n_218),
.B(n_219),
.Y(n_1614)
);

NAND4xp75_ASAP7_75t_SL g1615 ( 
.A(n_1515),
.B(n_223),
.C(n_221),
.D(n_222),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1555),
.A2(n_227),
.B1(n_224),
.B2(n_225),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1572),
.B(n_229),
.Y(n_1617)
);

AND2x2_ASAP7_75t_SL g1618 ( 
.A(n_1580),
.B(n_230),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_231),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1528),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1578),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1541),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1599),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1600),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1602),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1534),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1573),
.B(n_235),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1552),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1577),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1576),
.B(n_236),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1508),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1582),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1520),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1592),
.B(n_239),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1593),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1509),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1601),
.A2(n_1558),
.B1(n_1539),
.B2(n_1532),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1514),
.Y(n_1640)
);

AOI222xp33_ASAP7_75t_L g1641 ( 
.A1(n_1542),
.A2(n_245),
.B1(n_247),
.B2(n_242),
.C1(n_243),
.C2(n_246),
.Y(n_1641)
);

OAI31xp33_ASAP7_75t_L g1642 ( 
.A1(n_1554),
.A2(n_246),
.A3(n_242),
.B(n_243),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1546),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1519),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1559),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1522),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1524),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1577),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1529),
.Y(n_1649)
);

AND2x2_ASAP7_75t_SL g1650 ( 
.A(n_1548),
.B(n_1549),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1579),
.B(n_251),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1535),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1551),
.B(n_253),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1530),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1586),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1543),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1507),
.B(n_254),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1575),
.B(n_257),
.Y(n_1658)
);

AO21x1_ASAP7_75t_L g1659 ( 
.A1(n_1536),
.A2(n_257),
.B(n_258),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1544),
.B(n_258),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1512),
.B(n_259),
.Y(n_1661)
);

O2A1O1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1547),
.A2(n_262),
.B(n_260),
.C(n_261),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1561),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1583),
.B(n_266),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1556),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.C(n_269),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1568),
.B(n_270),
.C(n_271),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1518),
.B(n_272),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1531),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1525),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1557),
.B(n_274),
.Y(n_1670)
);

NAND2x1_ASAP7_75t_L g1671 ( 
.A(n_1505),
.B(n_275),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1510),
.B(n_277),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1560),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1595),
.B(n_280),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1596),
.B(n_283),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1504),
.A2(n_284),
.B(n_285),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1511),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1564),
.B(n_286),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1604),
.B(n_1570),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1612),
.B(n_1623),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1620),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1606),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1668),
.B(n_1574),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1630),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1618),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1622),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1643),
.B(n_1565),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1607),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1627),
.B(n_1584),
.Y(n_1689)
);

XNOR2xp5_ASAP7_75t_L g1690 ( 
.A(n_1650),
.B(n_1523),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1636),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1588),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1608),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1609),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1648),
.B(n_1589),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1639),
.B(n_1591),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1677),
.B(n_1598),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1631),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1633),
.B(n_1538),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1624),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1671),
.Y(n_1704)
);

OAI22xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1655),
.A2(n_1545),
.B1(n_1553),
.B2(n_1540),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1625),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1626),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1637),
.B(n_1517),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1526),
.Y(n_1709)
);

AOI31xp33_ASAP7_75t_L g1710 ( 
.A1(n_1603),
.A2(n_1587),
.A3(n_1569),
.B(n_1527),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1631),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1613),
.B(n_1506),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1628),
.B(n_288),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1634),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1653),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1676),
.B(n_290),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1672),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1659),
.B(n_291),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1646),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1675),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1647),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1649),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1611),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1614),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1641),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1652),
.B(n_296),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1656),
.B(n_296),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1661),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1638),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1635),
.B(n_297),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1642),
.B(n_297),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1617),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1660),
.B(n_298),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1640),
.B(n_298),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1644),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1711),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1692),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1720),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1681),
.Y(n_1739)
);

CKINVDCx14_ASAP7_75t_R g1740 ( 
.A(n_1690),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1680),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1734),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1701),
.Y(n_1744)
);

BUFx4f_ASAP7_75t_SL g1745 ( 
.A(n_1730),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1723),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1714),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1682),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1688),
.Y(n_1749)
);

INVx8_ASAP7_75t_L g1750 ( 
.A(n_1697),
.Y(n_1750)
);

INVx6_ASAP7_75t_L g1751 ( 
.A(n_1713),
.Y(n_1751)
);

INVx4_ASAP7_75t_L g1752 ( 
.A(n_1684),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1694),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1695),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1689),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1679),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1717),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1703),
.Y(n_1758)
);

CKINVDCx6p67_ASAP7_75t_R g1759 ( 
.A(n_1718),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1706),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1707),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1696),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1708),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1719),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1732),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1721),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1687),
.Y(n_1767)
);

BUFx4f_ASAP7_75t_SL g1768 ( 
.A(n_1686),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1722),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1702),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1728),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1729),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1735),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1712),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1709),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1683),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1700),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1727),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1691),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1698),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1733),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1716),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1699),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1693),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1731),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1705),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1710),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1725),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1724),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1685),
.B(n_1610),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1711),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1704),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1741),
.B(n_1663),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1738),
.A2(n_1662),
.B(n_1673),
.Y(n_1795)
);

AOI222xp33_ASAP7_75t_L g1796 ( 
.A1(n_1787),
.A2(n_1629),
.B1(n_1665),
.B2(n_1666),
.C1(n_1645),
.C2(n_1616),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1740),
.B(n_1651),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1759),
.B(n_1674),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1788),
.B(n_1670),
.C(n_1667),
.D(n_1678),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1745),
.B(n_1664),
.Y(n_1800)
);

NOR3xp33_ASAP7_75t_L g1801 ( 
.A(n_1791),
.B(n_1786),
.C(n_1785),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1784),
.A2(n_1658),
.B1(n_1657),
.B2(n_1615),
.C(n_300),
.Y(n_1802)
);

NAND4xp25_ASAP7_75t_L g1803 ( 
.A(n_1757),
.B(n_301),
.C(n_299),
.D(n_300),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_L g1804 ( 
.A(n_1767),
.B(n_1765),
.C(n_1752),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_L g1805 ( 
.A(n_1793),
.B(n_301),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1737),
.B(n_302),
.C(n_303),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1770),
.B(n_303),
.Y(n_1807)
);

NAND4xp25_ASAP7_75t_L g1808 ( 
.A(n_1755),
.B(n_306),
.C(n_304),
.D(n_305),
.Y(n_1808)
);

OAI211xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1780),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1736),
.B(n_307),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1789),
.B(n_308),
.C(n_309),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1790),
.A2(n_1750),
.B(n_1783),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1792),
.A2(n_1742),
.B1(n_1781),
.B2(n_1746),
.C(n_1774),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_L g1814 ( 
.A(n_1744),
.B(n_312),
.C(n_310),
.D(n_311),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1762),
.B(n_313),
.Y(n_1815)
);

AOI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1739),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1743),
.B(n_315),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1756),
.B(n_1763),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1751),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1768),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_1820)
);

O2A1O1Ixp5_ASAP7_75t_L g1821 ( 
.A1(n_1776),
.A2(n_1771),
.B(n_1775),
.C(n_1777),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1782),
.B(n_322),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1747),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1778),
.A2(n_1779),
.B(n_1749),
.C(n_1753),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1748),
.A2(n_326),
.B(n_323),
.C(n_325),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1754),
.B(n_325),
.Y(n_1826)
);

OAI211xp5_ASAP7_75t_SL g1827 ( 
.A1(n_1794),
.A2(n_1760),
.B(n_1761),
.C(n_1758),
.Y(n_1827)
);

OAI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1808),
.A2(n_1766),
.B1(n_1769),
.B2(n_1764),
.Y(n_1828)
);

AOI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1795),
.A2(n_1773),
.B(n_1772),
.C(n_329),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1804),
.B(n_327),
.C(n_328),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1813),
.A2(n_333),
.B(n_330),
.C(n_332),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1819),
.B(n_1799),
.Y(n_1832)
);

OAI211xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1801),
.A2(n_337),
.B(n_335),
.C(n_336),
.Y(n_1833)
);

AOI21xp33_ASAP7_75t_L g1834 ( 
.A1(n_1797),
.A2(n_1798),
.B(n_1800),
.Y(n_1834)
);

AOI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1821),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.C(n_341),
.Y(n_1835)
);

NOR4xp25_ASAP7_75t_L g1836 ( 
.A(n_1824),
.B(n_342),
.C(n_339),
.D(n_340),
.Y(n_1836)
);

OAI211xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1812),
.A2(n_346),
.B(n_343),
.C(n_345),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1823),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1796),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.C(n_350),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1810),
.Y(n_1840)
);

OAI211xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1802),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_1841)
);

AOI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1825),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.C(n_355),
.Y(n_1842)
);

AO22x2_ASAP7_75t_L g1843 ( 
.A1(n_1811),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1818),
.A2(n_361),
.B1(n_358),
.B2(n_360),
.Y(n_1844)
);

OAI311xp33_ASAP7_75t_L g1845 ( 
.A1(n_1803),
.A2(n_364),
.A3(n_362),
.B1(n_363),
.C1(n_365),
.Y(n_1845)
);

AOI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1809),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_1846)
);

OAI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1805),
.A2(n_367),
.B(n_368),
.Y(n_1847)
);

OAI211xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1816),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_1848)
);

NOR3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1814),
.B(n_372),
.C(n_373),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1806),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1820),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.C(n_379),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1839),
.A2(n_1815),
.B1(n_1817),
.B2(n_1807),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1832),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1841),
.A2(n_1822),
.B1(n_1826),
.B2(n_382),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1847),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1836),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1840),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1838),
.Y(n_1858)
);

NOR2x1_ASAP7_75t_L g1859 ( 
.A(n_1837),
.B(n_385),
.Y(n_1859)
);

NOR2x1_ASAP7_75t_L g1860 ( 
.A(n_1833),
.B(n_387),
.Y(n_1860)
);

NAND4xp75_ASAP7_75t_L g1861 ( 
.A(n_1834),
.B(n_389),
.C(n_387),
.D(n_388),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1830),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1831),
.B(n_391),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1843),
.Y(n_1864)
);

NOR4xp25_ASAP7_75t_L g1865 ( 
.A(n_1827),
.B(n_395),
.C(n_392),
.D(n_393),
.Y(n_1865)
);

NAND2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1844),
.B(n_396),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1865),
.B(n_1829),
.C(n_1835),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1858),
.B(n_1864),
.C(n_1863),
.Y(n_1868)
);

NAND2xp33_ASAP7_75t_SL g1869 ( 
.A(n_1856),
.B(n_1849),
.Y(n_1869)
);

NAND2xp33_ASAP7_75t_L g1870 ( 
.A(n_1859),
.B(n_1850),
.Y(n_1870)
);

XNOR2xp5_ASAP7_75t_L g1871 ( 
.A(n_1854),
.B(n_1846),
.Y(n_1871)
);

AOI211xp5_ASAP7_75t_L g1872 ( 
.A1(n_1868),
.A2(n_1828),
.B(n_1852),
.C(n_1845),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1870),
.Y(n_1873)
);

AOI32xp33_ASAP7_75t_L g1874 ( 
.A1(n_1869),
.A2(n_1860),
.A3(n_1848),
.B1(n_1853),
.B2(n_1857),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1873),
.B(n_1866),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1875),
.Y(n_1876)
);

AOI31xp33_ASAP7_75t_L g1877 ( 
.A1(n_1876),
.A2(n_1872),
.A3(n_1871),
.B(n_1867),
.Y(n_1877)
);

OAI322xp33_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1855),
.A3(n_1862),
.B1(n_1874),
.B2(n_1851),
.C1(n_1861),
.C2(n_1842),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1878),
.A2(n_401),
.B1(n_398),
.B2(n_400),
.Y(n_1879)
);

OAI222xp33_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.C1(n_403),
.C2(n_404),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.C(n_407),
.Y(n_1881)
);

AOI211xp5_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_1882)
);


endmodule