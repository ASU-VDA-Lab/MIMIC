module fake_jpeg_22297_n_299 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_19),
.B1(n_27),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_54),
.A2(n_75),
.B1(n_80),
.B2(n_52),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_19),
.B1(n_20),
.B2(n_27),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_60),
.B(n_73),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_18),
.B1(n_24),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_28),
.B1(n_3),
.B2(n_5),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_38),
.B1(n_25),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_35),
.B1(n_28),
.B2(n_5),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_70),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_26),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_13),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_72),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_27),
.B1(n_31),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_23),
.B1(n_37),
.B2(n_36),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_37),
.B1(n_38),
.B2(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_29),
.B1(n_32),
.B2(n_22),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_2),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_9),
.B(n_12),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_92),
.B1(n_61),
.B2(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_85),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_11),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_14),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_95),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_35),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_91),
.C(n_110),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_35),
.C(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_35),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_100),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_102),
.B1(n_105),
.B2(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_104),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_17),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_59),
.A3(n_52),
.B1(n_17),
.B2(n_14),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_8),
.C(n_9),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_54),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_15),
.B1(n_17),
.B2(n_64),
.Y(n_132)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_117),
.B(n_50),
.C(n_62),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_64),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_13),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_121),
.B(n_132),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_14),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_134),
.C(n_108),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_139),
.Y(n_161)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

BUFx4f_ASAP7_75t_SL g130 ( 
.A(n_112),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_87),
.B(n_115),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_70),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_72),
.B1(n_64),
.B2(n_49),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_109),
.B1(n_83),
.B2(n_93),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_84),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_49),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_62),
.B(n_114),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_117),
.B(n_110),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_62),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_104),
.Y(n_156)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_106),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_156),
.B(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_141),
.B(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_158),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_87),
.B1(n_117),
.B2(n_92),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_163),
.B1(n_148),
.B2(n_134),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_86),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_97),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_169),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_168),
.B(n_136),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_138),
.B(n_143),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_177),
.B(n_179),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_116),
.C(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_140),
.C(n_133),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_85),
.B(n_82),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_147),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_96),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_182),
.C(n_187),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_168),
.B(n_178),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_195),
.B(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_140),
.Y(n_182)
);

XNOR2x2_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_133),
.Y(n_185)
);

XOR2x2_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_120),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_203),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_198),
.B1(n_172),
.B2(n_156),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_185),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_120),
.B(n_127),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_96),
.B1(n_128),
.B2(n_106),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_139),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_129),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_139),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_146),
.B(n_113),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_94),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_174),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_154),
.B1(n_176),
.B2(n_163),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_211),
.A2(n_191),
.B1(n_190),
.B2(n_194),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_187),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_183),
.C(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_216),
.C(n_182),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_183),
.C(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_227),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_224),
.B1(n_199),
.B2(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_170),
.B1(n_169),
.B2(n_152),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_162),
.B(n_160),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_228),
.B(n_202),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_173),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_165),
.B(n_167),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_186),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_235),
.B1(n_207),
.B2(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_223),
.B1(n_221),
.B2(n_213),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_210),
.B(n_212),
.C(n_214),
.D(n_225),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_155),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_240),
.C(n_243),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_195),
.A3(n_164),
.B1(n_180),
.B2(n_187),
.C1(n_199),
.C2(n_190),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_208),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_224),
.B1(n_210),
.B2(n_216),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_195),
.C(n_194),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_164),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_214),
.C(n_211),
.Y(n_256)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_259),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_247),
.B1(n_236),
.B2(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_215),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_217),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_262),
.B(n_247),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_244),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_228),
.C(n_201),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_243),
.C(n_235),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_189),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_268),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_246),
.C(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_267),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_231),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_271),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_250),
.B1(n_253),
.B2(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_204),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_248),
.B1(n_238),
.B2(n_201),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_275),
.A2(n_280),
.B1(n_278),
.B2(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

BUFx4f_ASAP7_75t_SL g278 ( 
.A(n_263),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_255),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_261),
.B(n_230),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.C(n_286),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_264),
.B(n_266),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_271),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_256),
.B1(n_269),
.B2(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_274),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_291),
.B(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_249),
.C(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_200),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_293),
.A3(n_294),
.B1(n_206),
.B2(n_161),
.C1(n_173),
.C2(n_159),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_249),
.B(n_218),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_292),
.A2(n_290),
.B1(n_167),
.B2(n_173),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_296),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_159),
.Y(n_299)
);


endmodule