module real_jpeg_13096_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_5),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_68),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_7),
.A2(n_61),
.B1(n_65),
.B2(n_70),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_70),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_37),
.B(n_38),
.C(n_44),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_8),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_8),
.B(n_41),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_41),
.B(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_26),
.C(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_40),
.B1(n_61),
.B2(n_65),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_166),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_11),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_61),
.B1(n_65),
.B2(n_84),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_84),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_13),
.A2(n_26),
.B1(n_32),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_13),
.A2(n_53),
.B1(n_61),
.B2(n_65),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_61),
.B1(n_65),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_26),
.B1(n_32),
.B2(n_96),
.Y(n_116)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_101),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_19),
.B(n_101),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_48),
.B1(n_71),
.B2(n_72),
.Y(n_20)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_35),
.B2(n_36),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_24),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_24),
.A2(n_29),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_25),
.A2(n_28),
.B1(n_144),
.B2(n_152),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_25),
.A2(n_146),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_26),
.A2(n_32),
.B1(n_90),
.B2(n_91),
.Y(n_93)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_52),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_28),
.B(n_40),
.Y(n_150)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_30),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_29),
.B(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_32),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_37),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_40),
.B(n_93),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_66)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_SL g113 ( 
.A(n_42),
.B(n_63),
.C(n_65),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_58),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_69),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_65),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_64),
.B(n_111),
.C(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_81),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_100),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_94),
.B(n_97),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_99),
.B1(n_106),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_88),
.A2(n_99),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_88),
.A2(n_99),
.B1(n_131),
.B2(n_141),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.C(n_108),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_132),
.B(n_176),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_124),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_130),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_170),
.B(n_175),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_158),
.B(n_169),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_147),
.B(n_157),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_142),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_139),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_153),
.B(n_156),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_164),
.C(n_168),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_174),
.Y(n_175)
);


endmodule