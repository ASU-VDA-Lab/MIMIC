module fake_jpeg_9461_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_3),
.B(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_20),
.C(n_12),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_19),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_18),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_23),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_21),
.B1(n_14),
.B2(n_15),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_58),
.B(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_15),
.B1(n_22),
.B2(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_46),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_36),
.B(n_24),
.C(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_75),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_57),
.C(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_74),
.C(n_71),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_56),
.B1(n_45),
.B2(n_62),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_62),
.B(n_61),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_76),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_89),
.C(n_93),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_74),
.C(n_67),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_67),
.C(n_59),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_85),
.B1(n_80),
.B2(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.C(n_99),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_83),
.B(n_69),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_84),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_64),
.C(n_79),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_94),
.C(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_64),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.C(n_13),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_13),
.B(n_17),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.A3(n_8),
.B1(n_10),
.B2(n_4),
.C1(n_0),
.C2(n_1),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_107),
.A2(n_17),
.B1(n_45),
.B2(n_16),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_108),
.C(n_10),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_47),
.B(n_1),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_0),
.C(n_4),
.Y(n_114)
);


endmodule