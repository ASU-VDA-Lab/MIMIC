module fake_jpeg_9407_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_24),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_10),
.Y(n_35)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_12),
.Y(n_38)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_25),
.B1(n_23),
.B2(n_11),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_1),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_37),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_10),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_22),
.A2(n_16),
.B1(n_11),
.B2(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_19),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_31),
.C(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_15),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_28),
.B(n_33),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_51),
.C(n_58),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_41),
.C(n_15),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_3),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_54),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_34),
.C(n_30),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_60),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_67),
.C(n_68),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_56),
.Y(n_72)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_34),
.C(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_46),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_49),
.B(n_52),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_29),
.C(n_32),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.C(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_51),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_26),
.Y(n_82)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_55),
.B(n_59),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_59),
.B1(n_25),
.B2(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_27),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.C(n_18),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_47),
.Y(n_80)
);

AO221x1_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_65),
.B1(n_26),
.B2(n_18),
.C(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.C(n_72),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_80),
.B1(n_23),
.B2(n_27),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_27),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_93),
.C(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_85),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_83),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_9),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_4),
.C(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_8),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_100),
.C(n_7),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);


endmodule