module fake_jpeg_2288_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_58),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_48),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_56),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_2),
.CON(n_57),
.SN(n_57)
);

OR2x4_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_57),
.B(n_53),
.C(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_73),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_42),
.C(n_44),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_35),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_40),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_66),
.B(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_87),
.B1(n_66),
.B2(n_52),
.Y(n_100)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_58),
.B1(n_40),
.B2(n_39),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_43),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_66),
.Y(n_101)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_103),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_104),
.B1(n_111),
.B2(n_6),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_41),
.B1(n_38),
.B2(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_3),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_5),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_21),
.B(n_34),
.C(n_33),
.D(n_32),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_110),
.B(n_113),
.C(n_22),
.D(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_41),
.B1(n_8),
.B2(n_9),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_100),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_122),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_20),
.C(n_29),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_125),
.C(n_111),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.C(n_31),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_24),
.C(n_13),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_127),
.B(n_119),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_98),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_123),
.B1(n_115),
.B2(n_118),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_130),
.C(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_122),
.C(n_14),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_136),
.B(n_16),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_18),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_25),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_26),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_27),
.Y(n_142)
);


endmodule